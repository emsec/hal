library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

entity sha_256_core is
  port (
clk : in STD_LOGIC := 'X'; 
  data_ready : in STD_LOGIC := 'X'; 
  msg_block_in_0 : in STD_LOGIC := 'X'; 
  msg_block_in_1 : in STD_LOGIC := 'X'; 
  msg_block_in_10 : in STD_LOGIC := 'X'; 
  msg_block_in_100 : in STD_LOGIC := 'X'; 
  msg_block_in_101 : in STD_LOGIC := 'X'; 
  msg_block_in_102 : in STD_LOGIC := 'X'; 
  msg_block_in_103 : in STD_LOGIC := 'X'; 
  msg_block_in_104 : in STD_LOGIC := 'X'; 
  msg_block_in_105 : in STD_LOGIC := 'X'; 
  msg_block_in_106 : in STD_LOGIC := 'X'; 
  msg_block_in_107 : in STD_LOGIC := 'X'; 
  msg_block_in_108 : in STD_LOGIC := 'X'; 
  msg_block_in_109 : in STD_LOGIC := 'X'; 
  msg_block_in_11 : in STD_LOGIC := 'X'; 
  msg_block_in_110 : in STD_LOGIC := 'X'; 
  msg_block_in_111 : in STD_LOGIC := 'X'; 
  msg_block_in_112 : in STD_LOGIC := 'X'; 
  msg_block_in_113 : in STD_LOGIC := 'X'; 
  msg_block_in_114 : in STD_LOGIC := 'X'; 
  msg_block_in_115 : in STD_LOGIC := 'X'; 
  msg_block_in_116 : in STD_LOGIC := 'X'; 
  msg_block_in_117 : in STD_LOGIC := 'X'; 
  msg_block_in_118 : in STD_LOGIC := 'X'; 
  msg_block_in_119 : in STD_LOGIC := 'X'; 
  msg_block_in_12 : in STD_LOGIC := 'X'; 
  msg_block_in_120 : in STD_LOGIC := 'X'; 
  msg_block_in_121 : in STD_LOGIC := 'X'; 
  msg_block_in_122 : in STD_LOGIC := 'X'; 
  msg_block_in_123 : in STD_LOGIC := 'X'; 
  msg_block_in_124 : in STD_LOGIC := 'X'; 
  msg_block_in_125 : in STD_LOGIC := 'X'; 
  msg_block_in_126 : in STD_LOGIC := 'X'; 
  msg_block_in_127 : in STD_LOGIC := 'X'; 
  msg_block_in_128 : in STD_LOGIC := 'X'; 
  msg_block_in_129 : in STD_LOGIC := 'X'; 
  msg_block_in_13 : in STD_LOGIC := 'X'; 
  msg_block_in_130 : in STD_LOGIC := 'X'; 
  msg_block_in_131 : in STD_LOGIC := 'X'; 
  msg_block_in_132 : in STD_LOGIC := 'X'; 
  msg_block_in_133 : in STD_LOGIC := 'X'; 
  msg_block_in_134 : in STD_LOGIC := 'X'; 
  msg_block_in_135 : in STD_LOGIC := 'X'; 
  msg_block_in_136 : in STD_LOGIC := 'X'; 
  msg_block_in_137 : in STD_LOGIC := 'X'; 
  msg_block_in_138 : in STD_LOGIC := 'X'; 
  msg_block_in_139 : in STD_LOGIC := 'X'; 
  msg_block_in_14 : in STD_LOGIC := 'X'; 
  msg_block_in_140 : in STD_LOGIC := 'X'; 
  msg_block_in_141 : in STD_LOGIC := 'X'; 
  msg_block_in_142 : in STD_LOGIC := 'X'; 
  msg_block_in_143 : in STD_LOGIC := 'X'; 
  msg_block_in_144 : in STD_LOGIC := 'X'; 
  msg_block_in_145 : in STD_LOGIC := 'X'; 
  msg_block_in_146 : in STD_LOGIC := 'X'; 
  msg_block_in_147 : in STD_LOGIC := 'X'; 
  msg_block_in_148 : in STD_LOGIC := 'X'; 
  msg_block_in_149 : in STD_LOGIC := 'X'; 
  msg_block_in_15 : in STD_LOGIC := 'X'; 
  msg_block_in_150 : in STD_LOGIC := 'X'; 
  msg_block_in_151 : in STD_LOGIC := 'X'; 
  msg_block_in_152 : in STD_LOGIC := 'X'; 
  msg_block_in_153 : in STD_LOGIC := 'X'; 
  msg_block_in_154 : in STD_LOGIC := 'X'; 
  msg_block_in_155 : in STD_LOGIC := 'X'; 
  msg_block_in_156 : in STD_LOGIC := 'X'; 
  msg_block_in_157 : in STD_LOGIC := 'X'; 
  msg_block_in_158 : in STD_LOGIC := 'X'; 
  msg_block_in_159 : in STD_LOGIC := 'X'; 
  msg_block_in_16 : in STD_LOGIC := 'X'; 
  msg_block_in_160 : in STD_LOGIC := 'X'; 
  msg_block_in_161 : in STD_LOGIC := 'X'; 
  msg_block_in_162 : in STD_LOGIC := 'X'; 
  msg_block_in_163 : in STD_LOGIC := 'X'; 
  msg_block_in_164 : in STD_LOGIC := 'X'; 
  msg_block_in_165 : in STD_LOGIC := 'X'; 
  msg_block_in_166 : in STD_LOGIC := 'X'; 
  msg_block_in_167 : in STD_LOGIC := 'X'; 
  msg_block_in_168 : in STD_LOGIC := 'X'; 
  msg_block_in_169 : in STD_LOGIC := 'X'; 
  msg_block_in_17 : in STD_LOGIC := 'X'; 
  msg_block_in_170 : in STD_LOGIC := 'X'; 
  msg_block_in_171 : in STD_LOGIC := 'X'; 
  msg_block_in_172 : in STD_LOGIC := 'X'; 
  msg_block_in_173 : in STD_LOGIC := 'X'; 
  msg_block_in_174 : in STD_LOGIC := 'X'; 
  msg_block_in_175 : in STD_LOGIC := 'X'; 
  msg_block_in_176 : in STD_LOGIC := 'X'; 
  msg_block_in_177 : in STD_LOGIC := 'X'; 
  msg_block_in_178 : in STD_LOGIC := 'X'; 
  msg_block_in_179 : in STD_LOGIC := 'X'; 
  msg_block_in_18 : in STD_LOGIC := 'X'; 
  msg_block_in_180 : in STD_LOGIC := 'X'; 
  msg_block_in_181 : in STD_LOGIC := 'X'; 
  msg_block_in_182 : in STD_LOGIC := 'X'; 
  msg_block_in_183 : in STD_LOGIC := 'X'; 
  msg_block_in_184 : in STD_LOGIC := 'X'; 
  msg_block_in_185 : in STD_LOGIC := 'X'; 
  msg_block_in_186 : in STD_LOGIC := 'X'; 
  msg_block_in_187 : in STD_LOGIC := 'X'; 
  msg_block_in_188 : in STD_LOGIC := 'X'; 
  msg_block_in_189 : in STD_LOGIC := 'X'; 
  msg_block_in_19 : in STD_LOGIC := 'X'; 
  msg_block_in_190 : in STD_LOGIC := 'X'; 
  msg_block_in_191 : in STD_LOGIC := 'X'; 
  msg_block_in_192 : in STD_LOGIC := 'X'; 
  msg_block_in_193 : in STD_LOGIC := 'X'; 
  msg_block_in_194 : in STD_LOGIC := 'X'; 
  msg_block_in_195 : in STD_LOGIC := 'X'; 
  msg_block_in_196 : in STD_LOGIC := 'X'; 
  msg_block_in_197 : in STD_LOGIC := 'X'; 
  msg_block_in_198 : in STD_LOGIC := 'X'; 
  msg_block_in_199 : in STD_LOGIC := 'X'; 
  msg_block_in_2 : in STD_LOGIC := 'X'; 
  msg_block_in_20 : in STD_LOGIC := 'X'; 
  msg_block_in_200 : in STD_LOGIC := 'X'; 
  msg_block_in_201 : in STD_LOGIC := 'X'; 
  msg_block_in_202 : in STD_LOGIC := 'X'; 
  msg_block_in_203 : in STD_LOGIC := 'X'; 
  msg_block_in_204 : in STD_LOGIC := 'X'; 
  msg_block_in_205 : in STD_LOGIC := 'X'; 
  msg_block_in_206 : in STD_LOGIC := 'X'; 
  msg_block_in_207 : in STD_LOGIC := 'X'; 
  msg_block_in_208 : in STD_LOGIC := 'X'; 
  msg_block_in_209 : in STD_LOGIC := 'X'; 
  msg_block_in_21 : in STD_LOGIC := 'X'; 
  msg_block_in_210 : in STD_LOGIC := 'X'; 
  msg_block_in_211 : in STD_LOGIC := 'X'; 
  msg_block_in_212 : in STD_LOGIC := 'X'; 
  msg_block_in_213 : in STD_LOGIC := 'X'; 
  msg_block_in_214 : in STD_LOGIC := 'X'; 
  msg_block_in_215 : in STD_LOGIC := 'X'; 
  msg_block_in_216 : in STD_LOGIC := 'X'; 
  msg_block_in_217 : in STD_LOGIC := 'X'; 
  msg_block_in_218 : in STD_LOGIC := 'X'; 
  msg_block_in_219 : in STD_LOGIC := 'X'; 
  msg_block_in_22 : in STD_LOGIC := 'X'; 
  msg_block_in_220 : in STD_LOGIC := 'X'; 
  msg_block_in_221 : in STD_LOGIC := 'X'; 
  msg_block_in_222 : in STD_LOGIC := 'X'; 
  msg_block_in_223 : in STD_LOGIC := 'X'; 
  msg_block_in_224 : in STD_LOGIC := 'X'; 
  msg_block_in_225 : in STD_LOGIC := 'X'; 
  msg_block_in_226 : in STD_LOGIC := 'X'; 
  msg_block_in_227 : in STD_LOGIC := 'X'; 
  msg_block_in_228 : in STD_LOGIC := 'X'; 
  msg_block_in_229 : in STD_LOGIC := 'X'; 
  msg_block_in_23 : in STD_LOGIC := 'X'; 
  msg_block_in_230 : in STD_LOGIC := 'X'; 
  msg_block_in_231 : in STD_LOGIC := 'X'; 
  msg_block_in_232 : in STD_LOGIC := 'X'; 
  msg_block_in_233 : in STD_LOGIC := 'X'; 
  msg_block_in_234 : in STD_LOGIC := 'X'; 
  msg_block_in_235 : in STD_LOGIC := 'X'; 
  msg_block_in_236 : in STD_LOGIC := 'X'; 
  msg_block_in_237 : in STD_LOGIC := 'X'; 
  msg_block_in_238 : in STD_LOGIC := 'X'; 
  msg_block_in_239 : in STD_LOGIC := 'X'; 
  msg_block_in_24 : in STD_LOGIC := 'X'; 
  msg_block_in_240 : in STD_LOGIC := 'X'; 
  msg_block_in_241 : in STD_LOGIC := 'X'; 
  msg_block_in_242 : in STD_LOGIC := 'X'; 
  msg_block_in_243 : in STD_LOGIC := 'X'; 
  msg_block_in_244 : in STD_LOGIC := 'X'; 
  msg_block_in_245 : in STD_LOGIC := 'X'; 
  msg_block_in_246 : in STD_LOGIC := 'X'; 
  msg_block_in_247 : in STD_LOGIC := 'X'; 
  msg_block_in_248 : in STD_LOGIC := 'X'; 
  msg_block_in_249 : in STD_LOGIC := 'X'; 
  msg_block_in_25 : in STD_LOGIC := 'X'; 
  msg_block_in_250 : in STD_LOGIC := 'X'; 
  msg_block_in_251 : in STD_LOGIC := 'X'; 
  msg_block_in_252 : in STD_LOGIC := 'X'; 
  msg_block_in_253 : in STD_LOGIC := 'X'; 
  msg_block_in_254 : in STD_LOGIC := 'X'; 
  msg_block_in_255 : in STD_LOGIC := 'X'; 
  msg_block_in_256 : in STD_LOGIC := 'X'; 
  msg_block_in_257 : in STD_LOGIC := 'X'; 
  msg_block_in_258 : in STD_LOGIC := 'X'; 
  msg_block_in_259 : in STD_LOGIC := 'X'; 
  msg_block_in_26 : in STD_LOGIC := 'X'; 
  msg_block_in_260 : in STD_LOGIC := 'X'; 
  msg_block_in_261 : in STD_LOGIC := 'X'; 
  msg_block_in_262 : in STD_LOGIC := 'X'; 
  msg_block_in_263 : in STD_LOGIC := 'X'; 
  msg_block_in_264 : in STD_LOGIC := 'X'; 
  msg_block_in_265 : in STD_LOGIC := 'X'; 
  msg_block_in_266 : in STD_LOGIC := 'X'; 
  msg_block_in_267 : in STD_LOGIC := 'X'; 
  msg_block_in_268 : in STD_LOGIC := 'X'; 
  msg_block_in_269 : in STD_LOGIC := 'X'; 
  msg_block_in_27 : in STD_LOGIC := 'X'; 
  msg_block_in_270 : in STD_LOGIC := 'X'; 
  msg_block_in_271 : in STD_LOGIC := 'X'; 
  msg_block_in_272 : in STD_LOGIC := 'X'; 
  msg_block_in_273 : in STD_LOGIC := 'X'; 
  msg_block_in_274 : in STD_LOGIC := 'X'; 
  msg_block_in_275 : in STD_LOGIC := 'X'; 
  msg_block_in_276 : in STD_LOGIC := 'X'; 
  msg_block_in_277 : in STD_LOGIC := 'X'; 
  msg_block_in_278 : in STD_LOGIC := 'X'; 
  msg_block_in_279 : in STD_LOGIC := 'X'; 
  msg_block_in_28 : in STD_LOGIC := 'X'; 
  msg_block_in_280 : in STD_LOGIC := 'X'; 
  msg_block_in_281 : in STD_LOGIC := 'X'; 
  msg_block_in_282 : in STD_LOGIC := 'X'; 
  msg_block_in_283 : in STD_LOGIC := 'X'; 
  msg_block_in_284 : in STD_LOGIC := 'X'; 
  msg_block_in_285 : in STD_LOGIC := 'X'; 
  msg_block_in_286 : in STD_LOGIC := 'X'; 
  msg_block_in_287 : in STD_LOGIC := 'X'; 
  msg_block_in_288 : in STD_LOGIC := 'X'; 
  msg_block_in_289 : in STD_LOGIC := 'X'; 
  msg_block_in_29 : in STD_LOGIC := 'X'; 
  msg_block_in_290 : in STD_LOGIC := 'X'; 
  msg_block_in_291 : in STD_LOGIC := 'X'; 
  msg_block_in_292 : in STD_LOGIC := 'X'; 
  msg_block_in_293 : in STD_LOGIC := 'X'; 
  msg_block_in_294 : in STD_LOGIC := 'X'; 
  msg_block_in_295 : in STD_LOGIC := 'X'; 
  msg_block_in_296 : in STD_LOGIC := 'X'; 
  msg_block_in_297 : in STD_LOGIC := 'X'; 
  msg_block_in_298 : in STD_LOGIC := 'X'; 
  msg_block_in_299 : in STD_LOGIC := 'X'; 
  msg_block_in_3 : in STD_LOGIC := 'X'; 
  msg_block_in_30 : in STD_LOGIC := 'X'; 
  msg_block_in_300 : in STD_LOGIC := 'X'; 
  msg_block_in_301 : in STD_LOGIC := 'X'; 
  msg_block_in_302 : in STD_LOGIC := 'X'; 
  msg_block_in_303 : in STD_LOGIC := 'X'; 
  msg_block_in_304 : in STD_LOGIC := 'X'; 
  msg_block_in_305 : in STD_LOGIC := 'X'; 
  msg_block_in_306 : in STD_LOGIC := 'X'; 
  msg_block_in_307 : in STD_LOGIC := 'X'; 
  msg_block_in_308 : in STD_LOGIC := 'X'; 
  msg_block_in_309 : in STD_LOGIC := 'X'; 
  msg_block_in_31 : in STD_LOGIC := 'X'; 
  msg_block_in_310 : in STD_LOGIC := 'X'; 
  msg_block_in_311 : in STD_LOGIC := 'X'; 
  msg_block_in_312 : in STD_LOGIC := 'X'; 
  msg_block_in_313 : in STD_LOGIC := 'X'; 
  msg_block_in_314 : in STD_LOGIC := 'X'; 
  msg_block_in_315 : in STD_LOGIC := 'X'; 
  msg_block_in_316 : in STD_LOGIC := 'X'; 
  msg_block_in_317 : in STD_LOGIC := 'X'; 
  msg_block_in_318 : in STD_LOGIC := 'X'; 
  msg_block_in_319 : in STD_LOGIC := 'X'; 
  msg_block_in_32 : in STD_LOGIC := 'X'; 
  msg_block_in_320 : in STD_LOGIC := 'X'; 
  msg_block_in_321 : in STD_LOGIC := 'X'; 
  msg_block_in_322 : in STD_LOGIC := 'X'; 
  msg_block_in_323 : in STD_LOGIC := 'X'; 
  msg_block_in_324 : in STD_LOGIC := 'X'; 
  msg_block_in_325 : in STD_LOGIC := 'X'; 
  msg_block_in_326 : in STD_LOGIC := 'X'; 
  msg_block_in_327 : in STD_LOGIC := 'X'; 
  msg_block_in_328 : in STD_LOGIC := 'X'; 
  msg_block_in_329 : in STD_LOGIC := 'X'; 
  msg_block_in_33 : in STD_LOGIC := 'X'; 
  msg_block_in_330 : in STD_LOGIC := 'X'; 
  msg_block_in_331 : in STD_LOGIC := 'X'; 
  msg_block_in_332 : in STD_LOGIC := 'X'; 
  msg_block_in_333 : in STD_LOGIC := 'X'; 
  msg_block_in_334 : in STD_LOGIC := 'X'; 
  msg_block_in_335 : in STD_LOGIC := 'X'; 
  msg_block_in_336 : in STD_LOGIC := 'X'; 
  msg_block_in_337 : in STD_LOGIC := 'X'; 
  msg_block_in_338 : in STD_LOGIC := 'X'; 
  msg_block_in_339 : in STD_LOGIC := 'X'; 
  msg_block_in_34 : in STD_LOGIC := 'X'; 
  msg_block_in_340 : in STD_LOGIC := 'X'; 
  msg_block_in_341 : in STD_LOGIC := 'X'; 
  msg_block_in_342 : in STD_LOGIC := 'X'; 
  msg_block_in_343 : in STD_LOGIC := 'X'; 
  msg_block_in_344 : in STD_LOGIC := 'X'; 
  msg_block_in_345 : in STD_LOGIC := 'X'; 
  msg_block_in_346 : in STD_LOGIC := 'X'; 
  msg_block_in_347 : in STD_LOGIC := 'X'; 
  msg_block_in_348 : in STD_LOGIC := 'X'; 
  msg_block_in_349 : in STD_LOGIC := 'X'; 
  msg_block_in_35 : in STD_LOGIC := 'X'; 
  msg_block_in_350 : in STD_LOGIC := 'X'; 
  msg_block_in_351 : in STD_LOGIC := 'X'; 
  msg_block_in_352 : in STD_LOGIC := 'X'; 
  msg_block_in_353 : in STD_LOGIC := 'X'; 
  msg_block_in_354 : in STD_LOGIC := 'X'; 
  msg_block_in_355 : in STD_LOGIC := 'X'; 
  msg_block_in_356 : in STD_LOGIC := 'X'; 
  msg_block_in_357 : in STD_LOGIC := 'X'; 
  msg_block_in_358 : in STD_LOGIC := 'X'; 
  msg_block_in_359 : in STD_LOGIC := 'X'; 
  msg_block_in_36 : in STD_LOGIC := 'X'; 
  msg_block_in_360 : in STD_LOGIC := 'X'; 
  msg_block_in_361 : in STD_LOGIC := 'X'; 
  msg_block_in_362 : in STD_LOGIC := 'X'; 
  msg_block_in_363 : in STD_LOGIC := 'X'; 
  msg_block_in_364 : in STD_LOGIC := 'X'; 
  msg_block_in_365 : in STD_LOGIC := 'X'; 
  msg_block_in_366 : in STD_LOGIC := 'X'; 
  msg_block_in_367 : in STD_LOGIC := 'X'; 
  msg_block_in_368 : in STD_LOGIC := 'X'; 
  msg_block_in_369 : in STD_LOGIC := 'X'; 
  msg_block_in_37 : in STD_LOGIC := 'X'; 
  msg_block_in_370 : in STD_LOGIC := 'X'; 
  msg_block_in_371 : in STD_LOGIC := 'X'; 
  msg_block_in_372 : in STD_LOGIC := 'X'; 
  msg_block_in_373 : in STD_LOGIC := 'X'; 
  msg_block_in_374 : in STD_LOGIC := 'X'; 
  msg_block_in_375 : in STD_LOGIC := 'X'; 
  msg_block_in_376 : in STD_LOGIC := 'X'; 
  msg_block_in_377 : in STD_LOGIC := 'X'; 
  msg_block_in_378 : in STD_LOGIC := 'X'; 
  msg_block_in_379 : in STD_LOGIC := 'X'; 
  msg_block_in_38 : in STD_LOGIC := 'X'; 
  msg_block_in_380 : in STD_LOGIC := 'X'; 
  msg_block_in_381 : in STD_LOGIC := 'X'; 
  msg_block_in_382 : in STD_LOGIC := 'X'; 
  msg_block_in_383 : in STD_LOGIC := 'X'; 
  msg_block_in_384 : in STD_LOGIC := 'X'; 
  msg_block_in_385 : in STD_LOGIC := 'X'; 
  msg_block_in_386 : in STD_LOGIC := 'X'; 
  msg_block_in_387 : in STD_LOGIC := 'X'; 
  msg_block_in_388 : in STD_LOGIC := 'X'; 
  msg_block_in_389 : in STD_LOGIC := 'X'; 
  msg_block_in_39 : in STD_LOGIC := 'X'; 
  msg_block_in_390 : in STD_LOGIC := 'X'; 
  msg_block_in_391 : in STD_LOGIC := 'X'; 
  msg_block_in_392 : in STD_LOGIC := 'X'; 
  msg_block_in_393 : in STD_LOGIC := 'X'; 
  msg_block_in_394 : in STD_LOGIC := 'X'; 
  msg_block_in_395 : in STD_LOGIC := 'X'; 
  msg_block_in_396 : in STD_LOGIC := 'X'; 
  msg_block_in_397 : in STD_LOGIC := 'X'; 
  msg_block_in_398 : in STD_LOGIC := 'X'; 
  msg_block_in_399 : in STD_LOGIC := 'X'; 
  msg_block_in_4 : in STD_LOGIC := 'X'; 
  msg_block_in_40 : in STD_LOGIC := 'X'; 
  msg_block_in_400 : in STD_LOGIC := 'X'; 
  msg_block_in_401 : in STD_LOGIC := 'X'; 
  msg_block_in_402 : in STD_LOGIC := 'X'; 
  msg_block_in_403 : in STD_LOGIC := 'X'; 
  msg_block_in_404 : in STD_LOGIC := 'X'; 
  msg_block_in_405 : in STD_LOGIC := 'X'; 
  msg_block_in_406 : in STD_LOGIC := 'X'; 
  msg_block_in_407 : in STD_LOGIC := 'X'; 
  msg_block_in_408 : in STD_LOGIC := 'X'; 
  msg_block_in_409 : in STD_LOGIC := 'X'; 
  msg_block_in_41 : in STD_LOGIC := 'X'; 
  msg_block_in_410 : in STD_LOGIC := 'X'; 
  msg_block_in_411 : in STD_LOGIC := 'X'; 
  msg_block_in_412 : in STD_LOGIC := 'X'; 
  msg_block_in_413 : in STD_LOGIC := 'X'; 
  msg_block_in_414 : in STD_LOGIC := 'X'; 
  msg_block_in_415 : in STD_LOGIC := 'X'; 
  msg_block_in_416 : in STD_LOGIC := 'X'; 
  msg_block_in_417 : in STD_LOGIC := 'X'; 
  msg_block_in_418 : in STD_LOGIC := 'X'; 
  msg_block_in_419 : in STD_LOGIC := 'X'; 
  msg_block_in_42 : in STD_LOGIC := 'X'; 
  msg_block_in_420 : in STD_LOGIC := 'X'; 
  msg_block_in_421 : in STD_LOGIC := 'X'; 
  msg_block_in_422 : in STD_LOGIC := 'X'; 
  msg_block_in_423 : in STD_LOGIC := 'X'; 
  msg_block_in_424 : in STD_LOGIC := 'X'; 
  msg_block_in_425 : in STD_LOGIC := 'X'; 
  msg_block_in_426 : in STD_LOGIC := 'X'; 
  msg_block_in_427 : in STD_LOGIC := 'X'; 
  msg_block_in_428 : in STD_LOGIC := 'X'; 
  msg_block_in_429 : in STD_LOGIC := 'X'; 
  msg_block_in_43 : in STD_LOGIC := 'X'; 
  msg_block_in_430 : in STD_LOGIC := 'X'; 
  msg_block_in_431 : in STD_LOGIC := 'X'; 
  msg_block_in_432 : in STD_LOGIC := 'X'; 
  msg_block_in_433 : in STD_LOGIC := 'X'; 
  msg_block_in_434 : in STD_LOGIC := 'X'; 
  msg_block_in_435 : in STD_LOGIC := 'X'; 
  msg_block_in_436 : in STD_LOGIC := 'X'; 
  msg_block_in_437 : in STD_LOGIC := 'X'; 
  msg_block_in_438 : in STD_LOGIC := 'X'; 
  msg_block_in_439 : in STD_LOGIC := 'X'; 
  msg_block_in_44 : in STD_LOGIC := 'X'; 
  msg_block_in_440 : in STD_LOGIC := 'X'; 
  msg_block_in_441 : in STD_LOGIC := 'X'; 
  msg_block_in_442 : in STD_LOGIC := 'X'; 
  msg_block_in_443 : in STD_LOGIC := 'X'; 
  msg_block_in_444 : in STD_LOGIC := 'X'; 
  msg_block_in_445 : in STD_LOGIC := 'X'; 
  msg_block_in_446 : in STD_LOGIC := 'X'; 
  msg_block_in_447 : in STD_LOGIC := 'X'; 
  msg_block_in_448 : in STD_LOGIC := 'X'; 
  msg_block_in_449 : in STD_LOGIC := 'X'; 
  msg_block_in_45 : in STD_LOGIC := 'X'; 
  msg_block_in_450 : in STD_LOGIC := 'X'; 
  msg_block_in_451 : in STD_LOGIC := 'X'; 
  msg_block_in_452 : in STD_LOGIC := 'X'; 
  msg_block_in_453 : in STD_LOGIC := 'X'; 
  msg_block_in_454 : in STD_LOGIC := 'X'; 
  msg_block_in_455 : in STD_LOGIC := 'X'; 
  msg_block_in_456 : in STD_LOGIC := 'X'; 
  msg_block_in_457 : in STD_LOGIC := 'X'; 
  msg_block_in_458 : in STD_LOGIC := 'X'; 
  msg_block_in_459 : in STD_LOGIC := 'X'; 
  msg_block_in_46 : in STD_LOGIC := 'X'; 
  msg_block_in_460 : in STD_LOGIC := 'X'; 
  msg_block_in_461 : in STD_LOGIC := 'X'; 
  msg_block_in_462 : in STD_LOGIC := 'X'; 
  msg_block_in_463 : in STD_LOGIC := 'X'; 
  msg_block_in_464 : in STD_LOGIC := 'X'; 
  msg_block_in_465 : in STD_LOGIC := 'X'; 
  msg_block_in_466 : in STD_LOGIC := 'X'; 
  msg_block_in_467 : in STD_LOGIC := 'X'; 
  msg_block_in_468 : in STD_LOGIC := 'X'; 
  msg_block_in_469 : in STD_LOGIC := 'X'; 
  msg_block_in_47 : in STD_LOGIC := 'X'; 
  msg_block_in_470 : in STD_LOGIC := 'X'; 
  msg_block_in_471 : in STD_LOGIC := 'X'; 
  msg_block_in_472 : in STD_LOGIC := 'X'; 
  msg_block_in_473 : in STD_LOGIC := 'X'; 
  msg_block_in_474 : in STD_LOGIC := 'X'; 
  msg_block_in_475 : in STD_LOGIC := 'X'; 
  msg_block_in_476 : in STD_LOGIC := 'X'; 
  msg_block_in_477 : in STD_LOGIC := 'X'; 
  msg_block_in_478 : in STD_LOGIC := 'X'; 
  msg_block_in_479 : in STD_LOGIC := 'X'; 
  msg_block_in_48 : in STD_LOGIC := 'X'; 
  msg_block_in_480 : in STD_LOGIC := 'X'; 
  msg_block_in_481 : in STD_LOGIC := 'X'; 
  msg_block_in_482 : in STD_LOGIC := 'X'; 
  msg_block_in_483 : in STD_LOGIC := 'X'; 
  msg_block_in_484 : in STD_LOGIC := 'X'; 
  msg_block_in_485 : in STD_LOGIC := 'X'; 
  msg_block_in_486 : in STD_LOGIC := 'X'; 
  msg_block_in_487 : in STD_LOGIC := 'X'; 
  msg_block_in_488 : in STD_LOGIC := 'X'; 
  msg_block_in_489 : in STD_LOGIC := 'X'; 
  msg_block_in_49 : in STD_LOGIC := 'X'; 
  msg_block_in_490 : in STD_LOGIC := 'X'; 
  msg_block_in_491 : in STD_LOGIC := 'X'; 
  msg_block_in_492 : in STD_LOGIC := 'X'; 
  msg_block_in_493 : in STD_LOGIC := 'X'; 
  msg_block_in_494 : in STD_LOGIC := 'X'; 
  msg_block_in_495 : in STD_LOGIC := 'X'; 
  msg_block_in_496 : in STD_LOGIC := 'X'; 
  msg_block_in_497 : in STD_LOGIC := 'X'; 
  msg_block_in_498 : in STD_LOGIC := 'X'; 
  msg_block_in_499 : in STD_LOGIC := 'X'; 
  msg_block_in_5 : in STD_LOGIC := 'X'; 
  msg_block_in_50 : in STD_LOGIC := 'X'; 
  msg_block_in_500 : in STD_LOGIC := 'X'; 
  msg_block_in_501 : in STD_LOGIC := 'X'; 
  msg_block_in_502 : in STD_LOGIC := 'X'; 
  msg_block_in_503 : in STD_LOGIC := 'X'; 
  msg_block_in_504 : in STD_LOGIC := 'X'; 
  msg_block_in_505 : in STD_LOGIC := 'X'; 
  msg_block_in_506 : in STD_LOGIC := 'X'; 
  msg_block_in_507 : in STD_LOGIC := 'X'; 
  msg_block_in_508 : in STD_LOGIC := 'X'; 
  msg_block_in_509 : in STD_LOGIC := 'X'; 
  msg_block_in_51 : in STD_LOGIC := 'X'; 
  msg_block_in_510 : in STD_LOGIC := 'X'; 
  msg_block_in_511 : in STD_LOGIC := 'X'; 
  msg_block_in_52 : in STD_LOGIC := 'X'; 
  msg_block_in_53 : in STD_LOGIC := 'X'; 
  msg_block_in_54 : in STD_LOGIC := 'X'; 
  msg_block_in_55 : in STD_LOGIC := 'X'; 
  msg_block_in_56 : in STD_LOGIC := 'X'; 
  msg_block_in_57 : in STD_LOGIC := 'X'; 
  msg_block_in_58 : in STD_LOGIC := 'X'; 
  msg_block_in_59 : in STD_LOGIC := 'X'; 
  msg_block_in_6 : in STD_LOGIC := 'X'; 
  msg_block_in_60 : in STD_LOGIC := 'X'; 
  msg_block_in_61 : in STD_LOGIC := 'X'; 
  msg_block_in_62 : in STD_LOGIC := 'X'; 
  msg_block_in_63 : in STD_LOGIC := 'X'; 
  msg_block_in_64 : in STD_LOGIC := 'X'; 
  msg_block_in_65 : in STD_LOGIC := 'X'; 
  msg_block_in_66 : in STD_LOGIC := 'X'; 
  msg_block_in_67 : in STD_LOGIC := 'X'; 
  msg_block_in_68 : in STD_LOGIC := 'X'; 
  msg_block_in_69 : in STD_LOGIC := 'X'; 
  msg_block_in_7 : in STD_LOGIC := 'X'; 
  msg_block_in_70 : in STD_LOGIC := 'X'; 
  msg_block_in_71 : in STD_LOGIC := 'X'; 
  msg_block_in_72 : in STD_LOGIC := 'X'; 
  msg_block_in_73 : in STD_LOGIC := 'X'; 
  msg_block_in_74 : in STD_LOGIC := 'X'; 
  msg_block_in_75 : in STD_LOGIC := 'X'; 
  msg_block_in_76 : in STD_LOGIC := 'X'; 
  msg_block_in_77 : in STD_LOGIC := 'X'; 
  msg_block_in_78 : in STD_LOGIC := 'X'; 
  msg_block_in_79 : in STD_LOGIC := 'X'; 
  msg_block_in_8 : in STD_LOGIC := 'X'; 
  msg_block_in_80 : in STD_LOGIC := 'X'; 
  msg_block_in_81 : in STD_LOGIC := 'X'; 
  msg_block_in_82 : in STD_LOGIC := 'X'; 
  msg_block_in_83 : in STD_LOGIC := 'X'; 
  msg_block_in_84 : in STD_LOGIC := 'X'; 
  msg_block_in_85 : in STD_LOGIC := 'X'; 
  msg_block_in_86 : in STD_LOGIC := 'X'; 
  msg_block_in_87 : in STD_LOGIC := 'X'; 
  msg_block_in_88 : in STD_LOGIC := 'X'; 
  msg_block_in_89 : in STD_LOGIC := 'X'; 
  msg_block_in_9 : in STD_LOGIC := 'X'; 
  msg_block_in_90 : in STD_LOGIC := 'X'; 
  msg_block_in_91 : in STD_LOGIC := 'X'; 
  msg_block_in_92 : in STD_LOGIC := 'X'; 
  msg_block_in_93 : in STD_LOGIC := 'X'; 
  msg_block_in_94 : in STD_LOGIC := 'X'; 
  msg_block_in_95 : in STD_LOGIC := 'X'; 
  msg_block_in_96 : in STD_LOGIC := 'X'; 
  msg_block_in_97 : in STD_LOGIC := 'X'; 
  msg_block_in_98 : in STD_LOGIC := 'X'; 
  msg_block_in_99 : in STD_LOGIC := 'X'; 
  rst : in STD_LOGIC := 'X'; 
  data_out_0 : out STD_LOGIC; 
  data_out_1 : out STD_LOGIC; 
  data_out_10 : out STD_LOGIC; 
  data_out_100 : out STD_LOGIC; 
  data_out_101 : out STD_LOGIC; 
  data_out_102 : out STD_LOGIC; 
  data_out_103 : out STD_LOGIC; 
  data_out_104 : out STD_LOGIC; 
  data_out_105 : out STD_LOGIC; 
  data_out_106 : out STD_LOGIC; 
  data_out_107 : out STD_LOGIC; 
  data_out_108 : out STD_LOGIC; 
  data_out_109 : out STD_LOGIC; 
  data_out_11 : out STD_LOGIC; 
  data_out_110 : out STD_LOGIC; 
  data_out_111 : out STD_LOGIC; 
  data_out_112 : out STD_LOGIC; 
  data_out_113 : out STD_LOGIC; 
  data_out_114 : out STD_LOGIC; 
  data_out_115 : out STD_LOGIC; 
  data_out_116 : out STD_LOGIC; 
  data_out_117 : out STD_LOGIC; 
  data_out_118 : out STD_LOGIC; 
  data_out_119 : out STD_LOGIC; 
  data_out_12 : out STD_LOGIC; 
  data_out_120 : out STD_LOGIC; 
  data_out_121 : out STD_LOGIC; 
  data_out_122 : out STD_LOGIC; 
  data_out_123 : out STD_LOGIC; 
  data_out_124 : out STD_LOGIC; 
  data_out_125 : out STD_LOGIC; 
  data_out_126 : out STD_LOGIC; 
  data_out_127 : out STD_LOGIC; 
  data_out_128 : out STD_LOGIC; 
  data_out_129 : out STD_LOGIC; 
  data_out_13 : out STD_LOGIC; 
  data_out_130 : out STD_LOGIC; 
  data_out_131 : out STD_LOGIC; 
  data_out_132 : out STD_LOGIC; 
  data_out_133 : out STD_LOGIC; 
  data_out_134 : out STD_LOGIC; 
  data_out_135 : out STD_LOGIC; 
  data_out_136 : out STD_LOGIC; 
  data_out_137 : out STD_LOGIC; 
  data_out_138 : out STD_LOGIC; 
  data_out_139 : out STD_LOGIC; 
  data_out_14 : out STD_LOGIC; 
  data_out_140 : out STD_LOGIC; 
  data_out_141 : out STD_LOGIC; 
  data_out_142 : out STD_LOGIC; 
  data_out_143 : out STD_LOGIC; 
  data_out_144 : out STD_LOGIC; 
  data_out_145 : out STD_LOGIC; 
  data_out_146 : out STD_LOGIC; 
  data_out_147 : out STD_LOGIC; 
  data_out_148 : out STD_LOGIC; 
  data_out_149 : out STD_LOGIC; 
  data_out_15 : out STD_LOGIC; 
  data_out_150 : out STD_LOGIC; 
  data_out_151 : out STD_LOGIC; 
  data_out_152 : out STD_LOGIC; 
  data_out_153 : out STD_LOGIC; 
  data_out_154 : out STD_LOGIC; 
  data_out_155 : out STD_LOGIC; 
  data_out_156 : out STD_LOGIC; 
  data_out_157 : out STD_LOGIC; 
  data_out_158 : out STD_LOGIC; 
  data_out_159 : out STD_LOGIC; 
  data_out_16 : out STD_LOGIC; 
  data_out_160 : out STD_LOGIC; 
  data_out_161 : out STD_LOGIC; 
  data_out_162 : out STD_LOGIC; 
  data_out_163 : out STD_LOGIC; 
  data_out_164 : out STD_LOGIC; 
  data_out_165 : out STD_LOGIC; 
  data_out_166 : out STD_LOGIC; 
  data_out_167 : out STD_LOGIC; 
  data_out_168 : out STD_LOGIC; 
  data_out_169 : out STD_LOGIC; 
  data_out_17 : out STD_LOGIC; 
  data_out_170 : out STD_LOGIC; 
  data_out_171 : out STD_LOGIC; 
  data_out_172 : out STD_LOGIC; 
  data_out_173 : out STD_LOGIC; 
  data_out_174 : out STD_LOGIC; 
  data_out_175 : out STD_LOGIC; 
  data_out_176 : out STD_LOGIC; 
  data_out_177 : out STD_LOGIC; 
  data_out_178 : out STD_LOGIC; 
  data_out_179 : out STD_LOGIC; 
  data_out_18 : out STD_LOGIC; 
  data_out_180 : out STD_LOGIC; 
  data_out_181 : out STD_LOGIC; 
  data_out_182 : out STD_LOGIC; 
  data_out_183 : out STD_LOGIC; 
  data_out_184 : out STD_LOGIC; 
  data_out_185 : out STD_LOGIC; 
  data_out_186 : out STD_LOGIC; 
  data_out_187 : out STD_LOGIC; 
  data_out_188 : out STD_LOGIC; 
  data_out_189 : out STD_LOGIC; 
  data_out_19 : out STD_LOGIC; 
  data_out_190 : out STD_LOGIC; 
  data_out_191 : out STD_LOGIC; 
  data_out_192 : out STD_LOGIC; 
  data_out_193 : out STD_LOGIC; 
  data_out_194 : out STD_LOGIC; 
  data_out_195 : out STD_LOGIC; 
  data_out_196 : out STD_LOGIC; 
  data_out_197 : out STD_LOGIC; 
  data_out_198 : out STD_LOGIC; 
  data_out_199 : out STD_LOGIC; 
  data_out_2 : out STD_LOGIC; 
  data_out_20 : out STD_LOGIC; 
  data_out_200 : out STD_LOGIC; 
  data_out_201 : out STD_LOGIC; 
  data_out_202 : out STD_LOGIC; 
  data_out_203 : out STD_LOGIC; 
  data_out_204 : out STD_LOGIC; 
  data_out_205 : out STD_LOGIC; 
  data_out_206 : out STD_LOGIC; 
  data_out_207 : out STD_LOGIC; 
  data_out_208 : out STD_LOGIC; 
  data_out_209 : out STD_LOGIC; 
  data_out_21 : out STD_LOGIC; 
  data_out_210 : out STD_LOGIC; 
  data_out_211 : out STD_LOGIC; 
  data_out_212 : out STD_LOGIC; 
  data_out_213 : out STD_LOGIC; 
  data_out_214 : out STD_LOGIC; 
  data_out_215 : out STD_LOGIC; 
  data_out_216 : out STD_LOGIC; 
  data_out_217 : out STD_LOGIC; 
  data_out_218 : out STD_LOGIC; 
  data_out_219 : out STD_LOGIC; 
  data_out_22 : out STD_LOGIC; 
  data_out_220 : out STD_LOGIC; 
  data_out_221 : out STD_LOGIC; 
  data_out_222 : out STD_LOGIC; 
  data_out_223 : out STD_LOGIC; 
  data_out_224 : out STD_LOGIC; 
  data_out_225 : out STD_LOGIC; 
  data_out_226 : out STD_LOGIC; 
  data_out_227 : out STD_LOGIC; 
  data_out_228 : out STD_LOGIC; 
  data_out_229 : out STD_LOGIC; 
  data_out_23 : out STD_LOGIC; 
  data_out_230 : out STD_LOGIC; 
  data_out_231 : out STD_LOGIC; 
  data_out_232 : out STD_LOGIC; 
  data_out_233 : out STD_LOGIC; 
  data_out_234 : out STD_LOGIC; 
  data_out_235 : out STD_LOGIC; 
  data_out_236 : out STD_LOGIC; 
  data_out_237 : out STD_LOGIC; 
  data_out_238 : out STD_LOGIC; 
  data_out_239 : out STD_LOGIC; 
  data_out_24 : out STD_LOGIC; 
  data_out_240 : out STD_LOGIC; 
  data_out_241 : out STD_LOGIC; 
  data_out_242 : out STD_LOGIC; 
  data_out_243 : out STD_LOGIC; 
  data_out_244 : out STD_LOGIC; 
  data_out_245 : out STD_LOGIC; 
  data_out_246 : out STD_LOGIC; 
  data_out_247 : out STD_LOGIC; 
  data_out_248 : out STD_LOGIC; 
  data_out_249 : out STD_LOGIC; 
  data_out_25 : out STD_LOGIC; 
  data_out_250 : out STD_LOGIC; 
  data_out_251 : out STD_LOGIC; 
  data_out_252 : out STD_LOGIC; 
  data_out_253 : out STD_LOGIC; 
  data_out_254 : out STD_LOGIC; 
  data_out_255 : out STD_LOGIC; 
  data_out_26 : out STD_LOGIC; 
  data_out_27 : out STD_LOGIC; 
  data_out_28 : out STD_LOGIC; 
  data_out_29 : out STD_LOGIC; 
  data_out_3 : out STD_LOGIC; 
  data_out_30 : out STD_LOGIC; 
  data_out_31 : out STD_LOGIC; 
  data_out_32 : out STD_LOGIC; 
  data_out_33 : out STD_LOGIC; 
  data_out_34 : out STD_LOGIC; 
  data_out_35 : out STD_LOGIC; 
  data_out_36 : out STD_LOGIC; 
  data_out_37 : out STD_LOGIC; 
  data_out_38 : out STD_LOGIC; 
  data_out_39 : out STD_LOGIC; 
  data_out_4 : out STD_LOGIC; 
  data_out_40 : out STD_LOGIC; 
  data_out_41 : out STD_LOGIC; 
  data_out_42 : out STD_LOGIC; 
  data_out_43 : out STD_LOGIC; 
  data_out_44 : out STD_LOGIC; 
  data_out_45 : out STD_LOGIC; 
  data_out_46 : out STD_LOGIC; 
  data_out_47 : out STD_LOGIC; 
  data_out_48 : out STD_LOGIC; 
  data_out_49 : out STD_LOGIC; 
  data_out_5 : out STD_LOGIC; 
  data_out_50 : out STD_LOGIC; 
  data_out_51 : out STD_LOGIC; 
  data_out_52 : out STD_LOGIC; 
  data_out_53 : out STD_LOGIC; 
  data_out_54 : out STD_LOGIC; 
  data_out_55 : out STD_LOGIC; 
  data_out_56 : out STD_LOGIC; 
  data_out_57 : out STD_LOGIC; 
  data_out_58 : out STD_LOGIC; 
  data_out_59 : out STD_LOGIC; 
  data_out_6 : out STD_LOGIC; 
  data_out_60 : out STD_LOGIC; 
  data_out_61 : out STD_LOGIC; 
  data_out_62 : out STD_LOGIC; 
  data_out_63 : out STD_LOGIC; 
  data_out_64 : out STD_LOGIC; 
  data_out_65 : out STD_LOGIC; 
  data_out_66 : out STD_LOGIC; 
  data_out_67 : out STD_LOGIC; 
  data_out_68 : out STD_LOGIC; 
  data_out_69 : out STD_LOGIC; 
  data_out_7 : out STD_LOGIC; 
  data_out_70 : out STD_LOGIC; 
  data_out_71 : out STD_LOGIC; 
  data_out_72 : out STD_LOGIC; 
  data_out_73 : out STD_LOGIC; 
  data_out_74 : out STD_LOGIC; 
  data_out_75 : out STD_LOGIC; 
  data_out_76 : out STD_LOGIC; 
  data_out_77 : out STD_LOGIC; 
  data_out_78 : out STD_LOGIC; 
  data_out_79 : out STD_LOGIC; 
  data_out_8 : out STD_LOGIC; 
  data_out_80 : out STD_LOGIC; 
  data_out_81 : out STD_LOGIC; 
  data_out_82 : out STD_LOGIC; 
  data_out_83 : out STD_LOGIC; 
  data_out_84 : out STD_LOGIC; 
  data_out_85 : out STD_LOGIC; 
  data_out_86 : out STD_LOGIC; 
  data_out_87 : out STD_LOGIC; 
  data_out_88 : out STD_LOGIC; 
  data_out_89 : out STD_LOGIC; 
  data_out_9 : out STD_LOGIC; 
  data_out_90 : out STD_LOGIC; 
  data_out_91 : out STD_LOGIC; 
  data_out_92 : out STD_LOGIC; 
  data_out_93 : out STD_LOGIC; 
  data_out_94 : out STD_LOGIC; 
  data_out_95 : out STD_LOGIC; 
  data_out_96 : out STD_LOGIC; 
  data_out_97 : out STD_LOGIC; 
  data_out_98 : out STD_LOGIC; 
  data_out_99 : out STD_LOGIC; 
  finished : out STD_LOGIC
);
end sha_256_core;

architecture STRUCTURE of sha_256_core is
  signal a_0_i_1_n_0 : STD_LOGIC;
  signal a_10_i_1_n_0 : STD_LOGIC;
  signal a_11_i_1_n_0 : STD_LOGIC;
  signal a_11_i_3_n_0 : STD_LOGIC;
  signal a_11_i_4_n_0 : STD_LOGIC;
  signal a_11_i_5_n_0 : STD_LOGIC;
  signal a_11_i_6_n_0 : STD_LOGIC;
  signal a_12_i_1_n_0 : STD_LOGIC;
  signal a_13_i_1_n_0 : STD_LOGIC;
  signal a_14_i_1_n_0 : STD_LOGIC;
  signal a_15_i_1_n_0 : STD_LOGIC;
  signal a_15_i_3_n_0 : STD_LOGIC;
  signal a_15_i_4_n_0 : STD_LOGIC;
  signal a_15_i_5_n_0 : STD_LOGIC;
  signal a_15_i_6_n_0 : STD_LOGIC;
  signal a_16_i_1_n_0 : STD_LOGIC;
  signal a_17_i_1_n_0 : STD_LOGIC;
  signal a_18_i_1_n_0 : STD_LOGIC;
  signal a_19_i_1_n_0 : STD_LOGIC;
  signal a_19_i_3_n_0 : STD_LOGIC;
  signal a_19_i_4_n_0 : STD_LOGIC;
  signal a_19_i_5_n_0 : STD_LOGIC;
  signal a_19_i_6_n_0 : STD_LOGIC;
  signal a_1_i_1_n_0 : STD_LOGIC;
  signal a_20_i_1_n_0 : STD_LOGIC;
  signal a_21_i_1_n_0 : STD_LOGIC;
  signal a_22_i_1_n_0 : STD_LOGIC;
  signal a_23_i_1_n_0 : STD_LOGIC;
  signal a_23_i_3_n_0 : STD_LOGIC;
  signal a_23_i_4_n_0 : STD_LOGIC;
  signal a_23_i_5_n_0 : STD_LOGIC;
  signal a_23_i_6_n_0 : STD_LOGIC;
  signal a_24_i_1_n_0 : STD_LOGIC;
  signal a_25_i_1_n_0 : STD_LOGIC;
  signal a_26_i_1_n_0 : STD_LOGIC;
  signal a_27_i_1_n_0 : STD_LOGIC;
  signal a_27_i_3_n_0 : STD_LOGIC;
  signal a_27_i_4_n_0 : STD_LOGIC;
  signal a_27_i_5_n_0 : STD_LOGIC;
  signal a_27_i_6_n_0 : STD_LOGIC;
  signal a_28_i_1_n_0 : STD_LOGIC;
  signal a_29_i_1_n_0 : STD_LOGIC;
  signal a_2_i_1_n_0 : STD_LOGIC;
  signal a_30_i_1_n_0 : STD_LOGIC;
  signal a_31_i_1_n_0 : STD_LOGIC;
  signal a_31_i_2_n_0 : STD_LOGIC;
  signal a_31_i_4_n_0 : STD_LOGIC;
  signal a_31_i_5_n_0 : STD_LOGIC;
  signal a_31_i_6_n_0 : STD_LOGIC;
  signal a_31_i_7_n_0 : STD_LOGIC;
  signal a_3_i_1_n_0 : STD_LOGIC;
  signal a_3_i_3_n_0 : STD_LOGIC;
  signal a_3_i_4_n_0 : STD_LOGIC;
  signal a_3_i_5_n_0 : STD_LOGIC;
  signal a_3_i_6_n_0 : STD_LOGIC;
  signal a_4_i_1_n_0 : STD_LOGIC;
  signal a_5_i_1_n_0 : STD_LOGIC;
  signal a_6_i_1_n_0 : STD_LOGIC;
  signal a_7_i_1_n_0 : STD_LOGIC;
  signal a_7_i_3_n_0 : STD_LOGIC;
  signal a_7_i_4_n_0 : STD_LOGIC;
  signal a_7_i_5_n_0 : STD_LOGIC;
  signal a_7_i_6_n_0 : STD_LOGIC;
  signal a_8_i_1_n_0 : STD_LOGIC;
  signal a_9_i_1_n_0 : STD_LOGIC;
  signal a_reg_11_i_2_n_0 : STD_LOGIC;
  signal a_reg_11_i_2_n_1 : STD_LOGIC;
  signal a_reg_11_i_2_n_2 : STD_LOGIC;
  signal a_reg_11_i_2_n_3 : STD_LOGIC;
  signal a_reg_15_i_2_n_0 : STD_LOGIC;
  signal a_reg_15_i_2_n_1 : STD_LOGIC;
  signal a_reg_15_i_2_n_2 : STD_LOGIC;
  signal a_reg_15_i_2_n_3 : STD_LOGIC;
  signal a_reg_19_i_2_n_0 : STD_LOGIC;
  signal a_reg_19_i_2_n_1 : STD_LOGIC;
  signal a_reg_19_i_2_n_2 : STD_LOGIC;
  signal a_reg_19_i_2_n_3 : STD_LOGIC;
  signal a_reg_23_i_2_n_0 : STD_LOGIC;
  signal a_reg_23_i_2_n_1 : STD_LOGIC;
  signal a_reg_23_i_2_n_2 : STD_LOGIC;
  signal a_reg_23_i_2_n_3 : STD_LOGIC;
  signal a_reg_27_i_2_n_0 : STD_LOGIC;
  signal a_reg_27_i_2_n_1 : STD_LOGIC;
  signal a_reg_27_i_2_n_2 : STD_LOGIC;
  signal a_reg_27_i_2_n_3 : STD_LOGIC;
  signal a_reg_31_i_3_n_1 : STD_LOGIC;
  signal a_reg_31_i_3_n_2 : STD_LOGIC;
  signal a_reg_31_i_3_n_3 : STD_LOGIC;
  signal a_reg_3_i_2_n_0 : STD_LOGIC;
  signal a_reg_3_i_2_n_1 : STD_LOGIC;
  signal a_reg_3_i_2_n_2 : STD_LOGIC;
  signal a_reg_3_i_2_n_3 : STD_LOGIC;
  signal a_reg_7_i_2_n_0 : STD_LOGIC;
  signal a_reg_7_i_2_n_1 : STD_LOGIC;
  signal a_reg_7_i_2_n_2 : STD_LOGIC;
  signal a_reg_7_i_2_n_3 : STD_LOGIC;
  signal b_0_i_1_n_0 : STD_LOGIC;
  signal b_10_i_1_n_0 : STD_LOGIC;
  signal b_11_i_1_n_0 : STD_LOGIC;
  signal b_12_i_1_n_0 : STD_LOGIC;
  signal b_13_i_1_n_0 : STD_LOGIC;
  signal b_14_i_1_n_0 : STD_LOGIC;
  signal b_15_i_1_n_0 : STD_LOGIC;
  signal b_16_i_1_n_0 : STD_LOGIC;
  signal b_17_i_1_n_0 : STD_LOGIC;
  signal b_18_i_1_n_0 : STD_LOGIC;
  signal b_19_i_1_n_0 : STD_LOGIC;
  signal b_1_i_1_n_0 : STD_LOGIC;
  signal b_20_i_1_n_0 : STD_LOGIC;
  signal b_21_i_1_n_0 : STD_LOGIC;
  signal b_22_i_1_n_0 : STD_LOGIC;
  signal b_23_i_1_n_0 : STD_LOGIC;
  signal b_24_i_1_n_0 : STD_LOGIC;
  signal b_25_i_1_n_0 : STD_LOGIC;
  signal b_26_i_1_n_0 : STD_LOGIC;
  signal b_27_i_1_n_0 : STD_LOGIC;
  signal b_28_i_1_n_0 : STD_LOGIC;
  signal b_29_i_1_n_0 : STD_LOGIC;
  signal b_2_i_1_n_0 : STD_LOGIC;
  signal b_30_i_1_n_0 : STD_LOGIC;
  signal b_31_i_1_n_0 : STD_LOGIC;
  signal b_3_i_1_n_0 : STD_LOGIC;
  signal b_4_i_1_n_0 : STD_LOGIC;
  signal b_5_i_1_n_0 : STD_LOGIC;
  signal b_6_i_1_n_0 : STD_LOGIC;
  signal b_7_i_1_n_0 : STD_LOGIC;
  signal b_8_i_1_n_0 : STD_LOGIC;
  signal b_9_i_1_n_0 : STD_LOGIC;
  signal b_reg_n_0_0 : STD_LOGIC;
  signal b_reg_n_0_10 : STD_LOGIC;
  signal b_reg_n_0_11 : STD_LOGIC;
  signal b_reg_n_0_12 : STD_LOGIC;
  signal b_reg_n_0_13 : STD_LOGIC;
  signal b_reg_n_0_14 : STD_LOGIC;
  signal b_reg_n_0_15 : STD_LOGIC;
  signal b_reg_n_0_16 : STD_LOGIC;
  signal b_reg_n_0_17 : STD_LOGIC;
  signal b_reg_n_0_18 : STD_LOGIC;
  signal b_reg_n_0_19 : STD_LOGIC;
  signal b_reg_n_0_1 : STD_LOGIC;
  signal b_reg_n_0_20 : STD_LOGIC;
  signal b_reg_n_0_21 : STD_LOGIC;
  signal b_reg_n_0_22 : STD_LOGIC;
  signal b_reg_n_0_23 : STD_LOGIC;
  signal b_reg_n_0_24 : STD_LOGIC;
  signal b_reg_n_0_25 : STD_LOGIC;
  signal b_reg_n_0_26 : STD_LOGIC;
  signal b_reg_n_0_27 : STD_LOGIC;
  signal b_reg_n_0_28 : STD_LOGIC;
  signal b_reg_n_0_29 : STD_LOGIC;
  signal b_reg_n_0_2 : STD_LOGIC;
  signal b_reg_n_0_30 : STD_LOGIC;
  signal b_reg_n_0_31 : STD_LOGIC;
  signal b_reg_n_0_3 : STD_LOGIC;
  signal b_reg_n_0_4 : STD_LOGIC;
  signal b_reg_n_0_5 : STD_LOGIC;
  signal b_reg_n_0_6 : STD_LOGIC;
  signal b_reg_n_0_7 : STD_LOGIC;
  signal b_reg_n_0_8 : STD_LOGIC;
  signal b_reg_n_0_9 : STD_LOGIC;
  signal clk_IBUF : STD_LOGIC;
  signal clk_IBUF_BUFG : STD_LOGIC;
  signal c_0_i_1_n_0 : STD_LOGIC;
  signal c_10_i_1_n_0 : STD_LOGIC;
  signal c_11_i_1_n_0 : STD_LOGIC;
  signal c_12_i_1_n_0 : STD_LOGIC;
  signal c_13_i_1_n_0 : STD_LOGIC;
  signal c_14_i_1_n_0 : STD_LOGIC;
  signal c_15_i_1_n_0 : STD_LOGIC;
  signal c_16_i_1_n_0 : STD_LOGIC;
  signal c_17_i_1_n_0 : STD_LOGIC;
  signal c_18_i_1_n_0 : STD_LOGIC;
  signal c_19_i_1_n_0 : STD_LOGIC;
  signal c_1_i_1_n_0 : STD_LOGIC;
  signal c_20_i_1_n_0 : STD_LOGIC;
  signal c_21_i_1_n_0 : STD_LOGIC;
  signal c_22_i_1_n_0 : STD_LOGIC;
  signal c_23_i_1_n_0 : STD_LOGIC;
  signal c_24_i_1_n_0 : STD_LOGIC;
  signal c_25_i_1_n_0 : STD_LOGIC;
  signal c_26_i_1_n_0 : STD_LOGIC;
  signal c_27_i_1_n_0 : STD_LOGIC;
  signal c_28_i_1_n_0 : STD_LOGIC;
  signal c_29_i_1_n_0 : STD_LOGIC;
  signal c_2_i_1_n_0 : STD_LOGIC;
  signal c_30_i_1_n_0 : STD_LOGIC;
  signal c_31_i_1_n_0 : STD_LOGIC;
  signal c_3_i_1_n_0 : STD_LOGIC;
  signal c_4_i_1_n_0 : STD_LOGIC;
  signal c_5_i_1_n_0 : STD_LOGIC;
  signal c_6_i_1_n_0 : STD_LOGIC;
  signal c_7_i_1_n_0 : STD_LOGIC;
  signal c_8_i_1_n_0 : STD_LOGIC;
  signal c_9_i_1_n_0 : STD_LOGIC;
  signal c_reg_n_0_0 : STD_LOGIC;
  signal c_reg_n_0_10 : STD_LOGIC;
  signal c_reg_n_0_11 : STD_LOGIC;
  signal c_reg_n_0_12 : STD_LOGIC;
  signal c_reg_n_0_13 : STD_LOGIC;
  signal c_reg_n_0_14 : STD_LOGIC;
  signal c_reg_n_0_15 : STD_LOGIC;
  signal c_reg_n_0_16 : STD_LOGIC;
  signal c_reg_n_0_17 : STD_LOGIC;
  signal c_reg_n_0_18 : STD_LOGIC;
  signal c_reg_n_0_19 : STD_LOGIC;
  signal c_reg_n_0_1 : STD_LOGIC;
  signal c_reg_n_0_20 : STD_LOGIC;
  signal c_reg_n_0_21 : STD_LOGIC;
  signal c_reg_n_0_22 : STD_LOGIC;
  signal c_reg_n_0_23 : STD_LOGIC;
  signal c_reg_n_0_24 : STD_LOGIC;
  signal c_reg_n_0_25 : STD_LOGIC;
  signal c_reg_n_0_26 : STD_LOGIC;
  signal c_reg_n_0_27 : STD_LOGIC;
  signal c_reg_n_0_28 : STD_LOGIC;
  signal c_reg_n_0_29 : STD_LOGIC;
  signal c_reg_n_0_2 : STD_LOGIC;
  signal c_reg_n_0_30 : STD_LOGIC;
  signal c_reg_n_0_31 : STD_LOGIC;
  signal c_reg_n_0_3 : STD_LOGIC;
  signal c_reg_n_0_4 : STD_LOGIC;
  signal c_reg_n_0_5 : STD_LOGIC;
  signal c_reg_n_0_6 : STD_LOGIC;
  signal c_reg_n_0_7 : STD_LOGIC;
  signal c_reg_n_0_8 : STD_LOGIC;
  signal c_reg_n_0_9 : STD_LOGIC;
  signal d_31 : STD_LOGIC;
  signal d_30 : STD_LOGIC;
  signal d_29 : STD_LOGIC;
  signal d_28 : STD_LOGIC;
  signal d_27 : STD_LOGIC;
  signal d_26 : STD_LOGIC;
  signal d_25 : STD_LOGIC;
  signal d_24 : STD_LOGIC;
  signal d_23 : STD_LOGIC;
  signal d_22 : STD_LOGIC;
  signal d_21 : STD_LOGIC;
  signal d_20 : STD_LOGIC;
  signal d_19 : STD_LOGIC;
  signal d_18 : STD_LOGIC;
  signal d_17 : STD_LOGIC;
  signal d_16 : STD_LOGIC;
  signal d_15 : STD_LOGIC;
  signal d_14 : STD_LOGIC;
  signal d_13 : STD_LOGIC;
  signal d_12 : STD_LOGIC;
  signal d_11 : STD_LOGIC;
  signal d_10 : STD_LOGIC;
  signal d_9 : STD_LOGIC;
  signal d_8 : STD_LOGIC;
  signal d_7 : STD_LOGIC;
  signal d_6 : STD_LOGIC;
  signal d_5 : STD_LOGIC;
  signal d_4 : STD_LOGIC;
  signal d_3 : STD_LOGIC;
  signal d_2 : STD_LOGIC;
  signal d_1 : STD_LOGIC;
  signal d_0 : STD_LOGIC;
  signal data_out_OBUF_255 : STD_LOGIC;
  signal data_out_OBUF_254 : STD_LOGIC;
  signal data_out_OBUF_253 : STD_LOGIC;
  signal data_out_OBUF_252 : STD_LOGIC;
  signal data_out_OBUF_251 : STD_LOGIC;
  signal data_out_OBUF_250 : STD_LOGIC;
  signal data_out_OBUF_249 : STD_LOGIC;
  signal data_out_OBUF_248 : STD_LOGIC;
  signal data_out_OBUF_247 : STD_LOGIC;
  signal data_out_OBUF_246 : STD_LOGIC;
  signal data_out_OBUF_245 : STD_LOGIC;
  signal data_out_OBUF_244 : STD_LOGIC;
  signal data_out_OBUF_243 : STD_LOGIC;
  signal data_out_OBUF_242 : STD_LOGIC;
  signal data_out_OBUF_241 : STD_LOGIC;
  signal data_out_OBUF_240 : STD_LOGIC;
  signal data_out_OBUF_239 : STD_LOGIC;
  signal data_out_OBUF_238 : STD_LOGIC;
  signal data_out_OBUF_237 : STD_LOGIC;
  signal data_out_OBUF_236 : STD_LOGIC;
  signal data_out_OBUF_235 : STD_LOGIC;
  signal data_out_OBUF_234 : STD_LOGIC;
  signal data_out_OBUF_233 : STD_LOGIC;
  signal data_out_OBUF_232 : STD_LOGIC;
  signal data_out_OBUF_231 : STD_LOGIC;
  signal data_out_OBUF_230 : STD_LOGIC;
  signal data_out_OBUF_229 : STD_LOGIC;
  signal data_out_OBUF_228 : STD_LOGIC;
  signal data_out_OBUF_227 : STD_LOGIC;
  signal data_out_OBUF_226 : STD_LOGIC;
  signal data_out_OBUF_225 : STD_LOGIC;
  signal data_out_OBUF_224 : STD_LOGIC;
  signal data_out_OBUF_223 : STD_LOGIC;
  signal data_out_OBUF_222 : STD_LOGIC;
  signal data_out_OBUF_221 : STD_LOGIC;
  signal data_out_OBUF_220 : STD_LOGIC;
  signal data_out_OBUF_219 : STD_LOGIC;
  signal data_out_OBUF_218 : STD_LOGIC;
  signal data_out_OBUF_217 : STD_LOGIC;
  signal data_out_OBUF_216 : STD_LOGIC;
  signal data_out_OBUF_215 : STD_LOGIC;
  signal data_out_OBUF_214 : STD_LOGIC;
  signal data_out_OBUF_213 : STD_LOGIC;
  signal data_out_OBUF_212 : STD_LOGIC;
  signal data_out_OBUF_211 : STD_LOGIC;
  signal data_out_OBUF_210 : STD_LOGIC;
  signal data_out_OBUF_209 : STD_LOGIC;
  signal data_out_OBUF_208 : STD_LOGIC;
  signal data_out_OBUF_207 : STD_LOGIC;
  signal data_out_OBUF_206 : STD_LOGIC;
  signal data_out_OBUF_205 : STD_LOGIC;
  signal data_out_OBUF_204 : STD_LOGIC;
  signal data_out_OBUF_203 : STD_LOGIC;
  signal data_out_OBUF_202 : STD_LOGIC;
  signal data_out_OBUF_201 : STD_LOGIC;
  signal data_out_OBUF_200 : STD_LOGIC;
  signal data_out_OBUF_199 : STD_LOGIC;
  signal data_out_OBUF_198 : STD_LOGIC;
  signal data_out_OBUF_197 : STD_LOGIC;
  signal data_out_OBUF_196 : STD_LOGIC;
  signal data_out_OBUF_195 : STD_LOGIC;
  signal data_out_OBUF_194 : STD_LOGIC;
  signal data_out_OBUF_193 : STD_LOGIC;
  signal data_out_OBUF_192 : STD_LOGIC;
  signal data_out_OBUF_191 : STD_LOGIC;
  signal data_out_OBUF_190 : STD_LOGIC;
  signal data_out_OBUF_189 : STD_LOGIC;
  signal data_out_OBUF_188 : STD_LOGIC;
  signal data_out_OBUF_187 : STD_LOGIC;
  signal data_out_OBUF_186 : STD_LOGIC;
  signal data_out_OBUF_185 : STD_LOGIC;
  signal data_out_OBUF_184 : STD_LOGIC;
  signal data_out_OBUF_183 : STD_LOGIC;
  signal data_out_OBUF_182 : STD_LOGIC;
  signal data_out_OBUF_181 : STD_LOGIC;
  signal data_out_OBUF_180 : STD_LOGIC;
  signal data_out_OBUF_179 : STD_LOGIC;
  signal data_out_OBUF_178 : STD_LOGIC;
  signal data_out_OBUF_177 : STD_LOGIC;
  signal data_out_OBUF_176 : STD_LOGIC;
  signal data_out_OBUF_175 : STD_LOGIC;
  signal data_out_OBUF_174 : STD_LOGIC;
  signal data_out_OBUF_173 : STD_LOGIC;
  signal data_out_OBUF_172 : STD_LOGIC;
  signal data_out_OBUF_171 : STD_LOGIC;
  signal data_out_OBUF_170 : STD_LOGIC;
  signal data_out_OBUF_169 : STD_LOGIC;
  signal data_out_OBUF_168 : STD_LOGIC;
  signal data_out_OBUF_167 : STD_LOGIC;
  signal data_out_OBUF_166 : STD_LOGIC;
  signal data_out_OBUF_165 : STD_LOGIC;
  signal data_out_OBUF_164 : STD_LOGIC;
  signal data_out_OBUF_163 : STD_LOGIC;
  signal data_out_OBUF_162 : STD_LOGIC;
  signal data_out_OBUF_161 : STD_LOGIC;
  signal data_out_OBUF_160 : STD_LOGIC;
  signal data_out_OBUF_159 : STD_LOGIC;
  signal data_out_OBUF_158 : STD_LOGIC;
  signal data_out_OBUF_157 : STD_LOGIC;
  signal data_out_OBUF_156 : STD_LOGIC;
  signal data_out_OBUF_155 : STD_LOGIC;
  signal data_out_OBUF_154 : STD_LOGIC;
  signal data_out_OBUF_153 : STD_LOGIC;
  signal data_out_OBUF_152 : STD_LOGIC;
  signal data_out_OBUF_151 : STD_LOGIC;
  signal data_out_OBUF_150 : STD_LOGIC;
  signal data_out_OBUF_149 : STD_LOGIC;
  signal data_out_OBUF_148 : STD_LOGIC;
  signal data_out_OBUF_147 : STD_LOGIC;
  signal data_out_OBUF_146 : STD_LOGIC;
  signal data_out_OBUF_145 : STD_LOGIC;
  signal data_out_OBUF_144 : STD_LOGIC;
  signal data_out_OBUF_143 : STD_LOGIC;
  signal data_out_OBUF_142 : STD_LOGIC;
  signal data_out_OBUF_141 : STD_LOGIC;
  signal data_out_OBUF_140 : STD_LOGIC;
  signal data_out_OBUF_139 : STD_LOGIC;
  signal data_out_OBUF_138 : STD_LOGIC;
  signal data_out_OBUF_137 : STD_LOGIC;
  signal data_out_OBUF_136 : STD_LOGIC;
  signal data_out_OBUF_135 : STD_LOGIC;
  signal data_out_OBUF_134 : STD_LOGIC;
  signal data_out_OBUF_133 : STD_LOGIC;
  signal data_out_OBUF_132 : STD_LOGIC;
  signal data_out_OBUF_131 : STD_LOGIC;
  signal data_out_OBUF_130 : STD_LOGIC;
  signal data_out_OBUF_129 : STD_LOGIC;
  signal data_out_OBUF_128 : STD_LOGIC;
  signal data_out_OBUF_127 : STD_LOGIC;
  signal data_out_OBUF_126 : STD_LOGIC;
  signal data_out_OBUF_125 : STD_LOGIC;
  signal data_out_OBUF_124 : STD_LOGIC;
  signal data_out_OBUF_123 : STD_LOGIC;
  signal data_out_OBUF_122 : STD_LOGIC;
  signal data_out_OBUF_121 : STD_LOGIC;
  signal data_out_OBUF_120 : STD_LOGIC;
  signal data_out_OBUF_119 : STD_LOGIC;
  signal data_out_OBUF_118 : STD_LOGIC;
  signal data_out_OBUF_117 : STD_LOGIC;
  signal data_out_OBUF_116 : STD_LOGIC;
  signal data_out_OBUF_115 : STD_LOGIC;
  signal data_out_OBUF_114 : STD_LOGIC;
  signal data_out_OBUF_113 : STD_LOGIC;
  signal data_out_OBUF_112 : STD_LOGIC;
  signal data_out_OBUF_111 : STD_LOGIC;
  signal data_out_OBUF_110 : STD_LOGIC;
  signal data_out_OBUF_109 : STD_LOGIC;
  signal data_out_OBUF_108 : STD_LOGIC;
  signal data_out_OBUF_107 : STD_LOGIC;
  signal data_out_OBUF_106 : STD_LOGIC;
  signal data_out_OBUF_105 : STD_LOGIC;
  signal data_out_OBUF_104 : STD_LOGIC;
  signal data_out_OBUF_103 : STD_LOGIC;
  signal data_out_OBUF_102 : STD_LOGIC;
  signal data_out_OBUF_101 : STD_LOGIC;
  signal data_out_OBUF_100 : STD_LOGIC;
  signal data_out_OBUF_99 : STD_LOGIC;
  signal data_out_OBUF_98 : STD_LOGIC;
  signal data_out_OBUF_97 : STD_LOGIC;
  signal data_out_OBUF_96 : STD_LOGIC;
  signal data_out_OBUF_95 : STD_LOGIC;
  signal data_out_OBUF_94 : STD_LOGIC;
  signal data_out_OBUF_93 : STD_LOGIC;
  signal data_out_OBUF_92 : STD_LOGIC;
  signal data_out_OBUF_91 : STD_LOGIC;
  signal data_out_OBUF_90 : STD_LOGIC;
  signal data_out_OBUF_89 : STD_LOGIC;
  signal data_out_OBUF_88 : STD_LOGIC;
  signal data_out_OBUF_87 : STD_LOGIC;
  signal data_out_OBUF_86 : STD_LOGIC;
  signal data_out_OBUF_85 : STD_LOGIC;
  signal data_out_OBUF_84 : STD_LOGIC;
  signal data_out_OBUF_83 : STD_LOGIC;
  signal data_out_OBUF_82 : STD_LOGIC;
  signal data_out_OBUF_81 : STD_LOGIC;
  signal data_out_OBUF_80 : STD_LOGIC;
  signal data_out_OBUF_79 : STD_LOGIC;
  signal data_out_OBUF_78 : STD_LOGIC;
  signal data_out_OBUF_77 : STD_LOGIC;
  signal data_out_OBUF_76 : STD_LOGIC;
  signal data_out_OBUF_75 : STD_LOGIC;
  signal data_out_OBUF_74 : STD_LOGIC;
  signal data_out_OBUF_73 : STD_LOGIC;
  signal data_out_OBUF_72 : STD_LOGIC;
  signal data_out_OBUF_71 : STD_LOGIC;
  signal data_out_OBUF_70 : STD_LOGIC;
  signal data_out_OBUF_69 : STD_LOGIC;
  signal data_out_OBUF_68 : STD_LOGIC;
  signal data_out_OBUF_67 : STD_LOGIC;
  signal data_out_OBUF_66 : STD_LOGIC;
  signal data_out_OBUF_65 : STD_LOGIC;
  signal data_out_OBUF_64 : STD_LOGIC;
  signal data_out_OBUF_63 : STD_LOGIC;
  signal data_out_OBUF_62 : STD_LOGIC;
  signal data_out_OBUF_61 : STD_LOGIC;
  signal data_out_OBUF_60 : STD_LOGIC;
  signal data_out_OBUF_59 : STD_LOGIC;
  signal data_out_OBUF_58 : STD_LOGIC;
  signal data_out_OBUF_57 : STD_LOGIC;
  signal data_out_OBUF_56 : STD_LOGIC;
  signal data_out_OBUF_55 : STD_LOGIC;
  signal data_out_OBUF_54 : STD_LOGIC;
  signal data_out_OBUF_53 : STD_LOGIC;
  signal data_out_OBUF_52 : STD_LOGIC;
  signal data_out_OBUF_51 : STD_LOGIC;
  signal data_out_OBUF_50 : STD_LOGIC;
  signal data_out_OBUF_49 : STD_LOGIC;
  signal data_out_OBUF_48 : STD_LOGIC;
  signal data_out_OBUF_47 : STD_LOGIC;
  signal data_out_OBUF_46 : STD_LOGIC;
  signal data_out_OBUF_45 : STD_LOGIC;
  signal data_out_OBUF_44 : STD_LOGIC;
  signal data_out_OBUF_43 : STD_LOGIC;
  signal data_out_OBUF_42 : STD_LOGIC;
  signal data_out_OBUF_41 : STD_LOGIC;
  signal data_out_OBUF_40 : STD_LOGIC;
  signal data_out_OBUF_39 : STD_LOGIC;
  signal data_out_OBUF_38 : STD_LOGIC;
  signal data_out_OBUF_37 : STD_LOGIC;
  signal data_out_OBUF_36 : STD_LOGIC;
  signal data_out_OBUF_35 : STD_LOGIC;
  signal data_out_OBUF_34 : STD_LOGIC;
  signal data_out_OBUF_33 : STD_LOGIC;
  signal data_out_OBUF_32 : STD_LOGIC;
  signal data_out_OBUF_31 : STD_LOGIC;
  signal data_out_OBUF_30 : STD_LOGIC;
  signal data_out_OBUF_29 : STD_LOGIC;
  signal data_out_OBUF_28 : STD_LOGIC;
  signal data_out_OBUF_27 : STD_LOGIC;
  signal data_out_OBUF_26 : STD_LOGIC;
  signal data_out_OBUF_25 : STD_LOGIC;
  signal data_out_OBUF_24 : STD_LOGIC;
  signal data_out_OBUF_23 : STD_LOGIC;
  signal data_out_OBUF_22 : STD_LOGIC;
  signal data_out_OBUF_21 : STD_LOGIC;
  signal data_out_OBUF_20 : STD_LOGIC;
  signal data_out_OBUF_19 : STD_LOGIC;
  signal data_out_OBUF_18 : STD_LOGIC;
  signal data_out_OBUF_17 : STD_LOGIC;
  signal data_out_OBUF_16 : STD_LOGIC;
  signal data_out_OBUF_15 : STD_LOGIC;
  signal data_out_OBUF_14 : STD_LOGIC;
  signal data_out_OBUF_13 : STD_LOGIC;
  signal data_out_OBUF_12 : STD_LOGIC;
  signal data_out_OBUF_11 : STD_LOGIC;
  signal data_out_OBUF_10 : STD_LOGIC;
  signal data_out_OBUF_9 : STD_LOGIC;
  signal data_out_OBUF_8 : STD_LOGIC;
  signal data_out_OBUF_7 : STD_LOGIC;
  signal data_out_OBUF_6 : STD_LOGIC;
  signal data_out_OBUF_5 : STD_LOGIC;
  signal data_out_OBUF_4 : STD_LOGIC;
  signal data_out_OBUF_3 : STD_LOGIC;
  signal data_out_OBUF_2 : STD_LOGIC;
  signal data_out_OBUF_1 : STD_LOGIC;
  signal data_out_OBUF_0 : STD_LOGIC;
  signal data_ready_IBUF : STD_LOGIC;
  signal d_0_i_1_n_0 : STD_LOGIC;
  signal d_10_i_1_n_0 : STD_LOGIC;
  signal d_11_i_1_n_0 : STD_LOGIC;
  signal d_12_i_1_n_0 : STD_LOGIC;
  signal d_13_i_1_n_0 : STD_LOGIC;
  signal d_14_i_1_n_0 : STD_LOGIC;
  signal d_15_i_1_n_0 : STD_LOGIC;
  signal d_16_i_1_n_0 : STD_LOGIC;
  signal d_17_i_1_n_0 : STD_LOGIC;
  signal d_18_i_1_n_0 : STD_LOGIC;
  signal d_19_i_1_n_0 : STD_LOGIC;
  signal d_1_i_1_n_0 : STD_LOGIC;
  signal d_20_i_1_n_0 : STD_LOGIC;
  signal d_21_i_1_n_0 : STD_LOGIC;
  signal d_22_i_1_n_0 : STD_LOGIC;
  signal d_23_i_1_n_0 : STD_LOGIC;
  signal d_24_i_1_n_0 : STD_LOGIC;
  signal d_25_i_1_n_0 : STD_LOGIC;
  signal d_26_i_1_n_0 : STD_LOGIC;
  signal d_27_i_1_n_0 : STD_LOGIC;
  signal d_28_i_1_n_0 : STD_LOGIC;
  signal d_29_i_1_n_0 : STD_LOGIC;
  signal d_2_i_1_n_0 : STD_LOGIC;
  signal d_30_i_1_n_0 : STD_LOGIC;
  signal d_31_i_1_n_0 : STD_LOGIC;
  signal d_3_i_1_n_0 : STD_LOGIC;
  signal d_4_i_1_n_0 : STD_LOGIC;
  signal d_5_i_1_n_0 : STD_LOGIC;
  signal d_6_i_1_n_0 : STD_LOGIC;
  signal d_7_i_1_n_0 : STD_LOGIC;
  signal d_8_i_1_n_0 : STD_LOGIC;
  signal d_9_i_1_n_0 : STD_LOGIC;
  signal e_0_i_1_n_0 : STD_LOGIC;
  signal e_10_i_1_n_0 : STD_LOGIC;
  signal e_11_i_1_n_0 : STD_LOGIC;
  signal e_11_i_3_n_0 : STD_LOGIC;
  signal e_11_i_4_n_0 : STD_LOGIC;
  signal e_11_i_5_n_0 : STD_LOGIC;
  signal e_11_i_6_n_0 : STD_LOGIC;
  signal e_12_i_1_n_0 : STD_LOGIC;
  signal e_13_i_1_n_0 : STD_LOGIC;
  signal e_14_i_1_n_0 : STD_LOGIC;
  signal e_15_i_1_n_0 : STD_LOGIC;
  signal e_15_i_3_n_0 : STD_LOGIC;
  signal e_15_i_4_n_0 : STD_LOGIC;
  signal e_15_i_5_n_0 : STD_LOGIC;
  signal e_15_i_6_n_0 : STD_LOGIC;
  signal e_16_i_1_n_0 : STD_LOGIC;
  signal e_17_i_1_n_0 : STD_LOGIC;
  signal e_18_i_1_n_0 : STD_LOGIC;
  signal e_19_i_1_n_0 : STD_LOGIC;
  signal e_19_i_3_n_0 : STD_LOGIC;
  signal e_19_i_4_n_0 : STD_LOGIC;
  signal e_19_i_5_n_0 : STD_LOGIC;
  signal e_19_i_6_n_0 : STD_LOGIC;
  signal e_1_i_1_n_0 : STD_LOGIC;
  signal e_20_i_1_n_0 : STD_LOGIC;
  signal e_21_i_1_n_0 : STD_LOGIC;
  signal e_22_i_1_n_0 : STD_LOGIC;
  signal e_23_i_1_n_0 : STD_LOGIC;
  signal e_23_i_3_n_0 : STD_LOGIC;
  signal e_23_i_4_n_0 : STD_LOGIC;
  signal e_23_i_5_n_0 : STD_LOGIC;
  signal e_23_i_6_n_0 : STD_LOGIC;
  signal e_24_i_1_n_0 : STD_LOGIC;
  signal e_25_i_1_n_0 : STD_LOGIC;
  signal e_26_i_1_n_0 : STD_LOGIC;
  signal e_27_i_1_n_0 : STD_LOGIC;
  signal e_27_i_3_n_0 : STD_LOGIC;
  signal e_27_i_4_n_0 : STD_LOGIC;
  signal e_27_i_5_n_0 : STD_LOGIC;
  signal e_27_i_6_n_0 : STD_LOGIC;
  signal e_28_i_1_n_0 : STD_LOGIC;
  signal e_29_i_1_n_0 : STD_LOGIC;
  signal e_2_i_1_n_0 : STD_LOGIC;
  signal e_30_i_1_n_0 : STD_LOGIC;
  signal e_31_i_1_n_0 : STD_LOGIC;
  signal e_31_i_3_n_0 : STD_LOGIC;
  signal e_31_i_4_n_0 : STD_LOGIC;
  signal e_31_i_5_n_0 : STD_LOGIC;
  signal e_31_i_6_n_0 : STD_LOGIC;
  signal e_3_i_1_n_0 : STD_LOGIC;
  signal e_3_i_3_n_0 : STD_LOGIC;
  signal e_3_i_4_n_0 : STD_LOGIC;
  signal e_3_i_5_n_0 : STD_LOGIC;
  signal e_3_i_6_n_0 : STD_LOGIC;
  signal e_4_i_1_n_0 : STD_LOGIC;
  signal e_5_i_1_n_0 : STD_LOGIC;
  signal e_6_i_1_n_0 : STD_LOGIC;
  signal e_7_i_1_n_0 : STD_LOGIC;
  signal e_7_i_3_n_0 : STD_LOGIC;
  signal e_7_i_4_n_0 : STD_LOGIC;
  signal e_7_i_5_n_0 : STD_LOGIC;
  signal e_7_i_6_n_0 : STD_LOGIC;
  signal e_8_i_1_n_0 : STD_LOGIC;
  signal e_9_i_1_n_0 : STD_LOGIC;
  signal e_reg_11_i_2_n_0 : STD_LOGIC;
  signal e_reg_11_i_2_n_1 : STD_LOGIC;
  signal e_reg_11_i_2_n_2 : STD_LOGIC;
  signal e_reg_11_i_2_n_3 : STD_LOGIC;
  signal e_reg_15_i_2_n_0 : STD_LOGIC;
  signal e_reg_15_i_2_n_1 : STD_LOGIC;
  signal e_reg_15_i_2_n_2 : STD_LOGIC;
  signal e_reg_15_i_2_n_3 : STD_LOGIC;
  signal e_reg_19_i_2_n_0 : STD_LOGIC;
  signal e_reg_19_i_2_n_1 : STD_LOGIC;
  signal e_reg_19_i_2_n_2 : STD_LOGIC;
  signal e_reg_19_i_2_n_3 : STD_LOGIC;
  signal e_reg_23_i_2_n_0 : STD_LOGIC;
  signal e_reg_23_i_2_n_1 : STD_LOGIC;
  signal e_reg_23_i_2_n_2 : STD_LOGIC;
  signal e_reg_23_i_2_n_3 : STD_LOGIC;
  signal e_reg_27_i_2_n_0 : STD_LOGIC;
  signal e_reg_27_i_2_n_1 : STD_LOGIC;
  signal e_reg_27_i_2_n_2 : STD_LOGIC;
  signal e_reg_27_i_2_n_3 : STD_LOGIC;
  signal e_reg_31_i_2_n_1 : STD_LOGIC;
  signal e_reg_31_i_2_n_2 : STD_LOGIC;
  signal e_reg_31_i_2_n_3 : STD_LOGIC;
  signal e_reg_3_i_2_n_0 : STD_LOGIC;
  signal e_reg_3_i_2_n_1 : STD_LOGIC;
  signal e_reg_3_i_2_n_2 : STD_LOGIC;
  signal e_reg_3_i_2_n_3 : STD_LOGIC;
  signal e_reg_7_i_2_n_0 : STD_LOGIC;
  signal e_reg_7_i_2_n_1 : STD_LOGIC;
  signal e_reg_7_i_2_n_2 : STD_LOGIC;
  signal e_reg_7_i_2_n_3 : STD_LOGIC;
  signal finished_OBUF : STD_LOGIC;
  signal FSM_onehot_CURRENT_STATE_0_i_1_n_0 : STD_LOGIC;
  signal FSM_onehot_CURRENT_STATE_10_i_1_n_0 : STD_LOGIC;
  signal FSM_onehot_CURRENT_STATE_11_i_1_n_0 : STD_LOGIC;
  signal FSM_onehot_CURRENT_STATE_11_i_2_n_0 : STD_LOGIC;
  signal FSM_onehot_CURRENT_STATE_11_i_3_n_0 : STD_LOGIC;
  signal FSM_onehot_CURRENT_STATE_11_i_4_n_0 : STD_LOGIC;
  signal FSM_onehot_CURRENT_STATE_11_i_5_n_0 : STD_LOGIC;
  signal FSM_onehot_CURRENT_STATE_11_i_6_n_0 : STD_LOGIC;
  signal FSM_onehot_CURRENT_STATE_11_i_7_n_0 : STD_LOGIC;
  signal FSM_onehot_CURRENT_STATE_11_i_8_n_0 : STD_LOGIC;
  signal FSM_onehot_CURRENT_STATE_11_i_9_n_0 : STD_LOGIC;
  signal FSM_onehot_CURRENT_STATE_11_rep_i_1_n_0 : STD_LOGIC;
  signal FSM_onehot_CURRENT_STATE_1_i_1_n_0 : STD_LOGIC;
  signal FSM_onehot_CURRENT_STATE_2_i_1_n_0 : STD_LOGIC;
  signal FSM_onehot_CURRENT_STATE_8_i_1_n_0 : STD_LOGIC;
  signal FSM_onehot_CURRENT_STATE_9_i_1_n_0 : STD_LOGIC;
  signal FSM_onehot_CURRENT_STATE_reg_11_rep_n_0 : STD_LOGIC;
  signal FSM_onehot_CURRENT_STATE_reg_7_rep_n_0 : STD_LOGIC;
  signal FSM_onehot_CURRENT_STATE_reg_n_0_0 : STD_LOGIC;
  signal FSM_onehot_CURRENT_STATE_reg_n_0_11 : STD_LOGIC;
  signal FSM_onehot_CURRENT_STATE_reg_n_0_12 : STD_LOGIC;
  signal FSM_onehot_CURRENT_STATE_reg_n_0_1 : STD_LOGIC;
  signal FSM_onehot_CURRENT_STATE_reg_n_0_7 : STD_LOGIC;
  signal FSM_onehot_CURRENT_STATE_reg_n_0_8 : STD_LOGIC;
  signal FSM_onehot_CURRENT_STATE_reg_n_0_9 : STD_LOGIC;
  signal f_0_i_1_n_0 : STD_LOGIC;
  signal f_10_i_1_n_0 : STD_LOGIC;
  signal f_11_i_1_n_0 : STD_LOGIC;
  signal f_12_i_1_n_0 : STD_LOGIC;
  signal f_13_i_1_n_0 : STD_LOGIC;
  signal f_14_i_1_n_0 : STD_LOGIC;
  signal f_15_i_1_n_0 : STD_LOGIC;
  signal f_16_i_1_n_0 : STD_LOGIC;
  signal f_17_i_1_n_0 : STD_LOGIC;
  signal f_18_i_1_n_0 : STD_LOGIC;
  signal f_19_i_1_n_0 : STD_LOGIC;
  signal f_1_i_1_n_0 : STD_LOGIC;
  signal f_20_i_1_n_0 : STD_LOGIC;
  signal f_21_i_1_n_0 : STD_LOGIC;
  signal f_22_i_1_n_0 : STD_LOGIC;
  signal f_23_i_1_n_0 : STD_LOGIC;
  signal f_24_i_1_n_0 : STD_LOGIC;
  signal f_25_i_1_n_0 : STD_LOGIC;
  signal f_26_i_1_n_0 : STD_LOGIC;
  signal f_27_i_1_n_0 : STD_LOGIC;
  signal f_28_i_1_n_0 : STD_LOGIC;
  signal f_29_i_1_n_0 : STD_LOGIC;
  signal f_2_i_1_n_0 : STD_LOGIC;
  signal f_30_i_1_n_0 : STD_LOGIC;
  signal f_31_i_1_n_0 : STD_LOGIC;
  signal f_3_i_1_n_0 : STD_LOGIC;
  signal f_4_i_1_n_0 : STD_LOGIC;
  signal f_5_i_1_n_0 : STD_LOGIC;
  signal f_6_i_1_n_0 : STD_LOGIC;
  signal f_7_i_1_n_0 : STD_LOGIC;
  signal f_8_i_1_n_0 : STD_LOGIC;
  signal f_9_i_1_n_0 : STD_LOGIC;
  signal f_reg_n_0_0 : STD_LOGIC;
  signal f_reg_n_0_10 : STD_LOGIC;
  signal f_reg_n_0_11 : STD_LOGIC;
  signal f_reg_n_0_12 : STD_LOGIC;
  signal f_reg_n_0_13 : STD_LOGIC;
  signal f_reg_n_0_14 : STD_LOGIC;
  signal f_reg_n_0_15 : STD_LOGIC;
  signal f_reg_n_0_16 : STD_LOGIC;
  signal f_reg_n_0_17 : STD_LOGIC;
  signal f_reg_n_0_18 : STD_LOGIC;
  signal f_reg_n_0_19 : STD_LOGIC;
  signal f_reg_n_0_1 : STD_LOGIC;
  signal f_reg_n_0_20 : STD_LOGIC;
  signal f_reg_n_0_21 : STD_LOGIC;
  signal f_reg_n_0_22 : STD_LOGIC;
  signal f_reg_n_0_23 : STD_LOGIC;
  signal f_reg_n_0_24 : STD_LOGIC;
  signal f_reg_n_0_25 : STD_LOGIC;
  signal f_reg_n_0_26 : STD_LOGIC;
  signal f_reg_n_0_27 : STD_LOGIC;
  signal f_reg_n_0_28 : STD_LOGIC;
  signal f_reg_n_0_29 : STD_LOGIC;
  signal f_reg_n_0_2 : STD_LOGIC;
  signal f_reg_n_0_30 : STD_LOGIC;
  signal f_reg_n_0_31 : STD_LOGIC;
  signal f_reg_n_0_3 : STD_LOGIC;
  signal f_reg_n_0_4 : STD_LOGIC;
  signal f_reg_n_0_5 : STD_LOGIC;
  signal f_reg_n_0_6 : STD_LOGIC;
  signal f_reg_n_0_7 : STD_LOGIC;
  signal f_reg_n_0_8 : STD_LOGIC;
  signal f_reg_n_0_9 : STD_LOGIC;
  signal g0_b0_n_0 : STD_LOGIC;
  signal g0_b10_n_0 : STD_LOGIC;
  signal g0_b11_n_0 : STD_LOGIC;
  signal g0_b12_n_0 : STD_LOGIC;
  signal g0_b13_n_0 : STD_LOGIC;
  signal g0_b14_n_0 : STD_LOGIC;
  signal g0_b15_n_0 : STD_LOGIC;
  signal g0_b16_n_0 : STD_LOGIC;
  signal g0_b17_n_0 : STD_LOGIC;
  signal g0_b18_n_0 : STD_LOGIC;
  signal g0_b19_n_0 : STD_LOGIC;
  signal g0_b1_n_0 : STD_LOGIC;
  signal g0_b20_n_0 : STD_LOGIC;
  signal g0_b21_n_0 : STD_LOGIC;
  signal g0_b22_n_0 : STD_LOGIC;
  signal g0_b23_n_0 : STD_LOGIC;
  signal g0_b24_n_0 : STD_LOGIC;
  signal g0_b25_n_0 : STD_LOGIC;
  signal g0_b26_n_0 : STD_LOGIC;
  signal g0_b27_n_0 : STD_LOGIC;
  signal g0_b28_n_0 : STD_LOGIC;
  signal g0_b29_n_0 : STD_LOGIC;
  signal g0_b2_n_0 : STD_LOGIC;
  signal g0_b30_n_0 : STD_LOGIC;
  signal g0_b31_n_0 : STD_LOGIC;
  signal g0_b3_n_0 : STD_LOGIC;
  signal g0_b4_n_0 : STD_LOGIC;
  signal g0_b5_n_0 : STD_LOGIC;
  signal g0_b6_n_0 : STD_LOGIC;
  signal g0_b7_n_0 : STD_LOGIC;
  signal g0_b8_n_0 : STD_LOGIC;
  signal g0_b9_n_0 : STD_LOGIC;
  signal g_0_i_1_n_0 : STD_LOGIC;
  signal g_10_i_1_n_0 : STD_LOGIC;
  signal g_11_i_1_n_0 : STD_LOGIC;
  signal g_12_i_1_n_0 : STD_LOGIC;
  signal g_13_i_1_n_0 : STD_LOGIC;
  signal g_14_i_1_n_0 : STD_LOGIC;
  signal g_15_i_1_n_0 : STD_LOGIC;
  signal g_16_i_1_n_0 : STD_LOGIC;
  signal g_17_i_1_n_0 : STD_LOGIC;
  signal g_18_i_1_n_0 : STD_LOGIC;
  signal g_19_i_1_n_0 : STD_LOGIC;
  signal g_1_i_1_n_0 : STD_LOGIC;
  signal g_20_i_1_n_0 : STD_LOGIC;
  signal g_21_i_1_n_0 : STD_LOGIC;
  signal g_22_i_1_n_0 : STD_LOGIC;
  signal g_23_i_1_n_0 : STD_LOGIC;
  signal g_24_i_1_n_0 : STD_LOGIC;
  signal g_25_i_1_n_0 : STD_LOGIC;
  signal g_26_i_1_n_0 : STD_LOGIC;
  signal g_27_i_1_n_0 : STD_LOGIC;
  signal g_28_i_1_n_0 : STD_LOGIC;
  signal g_29_i_1_n_0 : STD_LOGIC;
  signal g_2_i_1_n_0 : STD_LOGIC;
  signal g_30_i_1_n_0 : STD_LOGIC;
  signal g_31_i_1_n_0 : STD_LOGIC;
  signal g_3_i_1_n_0 : STD_LOGIC;
  signal g_4_i_1_n_0 : STD_LOGIC;
  signal g_5_i_1_n_0 : STD_LOGIC;
  signal g_6_i_1_n_0 : STD_LOGIC;
  signal g_7_i_1_n_0 : STD_LOGIC;
  signal g_8_i_1_n_0 : STD_LOGIC;
  signal g_9_i_1_n_0 : STD_LOGIC;
  signal g_reg_n_0_0 : STD_LOGIC;
  signal g_reg_n_0_10 : STD_LOGIC;
  signal g_reg_n_0_11 : STD_LOGIC;
  signal g_reg_n_0_12 : STD_LOGIC;
  signal g_reg_n_0_13 : STD_LOGIC;
  signal g_reg_n_0_14 : STD_LOGIC;
  signal g_reg_n_0_15 : STD_LOGIC;
  signal g_reg_n_0_16 : STD_LOGIC;
  signal g_reg_n_0_17 : STD_LOGIC;
  signal g_reg_n_0_18 : STD_LOGIC;
  signal g_reg_n_0_19 : STD_LOGIC;
  signal g_reg_n_0_1 : STD_LOGIC;
  signal g_reg_n_0_20 : STD_LOGIC;
  signal g_reg_n_0_21 : STD_LOGIC;
  signal g_reg_n_0_22 : STD_LOGIC;
  signal g_reg_n_0_23 : STD_LOGIC;
  signal g_reg_n_0_24 : STD_LOGIC;
  signal g_reg_n_0_25 : STD_LOGIC;
  signal g_reg_n_0_26 : STD_LOGIC;
  signal g_reg_n_0_27 : STD_LOGIC;
  signal g_reg_n_0_28 : STD_LOGIC;
  signal g_reg_n_0_29 : STD_LOGIC;
  signal g_reg_n_0_2 : STD_LOGIC;
  signal g_reg_n_0_30 : STD_LOGIC;
  signal g_reg_n_0_31 : STD_LOGIC;
  signal g_reg_n_0_3 : STD_LOGIC;
  signal g_reg_n_0_4 : STD_LOGIC;
  signal g_reg_n_0_5 : STD_LOGIC;
  signal g_reg_n_0_6 : STD_LOGIC;
  signal g_reg_n_0_7 : STD_LOGIC;
  signal g_reg_n_0_8 : STD_LOGIC;
  signal g_reg_n_0_9 : STD_LOGIC;
  signal h_31 : STD_LOGIC;
  signal h_30 : STD_LOGIC;
  signal h_29 : STD_LOGIC;
  signal h_28 : STD_LOGIC;
  signal h_27 : STD_LOGIC;
  signal h_26 : STD_LOGIC;
  signal h_25 : STD_LOGIC;
  signal h_24 : STD_LOGIC;
  signal h_23 : STD_LOGIC;
  signal h_22 : STD_LOGIC;
  signal h_21 : STD_LOGIC;
  signal h_20 : STD_LOGIC;
  signal h_19 : STD_LOGIC;
  signal h_18 : STD_LOGIC;
  signal h_17 : STD_LOGIC;
  signal h_16 : STD_LOGIC;
  signal h_15 : STD_LOGIC;
  signal h_14 : STD_LOGIC;
  signal h_13 : STD_LOGIC;
  signal h_12 : STD_LOGIC;
  signal h_11 : STD_LOGIC;
  signal h_10 : STD_LOGIC;
  signal h_9 : STD_LOGIC;
  signal h_8 : STD_LOGIC;
  signal h_7 : STD_LOGIC;
  signal h_6 : STD_LOGIC;
  signal h_5 : STD_LOGIC;
  signal h_4 : STD_LOGIC;
  signal h_3 : STD_LOGIC;
  signal h_2 : STD_LOGIC;
  signal h_1 : STD_LOGIC;
  signal h_0 : STD_LOGIC;
  signal HASH_02_COUNTER_30 : STD_LOGIC;
  signal HASH_02_COUNTER_29 : STD_LOGIC;
  signal HASH_02_COUNTER_28 : STD_LOGIC;
  signal HASH_02_COUNTER_27 : STD_LOGIC;
  signal HASH_02_COUNTER_26 : STD_LOGIC;
  signal HASH_02_COUNTER_25 : STD_LOGIC;
  signal HASH_02_COUNTER_24 : STD_LOGIC;
  signal HASH_02_COUNTER_23 : STD_LOGIC;
  signal HASH_02_COUNTER_22 : STD_LOGIC;
  signal HASH_02_COUNTER_21 : STD_LOGIC;
  signal HASH_02_COUNTER_20 : STD_LOGIC;
  signal HASH_02_COUNTER_19 : STD_LOGIC;
  signal HASH_02_COUNTER_18 : STD_LOGIC;
  signal HASH_02_COUNTER_17 : STD_LOGIC;
  signal HASH_02_COUNTER_16 : STD_LOGIC;
  signal HASH_02_COUNTER_15 : STD_LOGIC;
  signal HASH_02_COUNTER_14 : STD_LOGIC;
  signal HASH_02_COUNTER_13 : STD_LOGIC;
  signal HASH_02_COUNTER_12 : STD_LOGIC;
  signal HASH_02_COUNTER_11 : STD_LOGIC;
  signal HASH_02_COUNTER_10 : STD_LOGIC;
  signal HASH_02_COUNTER_9 : STD_LOGIC;
  signal HASH_02_COUNTER_8 : STD_LOGIC;
  signal HASH_02_COUNTER_7 : STD_LOGIC;
  signal HASH_02_COUNTER_6 : STD_LOGIC;
  signal HASH_02_COUNTER_5 : STD_LOGIC;
  signal HASH_02_COUNTER_4 : STD_LOGIC;
  signal HASH_02_COUNTER_3 : STD_LOGIC;
  signal HASH_02_COUNTER_2 : STD_LOGIC;
  signal HASH_02_COUNTER_1 : STD_LOGIC;
  signal HASH_02_COUNTER_0 : STD_LOGIC;
  signal HASH_02_COUNTER_0_i_1_n_0 : STD_LOGIC;
  signal HASH_02_COUNTER_30_i_1_n_0 : STD_LOGIC;
  signal HASH_02_COUNTER_30_i_2_n_0 : STD_LOGIC;
  signal HASH_02_COUNTER_reg_12_i_1_n_0 : STD_LOGIC;
  signal HASH_02_COUNTER_reg_12_i_1_n_1 : STD_LOGIC;
  signal HASH_02_COUNTER_reg_12_i_1_n_2 : STD_LOGIC;
  signal HASH_02_COUNTER_reg_12_i_1_n_3 : STD_LOGIC;
  signal HASH_02_COUNTER_reg_16_i_1_n_0 : STD_LOGIC;
  signal HASH_02_COUNTER_reg_16_i_1_n_1 : STD_LOGIC;
  signal HASH_02_COUNTER_reg_16_i_1_n_2 : STD_LOGIC;
  signal HASH_02_COUNTER_reg_16_i_1_n_3 : STD_LOGIC;
  signal HASH_02_COUNTER_reg_20_i_1_n_0 : STD_LOGIC;
  signal HASH_02_COUNTER_reg_20_i_1_n_1 : STD_LOGIC;
  signal HASH_02_COUNTER_reg_20_i_1_n_2 : STD_LOGIC;
  signal HASH_02_COUNTER_reg_20_i_1_n_3 : STD_LOGIC;
  signal HASH_02_COUNTER_reg_24_i_1_n_0 : STD_LOGIC;
  signal HASH_02_COUNTER_reg_24_i_1_n_1 : STD_LOGIC;
  signal HASH_02_COUNTER_reg_24_i_1_n_2 : STD_LOGIC;
  signal HASH_02_COUNTER_reg_24_i_1_n_3 : STD_LOGIC;
  signal HASH_02_COUNTER_reg_28_i_1_n_0 : STD_LOGIC;
  signal HASH_02_COUNTER_reg_28_i_1_n_1 : STD_LOGIC;
  signal HASH_02_COUNTER_reg_28_i_1_n_2 : STD_LOGIC;
  signal HASH_02_COUNTER_reg_28_i_1_n_3 : STD_LOGIC;
  signal HASH_02_COUNTER_reg_30_i_3_n_3 : STD_LOGIC;
  signal HASH_02_COUNTER_reg_4_i_1_n_0 : STD_LOGIC;
  signal HASH_02_COUNTER_reg_4_i_1_n_1 : STD_LOGIC;
  signal HASH_02_COUNTER_reg_4_i_1_n_2 : STD_LOGIC;
  signal HASH_02_COUNTER_reg_4_i_1_n_3 : STD_LOGIC;
  signal HASH_02_COUNTER_reg_8_i_1_n_0 : STD_LOGIC;
  signal HASH_02_COUNTER_reg_8_i_1_n_1 : STD_LOGIC;
  signal HASH_02_COUNTER_reg_8_i_1_n_2 : STD_LOGIC;
  signal HASH_02_COUNTER_reg_8_i_1_n_3 : STD_LOGIC;
  signal HV_0_0_i_1_n_0 : STD_LOGIC;
  signal HV_0_10_i_1_n_0 : STD_LOGIC;
  signal HV_0_11_i_2_n_0 : STD_LOGIC;
  signal HV_0_11_i_3_n_0 : STD_LOGIC;
  signal HV_0_11_i_4_n_0 : STD_LOGIC;
  signal HV_0_11_i_5_n_0 : STD_LOGIC;
  signal HV_0_12_i_2_n_0 : STD_LOGIC;
  signal HV_0_12_i_3_n_0 : STD_LOGIC;
  signal HV_0_12_i_4_n_0 : STD_LOGIC;
  signal HV_0_12_i_5_n_0 : STD_LOGIC;
  signal HV_0_13_i_1_n_0 : STD_LOGIC;
  signal HV_0_14_i_1_n_0 : STD_LOGIC;
  signal HV_0_15_i_1_n_0 : STD_LOGIC;
  signal HV_0_16_i_1_n_0 : STD_LOGIC;
  signal HV_0_18_i_2_n_0 : STD_LOGIC;
  signal HV_0_18_i_3_n_0 : STD_LOGIC;
  signal HV_0_18_i_4_n_0 : STD_LOGIC;
  signal HV_0_18_i_5_n_0 : STD_LOGIC;
  signal HV_0_19_i_1_n_0 : STD_LOGIC;
  signal HV_0_1_i_1_n_0 : STD_LOGIC;
  signal HV_0_23_i_2_n_0 : STD_LOGIC;
  signal HV_0_23_i_3_n_0 : STD_LOGIC;
  signal HV_0_23_i_4_n_0 : STD_LOGIC;
  signal HV_0_23_i_5_n_0 : STD_LOGIC;
  signal HV_0_25_i_1_n_0 : STD_LOGIC;
  signal HV_0_26_i_2_n_0 : STD_LOGIC;
  signal HV_0_26_i_3_n_0 : STD_LOGIC;
  signal HV_0_26_i_4_n_0 : STD_LOGIC;
  signal HV_0_26_i_5_n_0 : STD_LOGIC;
  signal HV_0_27_i_1_n_0 : STD_LOGIC;
  signal HV_0_29_i_1_n_0 : STD_LOGIC;
  signal HV_0_2_i_1_n_0 : STD_LOGIC;
  signal HV_0_30_i_1_n_0 : STD_LOGIC;
  signal HV_0_31_i_2_n_0 : STD_LOGIC;
  signal HV_0_31_i_3_n_0 : STD_LOGIC;
  signal HV_0_31_i_4_n_0 : STD_LOGIC;
  signal HV_0_31_i_5_n_0 : STD_LOGIC;
  signal HV_0_3_i_2_n_0 : STD_LOGIC;
  signal HV_0_3_i_3_n_0 : STD_LOGIC;
  signal HV_0_3_i_4_n_0 : STD_LOGIC;
  signal HV_0_3_i_5_n_0 : STD_LOGIC;
  signal HV_0_5_i_1_n_0 : STD_LOGIC;
  signal HV_0_6_i_1_n_0 : STD_LOGIC;
  signal HV_0_7_i_2_n_0 : STD_LOGIC;
  signal HV_0_7_i_3_n_0 : STD_LOGIC;
  signal HV_0_7_i_4_n_0 : STD_LOGIC;
  signal HV_0_7_i_5_n_0 : STD_LOGIC;
  signal HV_0_9_i_1_n_0 : STD_LOGIC;
  signal HV_1_0_i_1_n_0 : STD_LOGIC;
  signal HV_1_10_i_1_n_0 : STD_LOGIC;
  signal HV_1_11_i_1_n_0 : STD_LOGIC;
  signal HV_1_13_i_1_n_0 : STD_LOGIC;
  signal HV_1_14_i_2_n_0 : STD_LOGIC;
  signal HV_1_14_i_3_n_0 : STD_LOGIC;
  signal HV_1_14_i_4_n_0 : STD_LOGIC;
  signal HV_1_14_i_5_n_0 : STD_LOGIC;
  signal HV_1_15_i_1_n_0 : STD_LOGIC;
  signal HV_1_16_i_1_n_0 : STD_LOGIC;
  signal HV_1_17_i_1_n_0 : STD_LOGIC;
  signal HV_1_18_i_1_n_0 : STD_LOGIC;
  signal HV_1_19_i_2_n_0 : STD_LOGIC;
  signal HV_1_19_i_3_n_0 : STD_LOGIC;
  signal HV_1_19_i_4_n_0 : STD_LOGIC;
  signal HV_1_19_i_5_n_0 : STD_LOGIC;
  signal HV_1_21_i_1_n_0 : STD_LOGIC;
  signal HV_1_22_i_1_n_0 : STD_LOGIC;
  signal HV_1_23_i_2_n_0 : STD_LOGIC;
  signal HV_1_23_i_3_n_0 : STD_LOGIC;
  signal HV_1_23_i_4_n_0 : STD_LOGIC;
  signal HV_1_23_i_5_n_0 : STD_LOGIC;
  signal HV_1_24_i_1_n_0 : STD_LOGIC;
  signal HV_1_25_i_1_n_0 : STD_LOGIC;
  signal HV_1_26_i_2_n_0 : STD_LOGIC;
  signal HV_1_26_i_3_n_0 : STD_LOGIC;
  signal HV_1_26_i_4_n_0 : STD_LOGIC;
  signal HV_1_26_i_5_n_0 : STD_LOGIC;
  signal HV_1_27_i_1_n_0 : STD_LOGIC;
  signal HV_1_28_i_1_n_0 : STD_LOGIC;
  signal HV_1_29_i_1_n_0 : STD_LOGIC;
  signal HV_1_2_i_1_n_0 : STD_LOGIC;
  signal HV_1_30_i_2_n_0 : STD_LOGIC;
  signal HV_1_30_i_3_n_0 : STD_LOGIC;
  signal HV_1_30_i_4_n_0 : STD_LOGIC;
  signal HV_1_30_i_5_n_0 : STD_LOGIC;
  signal HV_1_31_i_1_n_0 : STD_LOGIC;
  signal HV_1_3_i_2_n_0 : STD_LOGIC;
  signal HV_1_3_i_3_n_0 : STD_LOGIC;
  signal HV_1_3_i_4_n_0 : STD_LOGIC;
  signal HV_1_3_i_5_n_0 : STD_LOGIC;
  signal HV_1_6_i_2_n_0 : STD_LOGIC;
  signal HV_1_6_i_3_n_0 : STD_LOGIC;
  signal HV_1_6_i_4_n_0 : STD_LOGIC;
  signal HV_1_6_i_5_n_0 : STD_LOGIC;
  signal HV_1_7_i_1_n_0 : STD_LOGIC;
  signal HV_1_8_i_2_n_0 : STD_LOGIC;
  signal HV_1_8_i_3_n_0 : STD_LOGIC;
  signal HV_1_8_i_4_n_0 : STD_LOGIC;
  signal HV_1_8_i_5_n_0 : STD_LOGIC;
  signal HV_1_9_i_1_n_0 : STD_LOGIC;
  signal HV_2_11_i_2_n_0 : STD_LOGIC;
  signal HV_2_11_i_3_n_0 : STD_LOGIC;
  signal HV_2_11_i_4_n_0 : STD_LOGIC;
  signal HV_2_11_i_5_n_0 : STD_LOGIC;
  signal HV_2_12_i_1_n_0 : STD_LOGIC;
  signal HV_2_13_i_1_n_0 : STD_LOGIC;
  signal HV_2_14_i_1_n_0 : STD_LOGIC;
  signal HV_2_15_i_1_n_0 : STD_LOGIC;
  signal HV_2_16_i_10_n_0 : STD_LOGIC;
  signal HV_2_16_i_3_n_0 : STD_LOGIC;
  signal HV_2_16_i_4_n_0 : STD_LOGIC;
  signal HV_2_16_i_5_n_0 : STD_LOGIC;
  signal HV_2_16_i_6_n_0 : STD_LOGIC;
  signal HV_2_16_i_7_n_0 : STD_LOGIC;
  signal HV_2_16_i_8_n_0 : STD_LOGIC;
  signal HV_2_16_i_9_n_0 : STD_LOGIC;
  signal HV_2_17_i_1_n_0 : STD_LOGIC;
  signal HV_2_18_i_1_n_0 : STD_LOGIC;
  signal HV_2_19_i_1_n_0 : STD_LOGIC;
  signal HV_2_1_i_1_n_0 : STD_LOGIC;
  signal HV_2_21_i_1_n_0 : STD_LOGIC;
  signal HV_2_22_i_1_n_0 : STD_LOGIC;
  signal HV_2_23_i_2_n_0 : STD_LOGIC;
  signal HV_2_23_i_3_n_0 : STD_LOGIC;
  signal HV_2_23_i_4_n_0 : STD_LOGIC;
  signal HV_2_23_i_5_n_0 : STD_LOGIC;
  signal HV_2_25_i_2_n_0 : STD_LOGIC;
  signal HV_2_25_i_3_n_0 : STD_LOGIC;
  signal HV_2_25_i_4_n_0 : STD_LOGIC;
  signal HV_2_25_i_5_n_0 : STD_LOGIC;
  signal HV_2_26_i_1_n_0 : STD_LOGIC;
  signal HV_2_27_i_1_n_0 : STD_LOGIC;
  signal HV_2_28_i_1_n_0 : STD_LOGIC;
  signal HV_2_29_i_1_n_0 : STD_LOGIC;
  signal HV_2_31_i_2_n_0 : STD_LOGIC;
  signal HV_2_31_i_3_n_0 : STD_LOGIC;
  signal HV_2_31_i_4_n_0 : STD_LOGIC;
  signal HV_2_31_i_5_n_0 : STD_LOGIC;
  signal HV_2_3_i_2_n_0 : STD_LOGIC;
  signal HV_2_3_i_3_n_0 : STD_LOGIC;
  signal HV_2_3_i_4_n_0 : STD_LOGIC;
  signal HV_2_3_i_5_n_0 : STD_LOGIC;
  signal HV_2_4_i_1_n_0 : STD_LOGIC;
  signal HV_2_5_i_1_n_0 : STD_LOGIC;
  signal HV_2_6_i_1_n_0 : STD_LOGIC;
  signal HV_2_7_i_2_n_0 : STD_LOGIC;
  signal HV_2_7_i_3_n_0 : STD_LOGIC;
  signal HV_2_7_i_4_n_0 : STD_LOGIC;
  signal HV_2_7_i_5_n_0 : STD_LOGIC;
  signal HV_2_8_i_1_n_0 : STD_LOGIC;
  signal HV_2_9_i_1_n_0 : STD_LOGIC;
  signal HV_3_10_i_1_n_0 : STD_LOGIC;
  signal HV_3_11_i_2_n_0 : STD_LOGIC;
  signal HV_3_11_i_3_n_0 : STD_LOGIC;
  signal HV_3_11_i_4_n_0 : STD_LOGIC;
  signal HV_3_11_i_5_n_0 : STD_LOGIC;
  signal HV_3_12_i_1_n_0 : STD_LOGIC;
  signal HV_3_13_i_1_n_0 : STD_LOGIC;
  signal HV_3_14_i_1_n_0 : STD_LOGIC;
  signal HV_3_15_i_1_n_0 : STD_LOGIC;
  signal HV_3_15_i_3_n_0 : STD_LOGIC;
  signal HV_3_15_i_4_n_0 : STD_LOGIC;
  signal HV_3_15_i_5_n_0 : STD_LOGIC;
  signal HV_3_15_i_6_n_0 : STD_LOGIC;
  signal HV_3_16_i_1_n_0 : STD_LOGIC;
  signal HV_3_17_i_1_n_0 : STD_LOGIC;
  signal HV_3_18_i_1_n_0 : STD_LOGIC;
  signal HV_3_19_i_1_n_0 : STD_LOGIC;
  signal HV_3_1_i_1_n_0 : STD_LOGIC;
  signal HV_3_22_i_1_n_0 : STD_LOGIC;
  signal HV_3_23_i_10_n_0 : STD_LOGIC;
  signal HV_3_23_i_3_n_0 : STD_LOGIC;
  signal HV_3_23_i_4_n_0 : STD_LOGIC;
  signal HV_3_23_i_5_n_0 : STD_LOGIC;
  signal HV_3_23_i_6_n_0 : STD_LOGIC;
  signal HV_3_23_i_7_n_0 : STD_LOGIC;
  signal HV_3_23_i_8_n_0 : STD_LOGIC;
  signal HV_3_23_i_9_n_0 : STD_LOGIC;
  signal HV_3_24_i_1_n_0 : STD_LOGIC;
  signal HV_3_26_i_1_n_0 : STD_LOGIC;
  signal HV_3_27_i_2_n_0 : STD_LOGIC;
  signal HV_3_27_i_3_n_0 : STD_LOGIC;
  signal HV_3_27_i_4_n_0 : STD_LOGIC;
  signal HV_3_27_i_5_n_0 : STD_LOGIC;
  signal HV_3_29_i_1_n_0 : STD_LOGIC;
  signal HV_3_2_i_2_n_0 : STD_LOGIC;
  signal HV_3_2_i_3_n_0 : STD_LOGIC;
  signal HV_3_2_i_4_n_0 : STD_LOGIC;
  signal HV_3_2_i_5_n_0 : STD_LOGIC;
  signal HV_3_30_i_2_n_0 : STD_LOGIC;
  signal HV_3_30_i_3_n_0 : STD_LOGIC;
  signal HV_3_30_i_4_n_0 : STD_LOGIC;
  signal HV_3_30_i_5_n_0 : STD_LOGIC;
  signal HV_3_31_i_1_n_0 : STD_LOGIC;
  signal HV_3_3_i_1_n_0 : STD_LOGIC;
  signal HV_3_4_i_1_n_0 : STD_LOGIC;
  signal HV_3_5_i_1_n_0 : STD_LOGIC;
  signal HV_3_7_i_2_n_0 : STD_LOGIC;
  signal HV_3_7_i_3_n_0 : STD_LOGIC;
  signal HV_3_7_i_4_n_0 : STD_LOGIC;
  signal HV_3_7_i_5_n_0 : STD_LOGIC;
  signal HV_3_8_i_1_n_0 : STD_LOGIC;
  signal HV_4_0_i_1_n_0 : STD_LOGIC;
  signal HV_4_11_i_2_n_0 : STD_LOGIC;
  signal HV_4_11_i_3_n_0 : STD_LOGIC;
  signal HV_4_11_i_4_n_0 : STD_LOGIC;
  signal HV_4_11_i_5_n_0 : STD_LOGIC;
  signal HV_4_12_i_1_n_0 : STD_LOGIC;
  signal HV_4_14_i_1_n_0 : STD_LOGIC;
  signal HV_4_15_i_2_n_0 : STD_LOGIC;
  signal HV_4_15_i_3_n_0 : STD_LOGIC;
  signal HV_4_15_i_4_n_0 : STD_LOGIC;
  signal HV_4_15_i_5_n_0 : STD_LOGIC;
  signal HV_4_16_i_2_n_0 : STD_LOGIC;
  signal HV_4_16_i_3_n_0 : STD_LOGIC;
  signal HV_4_16_i_4_n_0 : STD_LOGIC;
  signal HV_4_16_i_5_n_0 : STD_LOGIC;
  signal HV_4_17_i_1_n_0 : STD_LOGIC;
  signal HV_4_18_i_1_n_0 : STD_LOGIC;
  signal HV_4_19_i_1_n_0 : STD_LOGIC;
  signal HV_4_1_i_1_n_0 : STD_LOGIC;
  signal HV_4_23_i_2_n_0 : STD_LOGIC;
  signal HV_4_23_i_3_n_0 : STD_LOGIC;
  signal HV_4_23_i_4_n_0 : STD_LOGIC;
  signal HV_4_23_i_5_n_0 : STD_LOGIC;
  signal HV_4_24_i_1_n_0 : STD_LOGIC;
  signal HV_4_27_i_2_n_0 : STD_LOGIC;
  signal HV_4_27_i_3_n_0 : STD_LOGIC;
  signal HV_4_27_i_4_n_0 : STD_LOGIC;
  signal HV_4_27_i_5_n_0 : STD_LOGIC;
  signal HV_4_28_i_1_n_0 : STD_LOGIC;
  signal HV_4_2_i_1_n_0 : STD_LOGIC;
  signal HV_4_30_i_1_n_0 : STD_LOGIC;
  signal HV_4_31_i_2_n_0 : STD_LOGIC;
  signal HV_4_31_i_3_n_0 : STD_LOGIC;
  signal HV_4_31_i_4_n_0 : STD_LOGIC;
  signal HV_4_31_i_5_n_0 : STD_LOGIC;
  signal HV_4_3_i_1_n_0 : STD_LOGIC;
  signal HV_4_4_i_1_n_0 : STD_LOGIC;
  signal HV_4_5_i_1_n_0 : STD_LOGIC;
  signal HV_4_6_i_1_n_0 : STD_LOGIC;
  signal HV_4_7_i_10_n_0 : STD_LOGIC;
  signal HV_4_7_i_3_n_0 : STD_LOGIC;
  signal HV_4_7_i_4_n_0 : STD_LOGIC;
  signal HV_4_7_i_5_n_0 : STD_LOGIC;
  signal HV_4_7_i_6_n_0 : STD_LOGIC;
  signal HV_4_7_i_7_n_0 : STD_LOGIC;
  signal HV_4_7_i_8_n_0 : STD_LOGIC;
  signal HV_4_7_i_9_n_0 : STD_LOGIC;
  signal HV_4_9_i_1_n_0 : STD_LOGIC;
  signal HV_5_10_i_2_n_0 : STD_LOGIC;
  signal HV_5_10_i_3_n_0 : STD_LOGIC;
  signal HV_5_10_i_4_n_0 : STD_LOGIC;
  signal HV_5_10_i_5_n_0 : STD_LOGIC;
  signal HV_5_11_i_1_n_0 : STD_LOGIC;
  signal HV_5_13_i_1_n_0 : STD_LOGIC;
  signal HV_5_14_i_1_n_0 : STD_LOGIC;
  signal HV_5_15_i_2_n_0 : STD_LOGIC;
  signal HV_5_15_i_3_n_0 : STD_LOGIC;
  signal HV_5_15_i_4_n_0 : STD_LOGIC;
  signal HV_5_15_i_5_n_0 : STD_LOGIC;
  signal HV_5_16_i_1_n_0 : STD_LOGIC;
  signal HV_5_18_i_1_n_0 : STD_LOGIC;
  signal HV_5_19_i_2_n_0 : STD_LOGIC;
  signal HV_5_19_i_3_n_0 : STD_LOGIC;
  signal HV_5_19_i_4_n_0 : STD_LOGIC;
  signal HV_5_19_i_5_n_0 : STD_LOGIC;
  signal HV_5_1_i_2_n_0 : STD_LOGIC;
  signal HV_5_1_i_3_n_0 : STD_LOGIC;
  signal HV_5_1_i_4_n_0 : STD_LOGIC;
  signal HV_5_1_i_5_n_0 : STD_LOGIC;
  signal HV_5_23_i_2_n_0 : STD_LOGIC;
  signal HV_5_23_i_3_n_0 : STD_LOGIC;
  signal HV_5_23_i_4_n_0 : STD_LOGIC;
  signal HV_5_23_i_5_n_0 : STD_LOGIC;
  signal HV_5_24_i_1_n_0 : STD_LOGIC;
  signal HV_5_25_i_1_n_0 : STD_LOGIC;
  signal HV_5_26_i_2_n_0 : STD_LOGIC;
  signal HV_5_26_i_3_n_0 : STD_LOGIC;
  signal HV_5_26_i_4_n_0 : STD_LOGIC;
  signal HV_5_26_i_5_n_0 : STD_LOGIC;
  signal HV_5_27_i_1_n_0 : STD_LOGIC;
  signal HV_5_28_i_1_n_0 : STD_LOGIC;
  signal HV_5_2_i_1_n_0 : STD_LOGIC;
  signal HV_5_30_i_2_n_0 : STD_LOGIC;
  signal HV_5_30_i_3_n_0 : STD_LOGIC;
  signal HV_5_30_i_4_n_0 : STD_LOGIC;
  signal HV_5_30_i_5_n_0 : STD_LOGIC;
  signal HV_5_31_i_1_n_0 : STD_LOGIC;
  signal HV_5_3_i_1_n_0 : STD_LOGIC;
  signal HV_5_6_i_2_n_0 : STD_LOGIC;
  signal HV_5_6_i_3_n_0 : STD_LOGIC;
  signal HV_5_6_i_4_n_0 : STD_LOGIC;
  signal HV_5_6_i_5_n_0 : STD_LOGIC;
  signal HV_5_7_i_1_n_0 : STD_LOGIC;
  signal HV_6_0_i_1_n_0 : STD_LOGIC;
  signal HV_6_10_i_2_n_0 : STD_LOGIC;
  signal HV_6_10_i_3_n_0 : STD_LOGIC;
  signal HV_6_10_i_4_n_0 : STD_LOGIC;
  signal HV_6_10_i_5_n_0 : STD_LOGIC;
  signal HV_6_11_i_1_n_0 : STD_LOGIC;
  signal HV_6_12_i_1_n_0 : STD_LOGIC;
  signal HV_6_13_i_2_n_0 : STD_LOGIC;
  signal HV_6_13_i_3_n_0 : STD_LOGIC;
  signal HV_6_13_i_4_n_0 : STD_LOGIC;
  signal HV_6_13_i_5_n_0 : STD_LOGIC;
  signal HV_6_14_i_1_n_0 : STD_LOGIC;
  signal HV_6_15_i_1_n_0 : STD_LOGIC;
  signal HV_6_16_i_1_n_0 : STD_LOGIC;
  signal HV_6_17_i_1_n_0 : STD_LOGIC;
  signal HV_6_19_i_2_n_0 : STD_LOGIC;
  signal HV_6_19_i_3_n_0 : STD_LOGIC;
  signal HV_6_19_i_4_n_0 : STD_LOGIC;
  signal HV_6_19_i_5_n_0 : STD_LOGIC;
  signal HV_6_1_i_1_n_0 : STD_LOGIC;
  signal HV_6_22_i_2_n_0 : STD_LOGIC;
  signal HV_6_22_i_3_n_0 : STD_LOGIC;
  signal HV_6_22_i_4_n_0 : STD_LOGIC;
  signal HV_6_22_i_5_n_0 : STD_LOGIC;
  signal HV_6_23_i_1_n_0 : STD_LOGIC;
  signal HV_6_24_i_1_n_0 : STD_LOGIC;
  signal HV_6_25_i_1_n_0 : STD_LOGIC;
  signal HV_6_26_i_1_n_0 : STD_LOGIC;
  signal HV_6_27_i_1_n_0 : STD_LOGIC;
  signal HV_6_28_i_1_n_0 : STD_LOGIC;
  signal HV_6_28_i_2_n_0 : STD_LOGIC;
  signal HV_6_2_i_2_n_0 : STD_LOGIC;
  signal HV_6_2_i_3_n_0 : STD_LOGIC;
  signal HV_6_2_i_4_n_0 : STD_LOGIC;
  signal HV_6_2_i_5_n_0 : STD_LOGIC;
  signal HV_6_31_i_10_n_0 : STD_LOGIC;
  signal HV_6_31_i_11_n_0 : STD_LOGIC;
  signal HV_6_31_i_12_n_0 : STD_LOGIC;
  signal HV_6_31_i_1_n_0 : STD_LOGIC;
  signal HV_6_31_i_5_n_0 : STD_LOGIC;
  signal HV_6_31_i_6_n_0 : STD_LOGIC;
  signal HV_6_31_i_7_n_0 : STD_LOGIC;
  signal HV_6_31_i_8_n_0 : STD_LOGIC;
  signal HV_6_31_i_9_n_0 : STD_LOGIC;
  signal HV_6_3_i_1_n_0 : STD_LOGIC;
  signal HV_6_5_i_1_n_0 : STD_LOGIC;
  signal HV_6_6_i_2_n_0 : STD_LOGIC;
  signal HV_6_6_i_3_n_0 : STD_LOGIC;
  signal HV_6_6_i_4_n_0 : STD_LOGIC;
  signal HV_6_6_i_5_n_0 : STD_LOGIC;
  signal HV_6_7_i_1_n_0 : STD_LOGIC;
  signal HV_6_8_i_1_n_0 : STD_LOGIC;
  signal HV_7_0_i_1_n_0 : STD_LOGIC;
  signal HV_7_10_i_1_n_0 : STD_LOGIC;
  signal HV_7_11_i_1_n_0 : STD_LOGIC;
  signal HV_7_13_i_2_n_0 : STD_LOGIC;
  signal HV_7_13_i_3_n_0 : STD_LOGIC;
  signal HV_7_13_i_4_n_0 : STD_LOGIC;
  signal HV_7_13_i_5_n_0 : STD_LOGIC;
  signal HV_7_14_i_1_n_0 : STD_LOGIC;
  signal HV_7_15_i_1_n_0 : STD_LOGIC;
  signal HV_7_19_i_2_n_0 : STD_LOGIC;
  signal HV_7_19_i_3_n_0 : STD_LOGIC;
  signal HV_7_19_i_4_n_0 : STD_LOGIC;
  signal HV_7_19_i_5_n_0 : STD_LOGIC;
  signal HV_7_20_i_2_n_0 : STD_LOGIC;
  signal HV_7_20_i_3_n_0 : STD_LOGIC;
  signal HV_7_20_i_4_n_0 : STD_LOGIC;
  signal HV_7_20_i_5_n_0 : STD_LOGIC;
  signal HV_7_21_i_1_n_0 : STD_LOGIC;
  signal HV_7_22_i_1_n_0 : STD_LOGIC;
  signal HV_7_23_i_1_n_0 : STD_LOGIC;
  signal HV_7_24_i_1_n_0 : STD_LOGIC;
  signal HV_7_25_i_1_n_0 : STD_LOGIC;
  signal HV_7_26_i_2_n_0 : STD_LOGIC;
  signal HV_7_26_i_3_n_0 : STD_LOGIC;
  signal HV_7_26_i_4_n_0 : STD_LOGIC;
  signal HV_7_26_i_5_n_0 : STD_LOGIC;
  signal HV_7_27_i_1_n_0 : STD_LOGIC;
  signal HV_7_28_i_1_n_0 : STD_LOGIC;
  signal HV_7_2_i_2_n_0 : STD_LOGIC;
  signal HV_7_2_i_3_n_0 : STD_LOGIC;
  signal HV_7_2_i_4_n_0 : STD_LOGIC;
  signal HV_7_2_i_5_n_0 : STD_LOGIC;
  signal HV_7_30_i_1_n_0 : STD_LOGIC;
  signal HV_7_31_i_2_n_0 : STD_LOGIC;
  signal HV_7_31_i_3_n_0 : STD_LOGIC;
  signal HV_7_31_i_4_n_0 : STD_LOGIC;
  signal HV_7_31_i_5_n_0 : STD_LOGIC;
  signal HV_7_3_i_1_n_0 : STD_LOGIC;
  signal HV_7_4_i_1_n_0 : STD_LOGIC;
  signal HV_7_7_i_2_n_0 : STD_LOGIC;
  signal HV_7_7_i_3_n_0 : STD_LOGIC;
  signal HV_7_7_i_4_n_0 : STD_LOGIC;
  signal HV_7_7_i_5_n_0 : STD_LOGIC;
  signal HV_7_8_i_1_n_0 : STD_LOGIC;
  signal HV_7_9_i_2_n_0 : STD_LOGIC;
  signal HV_7_9_i_3_n_0 : STD_LOGIC;
  signal HV_7_9_i_4_n_0 : STD_LOGIC;
  signal HV_7_9_i_5_n_0 : STD_LOGIC;
  signal HV_reg_0_0 : STD_LOGIC;
  signal HV_reg_0_11_i_1_n_0 : STD_LOGIC;
  signal HV_reg_0_11_i_1_n_1 : STD_LOGIC;
  signal HV_reg_0_11_i_1_n_2 : STD_LOGIC;
  signal HV_reg_0_11_i_1_n_3 : STD_LOGIC;
  signal HV_reg_0_12_i_1_n_0 : STD_LOGIC;
  signal HV_reg_0_12_i_1_n_1 : STD_LOGIC;
  signal HV_reg_0_12_i_1_n_2 : STD_LOGIC;
  signal HV_reg_0_12_i_1_n_3 : STD_LOGIC;
  signal HV_reg_0_18_i_1_n_0 : STD_LOGIC;
  signal HV_reg_0_18_i_1_n_1 : STD_LOGIC;
  signal HV_reg_0_18_i_1_n_2 : STD_LOGIC;
  signal HV_reg_0_18_i_1_n_3 : STD_LOGIC;
  signal HV_reg_0_23_i_1_n_0 : STD_LOGIC;
  signal HV_reg_0_23_i_1_n_1 : STD_LOGIC;
  signal HV_reg_0_23_i_1_n_2 : STD_LOGIC;
  signal HV_reg_0_23_i_1_n_3 : STD_LOGIC;
  signal HV_reg_0_26_i_1_n_0 : STD_LOGIC;
  signal HV_reg_0_26_i_1_n_1 : STD_LOGIC;
  signal HV_reg_0_26_i_1_n_2 : STD_LOGIC;
  signal HV_reg_0_26_i_1_n_3 : STD_LOGIC;
  signal HV_reg_0_31_i_1_n_1 : STD_LOGIC;
  signal HV_reg_0_31_i_1_n_2 : STD_LOGIC;
  signal HV_reg_0_31_i_1_n_3 : STD_LOGIC;
  signal HV_reg_0_3_i_1_n_0 : STD_LOGIC;
  signal HV_reg_0_3_i_1_n_1 : STD_LOGIC;
  signal HV_reg_0_3_i_1_n_2 : STD_LOGIC;
  signal HV_reg_0_3_i_1_n_3 : STD_LOGIC;
  signal HV_reg_0_7_i_1_n_0 : STD_LOGIC;
  signal HV_reg_0_7_i_1_n_1 : STD_LOGIC;
  signal HV_reg_0_7_i_1_n_2 : STD_LOGIC;
  signal HV_reg_0_7_i_1_n_3 : STD_LOGIC;
  signal HV_reg_1_14_i_1_n_0 : STD_LOGIC;
  signal HV_reg_1_14_i_1_n_1 : STD_LOGIC;
  signal HV_reg_1_14_i_1_n_2 : STD_LOGIC;
  signal HV_reg_1_14_i_1_n_3 : STD_LOGIC;
  signal HV_reg_1_19_i_1_n_0 : STD_LOGIC;
  signal HV_reg_1_19_i_1_n_1 : STD_LOGIC;
  signal HV_reg_1_19_i_1_n_2 : STD_LOGIC;
  signal HV_reg_1_19_i_1_n_3 : STD_LOGIC;
  signal HV_reg_1_23_i_1_n_0 : STD_LOGIC;
  signal HV_reg_1_23_i_1_n_1 : STD_LOGIC;
  signal HV_reg_1_23_i_1_n_2 : STD_LOGIC;
  signal HV_reg_1_23_i_1_n_3 : STD_LOGIC;
  signal HV_reg_1_26_i_1_n_0 : STD_LOGIC;
  signal HV_reg_1_26_i_1_n_1 : STD_LOGIC;
  signal HV_reg_1_26_i_1_n_2 : STD_LOGIC;
  signal HV_reg_1_26_i_1_n_3 : STD_LOGIC;
  signal HV_reg_1_30_i_1_n_1 : STD_LOGIC;
  signal HV_reg_1_30_i_1_n_2 : STD_LOGIC;
  signal HV_reg_1_30_i_1_n_3 : STD_LOGIC;
  signal HV_reg_1_3_i_1_n_0 : STD_LOGIC;
  signal HV_reg_1_3_i_1_n_1 : STD_LOGIC;
  signal HV_reg_1_3_i_1_n_2 : STD_LOGIC;
  signal HV_reg_1_3_i_1_n_3 : STD_LOGIC;
  signal HV_reg_1_6_i_1_n_0 : STD_LOGIC;
  signal HV_reg_1_6_i_1_n_1 : STD_LOGIC;
  signal HV_reg_1_6_i_1_n_2 : STD_LOGIC;
  signal HV_reg_1_6_i_1_n_3 : STD_LOGIC;
  signal HV_reg_1_8_i_1_n_0 : STD_LOGIC;
  signal HV_reg_1_8_i_1_n_1 : STD_LOGIC;
  signal HV_reg_1_8_i_1_n_2 : STD_LOGIC;
  signal HV_reg_1_8_i_1_n_3 : STD_LOGIC;
  signal HV_reg_2_11_i_1_n_0 : STD_LOGIC;
  signal HV_reg_2_11_i_1_n_1 : STD_LOGIC;
  signal HV_reg_2_11_i_1_n_2 : STD_LOGIC;
  signal HV_reg_2_11_i_1_n_3 : STD_LOGIC;
  signal HV_reg_2_16_i_1_n_0 : STD_LOGIC;
  signal HV_reg_2_16_i_1_n_1 : STD_LOGIC;
  signal HV_reg_2_16_i_1_n_2 : STD_LOGIC;
  signal HV_reg_2_16_i_1_n_3 : STD_LOGIC;
  signal HV_reg_2_16_i_2_n_0 : STD_LOGIC;
  signal HV_reg_2_16_i_2_n_1 : STD_LOGIC;
  signal HV_reg_2_16_i_2_n_2 : STD_LOGIC;
  signal HV_reg_2_16_i_2_n_3 : STD_LOGIC;
  signal HV_reg_2_23_i_1_n_0 : STD_LOGIC;
  signal HV_reg_2_23_i_1_n_1 : STD_LOGIC;
  signal HV_reg_2_23_i_1_n_2 : STD_LOGIC;
  signal HV_reg_2_23_i_1_n_3 : STD_LOGIC;
  signal HV_reg_2_25_i_1_n_0 : STD_LOGIC;
  signal HV_reg_2_25_i_1_n_1 : STD_LOGIC;
  signal HV_reg_2_25_i_1_n_2 : STD_LOGIC;
  signal HV_reg_2_25_i_1_n_3 : STD_LOGIC;
  signal HV_reg_2_31_i_1_n_1 : STD_LOGIC;
  signal HV_reg_2_31_i_1_n_2 : STD_LOGIC;
  signal HV_reg_2_31_i_1_n_3 : STD_LOGIC;
  signal HV_reg_2_3_i_1_n_0 : STD_LOGIC;
  signal HV_reg_2_3_i_1_n_1 : STD_LOGIC;
  signal HV_reg_2_3_i_1_n_2 : STD_LOGIC;
  signal HV_reg_2_3_i_1_n_3 : STD_LOGIC;
  signal HV_reg_2_7_i_1_n_0 : STD_LOGIC;
  signal HV_reg_2_7_i_1_n_1 : STD_LOGIC;
  signal HV_reg_2_7_i_1_n_2 : STD_LOGIC;
  signal HV_reg_2_7_i_1_n_3 : STD_LOGIC;
  signal HV_reg_3_11_i_1_n_0 : STD_LOGIC;
  signal HV_reg_3_11_i_1_n_1 : STD_LOGIC;
  signal HV_reg_3_11_i_1_n_2 : STD_LOGIC;
  signal HV_reg_3_11_i_1_n_3 : STD_LOGIC;
  signal HV_reg_3_15_i_2_n_0 : STD_LOGIC;
  signal HV_reg_3_15_i_2_n_1 : STD_LOGIC;
  signal HV_reg_3_15_i_2_n_2 : STD_LOGIC;
  signal HV_reg_3_15_i_2_n_3 : STD_LOGIC;
  signal HV_reg_3_23_i_1_n_0 : STD_LOGIC;
  signal HV_reg_3_23_i_1_n_1 : STD_LOGIC;
  signal HV_reg_3_23_i_1_n_2 : STD_LOGIC;
  signal HV_reg_3_23_i_1_n_3 : STD_LOGIC;
  signal HV_reg_3_23_i_2_n_0 : STD_LOGIC;
  signal HV_reg_3_23_i_2_n_1 : STD_LOGIC;
  signal HV_reg_3_23_i_2_n_2 : STD_LOGIC;
  signal HV_reg_3_23_i_2_n_3 : STD_LOGIC;
  signal HV_reg_3_27_i_1_n_0 : STD_LOGIC;
  signal HV_reg_3_27_i_1_n_1 : STD_LOGIC;
  signal HV_reg_3_27_i_1_n_2 : STD_LOGIC;
  signal HV_reg_3_27_i_1_n_3 : STD_LOGIC;
  signal HV_reg_3_2_i_1_n_0 : STD_LOGIC;
  signal HV_reg_3_2_i_1_n_1 : STD_LOGIC;
  signal HV_reg_3_2_i_1_n_2 : STD_LOGIC;
  signal HV_reg_3_2_i_1_n_3 : STD_LOGIC;
  signal HV_reg_3_30_i_1_n_1 : STD_LOGIC;
  signal HV_reg_3_30_i_1_n_2 : STD_LOGIC;
  signal HV_reg_3_30_i_1_n_3 : STD_LOGIC;
  signal HV_reg_3_7_i_1_n_0 : STD_LOGIC;
  signal HV_reg_3_7_i_1_n_1 : STD_LOGIC;
  signal HV_reg_3_7_i_1_n_2 : STD_LOGIC;
  signal HV_reg_3_7_i_1_n_3 : STD_LOGIC;
  signal HV_reg_4_11_i_1_n_0 : STD_LOGIC;
  signal HV_reg_4_11_i_1_n_1 : STD_LOGIC;
  signal HV_reg_4_11_i_1_n_2 : STD_LOGIC;
  signal HV_reg_4_11_i_1_n_3 : STD_LOGIC;
  signal HV_reg_4_15_i_1_n_0 : STD_LOGIC;
  signal HV_reg_4_15_i_1_n_1 : STD_LOGIC;
  signal HV_reg_4_15_i_1_n_2 : STD_LOGIC;
  signal HV_reg_4_15_i_1_n_3 : STD_LOGIC;
  signal HV_reg_4_16_i_1_n_0 : STD_LOGIC;
  signal HV_reg_4_16_i_1_n_1 : STD_LOGIC;
  signal HV_reg_4_16_i_1_n_2 : STD_LOGIC;
  signal HV_reg_4_16_i_1_n_3 : STD_LOGIC;
  signal HV_reg_4_23_i_1_n_0 : STD_LOGIC;
  signal HV_reg_4_23_i_1_n_1 : STD_LOGIC;
  signal HV_reg_4_23_i_1_n_2 : STD_LOGIC;
  signal HV_reg_4_23_i_1_n_3 : STD_LOGIC;
  signal HV_reg_4_27_i_1_n_0 : STD_LOGIC;
  signal HV_reg_4_27_i_1_n_1 : STD_LOGIC;
  signal HV_reg_4_27_i_1_n_2 : STD_LOGIC;
  signal HV_reg_4_27_i_1_n_3 : STD_LOGIC;
  signal HV_reg_4_31_i_1_n_1 : STD_LOGIC;
  signal HV_reg_4_31_i_1_n_2 : STD_LOGIC;
  signal HV_reg_4_31_i_1_n_3 : STD_LOGIC;
  signal HV_reg_4_7_i_1_n_0 : STD_LOGIC;
  signal HV_reg_4_7_i_1_n_1 : STD_LOGIC;
  signal HV_reg_4_7_i_1_n_2 : STD_LOGIC;
  signal HV_reg_4_7_i_1_n_3 : STD_LOGIC;
  signal HV_reg_4_7_i_2_n_0 : STD_LOGIC;
  signal HV_reg_4_7_i_2_n_1 : STD_LOGIC;
  signal HV_reg_4_7_i_2_n_2 : STD_LOGIC;
  signal HV_reg_4_7_i_2_n_3 : STD_LOGIC;
  signal HV_reg_5_10_i_1_n_0 : STD_LOGIC;
  signal HV_reg_5_10_i_1_n_1 : STD_LOGIC;
  signal HV_reg_5_10_i_1_n_2 : STD_LOGIC;
  signal HV_reg_5_10_i_1_n_3 : STD_LOGIC;
  signal HV_reg_5_15_i_1_n_0 : STD_LOGIC;
  signal HV_reg_5_15_i_1_n_1 : STD_LOGIC;
  signal HV_reg_5_15_i_1_n_2 : STD_LOGIC;
  signal HV_reg_5_15_i_1_n_3 : STD_LOGIC;
  signal HV_reg_5_19_i_1_n_0 : STD_LOGIC;
  signal HV_reg_5_19_i_1_n_1 : STD_LOGIC;
  signal HV_reg_5_19_i_1_n_2 : STD_LOGIC;
  signal HV_reg_5_19_i_1_n_3 : STD_LOGIC;
  signal HV_reg_5_1_i_1_n_0 : STD_LOGIC;
  signal HV_reg_5_1_i_1_n_1 : STD_LOGIC;
  signal HV_reg_5_1_i_1_n_2 : STD_LOGIC;
  signal HV_reg_5_1_i_1_n_3 : STD_LOGIC;
  signal HV_reg_5_23_i_1_n_0 : STD_LOGIC;
  signal HV_reg_5_23_i_1_n_1 : STD_LOGIC;
  signal HV_reg_5_23_i_1_n_2 : STD_LOGIC;
  signal HV_reg_5_23_i_1_n_3 : STD_LOGIC;
  signal HV_reg_5_26_i_1_n_0 : STD_LOGIC;
  signal HV_reg_5_26_i_1_n_1 : STD_LOGIC;
  signal HV_reg_5_26_i_1_n_2 : STD_LOGIC;
  signal HV_reg_5_26_i_1_n_3 : STD_LOGIC;
  signal HV_reg_5_30_i_1_n_1 : STD_LOGIC;
  signal HV_reg_5_30_i_1_n_2 : STD_LOGIC;
  signal HV_reg_5_30_i_1_n_3 : STD_LOGIC;
  signal HV_reg_5_6_i_1_n_0 : STD_LOGIC;
  signal HV_reg_5_6_i_1_n_1 : STD_LOGIC;
  signal HV_reg_5_6_i_1_n_2 : STD_LOGIC;
  signal HV_reg_5_6_i_1_n_3 : STD_LOGIC;
  signal HV_reg_6_10_i_1_n_0 : STD_LOGIC;
  signal HV_reg_6_10_i_1_n_1 : STD_LOGIC;
  signal HV_reg_6_10_i_1_n_2 : STD_LOGIC;
  signal HV_reg_6_10_i_1_n_3 : STD_LOGIC;
  signal HV_reg_6_13_i_1_n_0 : STD_LOGIC;
  signal HV_reg_6_13_i_1_n_1 : STD_LOGIC;
  signal HV_reg_6_13_i_1_n_2 : STD_LOGIC;
  signal HV_reg_6_13_i_1_n_3 : STD_LOGIC;
  signal HV_reg_6_19_i_1_n_0 : STD_LOGIC;
  signal HV_reg_6_19_i_1_n_1 : STD_LOGIC;
  signal HV_reg_6_19_i_1_n_2 : STD_LOGIC;
  signal HV_reg_6_19_i_1_n_3 : STD_LOGIC;
  signal HV_reg_6_22_i_1_n_0 : STD_LOGIC;
  signal HV_reg_6_22_i_1_n_1 : STD_LOGIC;
  signal HV_reg_6_22_i_1_n_2 : STD_LOGIC;
  signal HV_reg_6_22_i_1_n_3 : STD_LOGIC;
  signal HV_reg_6_2_i_1_n_0 : STD_LOGIC;
  signal HV_reg_6_2_i_1_n_1 : STD_LOGIC;
  signal HV_reg_6_2_i_1_n_2 : STD_LOGIC;
  signal HV_reg_6_2_i_1_n_3 : STD_LOGIC;
  signal HV_reg_6_31_i_3_n_1 : STD_LOGIC;
  signal HV_reg_6_31_i_3_n_2 : STD_LOGIC;
  signal HV_reg_6_31_i_3_n_3 : STD_LOGIC;
  signal HV_reg_6_31_i_4_n_0 : STD_LOGIC;
  signal HV_reg_6_31_i_4_n_1 : STD_LOGIC;
  signal HV_reg_6_31_i_4_n_2 : STD_LOGIC;
  signal HV_reg_6_31_i_4_n_3 : STD_LOGIC;
  signal HV_reg_6_6_i_1_n_0 : STD_LOGIC;
  signal HV_reg_6_6_i_1_n_1 : STD_LOGIC;
  signal HV_reg_6_6_i_1_n_2 : STD_LOGIC;
  signal HV_reg_6_6_i_1_n_3 : STD_LOGIC;
  signal HV_reg_7_13_i_1_n_0 : STD_LOGIC;
  signal HV_reg_7_13_i_1_n_1 : STD_LOGIC;
  signal HV_reg_7_13_i_1_n_2 : STD_LOGIC;
  signal HV_reg_7_13_i_1_n_3 : STD_LOGIC;
  signal HV_reg_7_19_i_1_n_0 : STD_LOGIC;
  signal HV_reg_7_19_i_1_n_1 : STD_LOGIC;
  signal HV_reg_7_19_i_1_n_2 : STD_LOGIC;
  signal HV_reg_7_19_i_1_n_3 : STD_LOGIC;
  signal HV_reg_7_20_i_1_n_0 : STD_LOGIC;
  signal HV_reg_7_20_i_1_n_1 : STD_LOGIC;
  signal HV_reg_7_20_i_1_n_2 : STD_LOGIC;
  signal HV_reg_7_20_i_1_n_3 : STD_LOGIC;
  signal HV_reg_7_26_i_1_n_0 : STD_LOGIC;
  signal HV_reg_7_26_i_1_n_1 : STD_LOGIC;
  signal HV_reg_7_26_i_1_n_2 : STD_LOGIC;
  signal HV_reg_7_26_i_1_n_3 : STD_LOGIC;
  signal HV_reg_7_2_i_1_n_0 : STD_LOGIC;
  signal HV_reg_7_2_i_1_n_1 : STD_LOGIC;
  signal HV_reg_7_2_i_1_n_2 : STD_LOGIC;
  signal HV_reg_7_2_i_1_n_3 : STD_LOGIC;
  signal HV_reg_7_31_i_1_n_1 : STD_LOGIC;
  signal HV_reg_7_31_i_1_n_2 : STD_LOGIC;
  signal HV_reg_7_31_i_1_n_3 : STD_LOGIC;
  signal HV_reg_7_7_i_1_n_0 : STD_LOGIC;
  signal HV_reg_7_7_i_1_n_1 : STD_LOGIC;
  signal HV_reg_7_7_i_1_n_2 : STD_LOGIC;
  signal HV_reg_7_7_i_1_n_3 : STD_LOGIC;
  signal HV_reg_7_9_i_1_n_0 : STD_LOGIC;
  signal HV_reg_7_9_i_1_n_1 : STD_LOGIC;
  signal HV_reg_7_9_i_1_n_2 : STD_LOGIC;
  signal HV_reg_7_9_i_1_n_3 : STD_LOGIC;
  signal h_0_i_1_n_0 : STD_LOGIC;
  signal h_10_i_1_n_0 : STD_LOGIC;
  signal h_11_i_1_n_0 : STD_LOGIC;
  signal h_12_i_1_n_0 : STD_LOGIC;
  signal h_13_i_1_n_0 : STD_LOGIC;
  signal h_14_i_1_n_0 : STD_LOGIC;
  signal h_15_i_1_n_0 : STD_LOGIC;
  signal h_16_i_1_n_0 : STD_LOGIC;
  signal h_17_i_1_n_0 : STD_LOGIC;
  signal h_18_i_1_n_0 : STD_LOGIC;
  signal h_19_i_1_n_0 : STD_LOGIC;
  signal h_1_i_1_n_0 : STD_LOGIC;
  signal h_20_i_1_n_0 : STD_LOGIC;
  signal h_21_i_1_n_0 : STD_LOGIC;
  signal h_22_i_1_n_0 : STD_LOGIC;
  signal h_23_i_1_n_0 : STD_LOGIC;
  signal h_24_i_1_n_0 : STD_LOGIC;
  signal h_25_i_1_n_0 : STD_LOGIC;
  signal h_26_i_1_n_0 : STD_LOGIC;
  signal h_27_i_1_n_0 : STD_LOGIC;
  signal h_28_i_1_n_0 : STD_LOGIC;
  signal h_29_i_1_n_0 : STD_LOGIC;
  signal h_2_i_1_n_0 : STD_LOGIC;
  signal h_30_i_1_n_0 : STD_LOGIC;
  signal h_31_i_1_n_0 : STD_LOGIC;
  signal h_3_i_1_n_0 : STD_LOGIC;
  signal h_4_i_1_n_0 : STD_LOGIC;
  signal h_5_i_1_n_0 : STD_LOGIC;
  signal h_6_i_1_n_0 : STD_LOGIC;
  signal h_7_i_1_n_0 : STD_LOGIC;
  signal h_8_i_1_n_0 : STD_LOGIC;
  signal h_9_i_1_n_0 : STD_LOGIC;
  signal in15_31 : STD_LOGIC;
  signal in15_30 : STD_LOGIC;
  signal in15_29 : STD_LOGIC;
  signal in15_28 : STD_LOGIC;
  signal in15_27 : STD_LOGIC;
  signal in15_26 : STD_LOGIC;
  signal in15_25 : STD_LOGIC;
  signal in15_24 : STD_LOGIC;
  signal in15_23 : STD_LOGIC;
  signal in15_22 : STD_LOGIC;
  signal in15_21 : STD_LOGIC;
  signal in15_20 : STD_LOGIC;
  signal in15_19 : STD_LOGIC;
  signal in15_18 : STD_LOGIC;
  signal in15_17 : STD_LOGIC;
  signal in15_16 : STD_LOGIC;
  signal in15_15 : STD_LOGIC;
  signal in15_14 : STD_LOGIC;
  signal in15_13 : STD_LOGIC;
  signal in15_12 : STD_LOGIC;
  signal in15_11 : STD_LOGIC;
  signal in15_10 : STD_LOGIC;
  signal in15_9 : STD_LOGIC;
  signal in15_8 : STD_LOGIC;
  signal in15_7 : STD_LOGIC;
  signal in15_6 : STD_LOGIC;
  signal in15_5 : STD_LOGIC;
  signal in15_4 : STD_LOGIC;
  signal in15_3 : STD_LOGIC;
  signal in15_2 : STD_LOGIC;
  signal in15_1 : STD_LOGIC;
  signal in15_0 : STD_LOGIC;
  signal in23_31 : STD_LOGIC;
  signal in23_30 : STD_LOGIC;
  signal in23_29 : STD_LOGIC;
  signal in23_28 : STD_LOGIC;
  signal in23_27 : STD_LOGIC;
  signal in23_26 : STD_LOGIC;
  signal in23_25 : STD_LOGIC;
  signal in23_24 : STD_LOGIC;
  signal in23_23 : STD_LOGIC;
  signal in23_22 : STD_LOGIC;
  signal in23_21 : STD_LOGIC;
  signal in23_20 : STD_LOGIC;
  signal in23_19 : STD_LOGIC;
  signal in23_18 : STD_LOGIC;
  signal in23_17 : STD_LOGIC;
  signal in23_16 : STD_LOGIC;
  signal in23_15 : STD_LOGIC;
  signal in23_14 : STD_LOGIC;
  signal in23_13 : STD_LOGIC;
  signal in23_12 : STD_LOGIC;
  signal in23_11 : STD_LOGIC;
  signal in23_10 : STD_LOGIC;
  signal in23_9 : STD_LOGIC;
  signal in23_8 : STD_LOGIC;
  signal in23_7 : STD_LOGIC;
  signal in23_6 : STD_LOGIC;
  signal in23_5 : STD_LOGIC;
  signal in23_4 : STD_LOGIC;
  signal in23_3 : STD_LOGIC;
  signal in23_2 : STD_LOGIC;
  signal in23_1 : STD_LOGIC;
  signal in23_0 : STD_LOGIC;
  signal in25_31 : STD_LOGIC;
  signal in25_30 : STD_LOGIC;
  signal in25_29 : STD_LOGIC;
  signal in25_28 : STD_LOGIC;
  signal in25_27 : STD_LOGIC;
  signal in25_26 : STD_LOGIC;
  signal in25_25 : STD_LOGIC;
  signal in25_24 : STD_LOGIC;
  signal in25_23 : STD_LOGIC;
  signal in25_22 : STD_LOGIC;
  signal in25_21 : STD_LOGIC;
  signal in25_20 : STD_LOGIC;
  signal in25_19 : STD_LOGIC;
  signal in25_18 : STD_LOGIC;
  signal in25_17 : STD_LOGIC;
  signal in25_16 : STD_LOGIC;
  signal in25_15 : STD_LOGIC;
  signal in25_14 : STD_LOGIC;
  signal in25_13 : STD_LOGIC;
  signal in25_12 : STD_LOGIC;
  signal in25_11 : STD_LOGIC;
  signal in25_10 : STD_LOGIC;
  signal in25_9 : STD_LOGIC;
  signal in25_8 : STD_LOGIC;
  signal in25_7 : STD_LOGIC;
  signal in25_6 : STD_LOGIC;
  signal in25_5 : STD_LOGIC;
  signal in25_4 : STD_LOGIC;
  signal in25_3 : STD_LOGIC;
  signal in25_2 : STD_LOGIC;
  signal in25_1 : STD_LOGIC;
  signal in25_0 : STD_LOGIC;
  signal in26_31 : STD_LOGIC;
  signal in26_30 : STD_LOGIC;
  signal in26_29 : STD_LOGIC;
  signal in26_28 : STD_LOGIC;
  signal in26_27 : STD_LOGIC;
  signal in26_26 : STD_LOGIC;
  signal in26_25 : STD_LOGIC;
  signal in26_24 : STD_LOGIC;
  signal in26_23 : STD_LOGIC;
  signal in26_22 : STD_LOGIC;
  signal in26_21 : STD_LOGIC;
  signal in26_20 : STD_LOGIC;
  signal in26_19 : STD_LOGIC;
  signal in26_18 : STD_LOGIC;
  signal in26_17 : STD_LOGIC;
  signal in26_16 : STD_LOGIC;
  signal in26_15 : STD_LOGIC;
  signal in26_14 : STD_LOGIC;
  signal in26_13 : STD_LOGIC;
  signal in26_12 : STD_LOGIC;
  signal in26_11 : STD_LOGIC;
  signal in26_10 : STD_LOGIC;
  signal in26_9 : STD_LOGIC;
  signal in26_8 : STD_LOGIC;
  signal in26_7 : STD_LOGIC;
  signal in26_6 : STD_LOGIC;
  signal in26_5 : STD_LOGIC;
  signal in26_4 : STD_LOGIC;
  signal in26_3 : STD_LOGIC;
  signal in26_2 : STD_LOGIC;
  signal in26_1 : STD_LOGIC;
  signal in26_0 : STD_LOGIC;
  signal in27_31 : STD_LOGIC;
  signal in27_30 : STD_LOGIC;
  signal in27_29 : STD_LOGIC;
  signal in27_28 : STD_LOGIC;
  signal in27_27 : STD_LOGIC;
  signal in27_26 : STD_LOGIC;
  signal in27_25 : STD_LOGIC;
  signal in27_24 : STD_LOGIC;
  signal in27_23 : STD_LOGIC;
  signal in27_22 : STD_LOGIC;
  signal in27_21 : STD_LOGIC;
  signal in27_20 : STD_LOGIC;
  signal in27_19 : STD_LOGIC;
  signal in27_18 : STD_LOGIC;
  signal in27_17 : STD_LOGIC;
  signal in27_16 : STD_LOGIC;
  signal in27_15 : STD_LOGIC;
  signal in27_14 : STD_LOGIC;
  signal in27_13 : STD_LOGIC;
  signal in27_12 : STD_LOGIC;
  signal in27_11 : STD_LOGIC;
  signal in27_10 : STD_LOGIC;
  signal in27_9 : STD_LOGIC;
  signal in27_8 : STD_LOGIC;
  signal in27_7 : STD_LOGIC;
  signal in27_6 : STD_LOGIC;
  signal in27_5 : STD_LOGIC;
  signal in27_4 : STD_LOGIC;
  signal in27_3 : STD_LOGIC;
  signal in27_2 : STD_LOGIC;
  signal in27_1 : STD_LOGIC;
  signal in27_0 : STD_LOGIC;
  signal in28_31 : STD_LOGIC;
  signal in28_30 : STD_LOGIC;
  signal in28_29 : STD_LOGIC;
  signal in28_28 : STD_LOGIC;
  signal in28_27 : STD_LOGIC;
  signal in28_26 : STD_LOGIC;
  signal in28_25 : STD_LOGIC;
  signal in28_24 : STD_LOGIC;
  signal in28_23 : STD_LOGIC;
  signal in28_22 : STD_LOGIC;
  signal in28_21 : STD_LOGIC;
  signal in28_20 : STD_LOGIC;
  signal in28_19 : STD_LOGIC;
  signal in28_18 : STD_LOGIC;
  signal in28_17 : STD_LOGIC;
  signal in28_16 : STD_LOGIC;
  signal in28_15 : STD_LOGIC;
  signal in28_14 : STD_LOGIC;
  signal in28_13 : STD_LOGIC;
  signal in28_12 : STD_LOGIC;
  signal in28_11 : STD_LOGIC;
  signal in28_10 : STD_LOGIC;
  signal in28_9 : STD_LOGIC;
  signal in28_8 : STD_LOGIC;
  signal in28_7 : STD_LOGIC;
  signal in28_6 : STD_LOGIC;
  signal in28_5 : STD_LOGIC;
  signal in28_4 : STD_LOGIC;
  signal in28_3 : STD_LOGIC;
  signal in28_2 : STD_LOGIC;
  signal in28_1 : STD_LOGIC;
  signal in28_0 : STD_LOGIC;
  signal in29_31 : STD_LOGIC;
  signal in29_30 : STD_LOGIC;
  signal in29_29 : STD_LOGIC;
  signal in29_28 : STD_LOGIC;
  signal in29_27 : STD_LOGIC;
  signal in29_26 : STD_LOGIC;
  signal in29_25 : STD_LOGIC;
  signal in29_24 : STD_LOGIC;
  signal in29_23 : STD_LOGIC;
  signal in29_22 : STD_LOGIC;
  signal in29_21 : STD_LOGIC;
  signal in29_20 : STD_LOGIC;
  signal in29_19 : STD_LOGIC;
  signal in29_18 : STD_LOGIC;
  signal in29_17 : STD_LOGIC;
  signal in29_16 : STD_LOGIC;
  signal in29_15 : STD_LOGIC;
  signal in29_14 : STD_LOGIC;
  signal in29_13 : STD_LOGIC;
  signal in29_12 : STD_LOGIC;
  signal in29_11 : STD_LOGIC;
  signal in29_10 : STD_LOGIC;
  signal in29_9 : STD_LOGIC;
  signal in29_8 : STD_LOGIC;
  signal in29_7 : STD_LOGIC;
  signal in29_6 : STD_LOGIC;
  signal in29_5 : STD_LOGIC;
  signal in29_4 : STD_LOGIC;
  signal in29_3 : STD_LOGIC;
  signal in29_2 : STD_LOGIC;
  signal in29_1 : STD_LOGIC;
  signal in29_0 : STD_LOGIC;
  signal in30_31 : STD_LOGIC;
  signal in30_30 : STD_LOGIC;
  signal in30_29 : STD_LOGIC;
  signal in30_28 : STD_LOGIC;
  signal in30_27 : STD_LOGIC;
  signal in30_26 : STD_LOGIC;
  signal in30_25 : STD_LOGIC;
  signal in30_24 : STD_LOGIC;
  signal in30_23 : STD_LOGIC;
  signal in30_22 : STD_LOGIC;
  signal in30_21 : STD_LOGIC;
  signal in30_20 : STD_LOGIC;
  signal in30_19 : STD_LOGIC;
  signal in30_18 : STD_LOGIC;
  signal in30_17 : STD_LOGIC;
  signal in30_16 : STD_LOGIC;
  signal in30_15 : STD_LOGIC;
  signal in30_14 : STD_LOGIC;
  signal in30_13 : STD_LOGIC;
  signal in30_12 : STD_LOGIC;
  signal in30_11 : STD_LOGIC;
  signal in30_10 : STD_LOGIC;
  signal in30_9 : STD_LOGIC;
  signal in30_8 : STD_LOGIC;
  signal in30_7 : STD_LOGIC;
  signal in30_6 : STD_LOGIC;
  signal in30_5 : STD_LOGIC;
  signal in30_4 : STD_LOGIC;
  signal in30_3 : STD_LOGIC;
  signal in30_2 : STD_LOGIC;
  signal in30_1 : STD_LOGIC;
  signal in30_0 : STD_LOGIC;
  signal in31_31 : STD_LOGIC;
  signal in31_30 : STD_LOGIC;
  signal in31_29 : STD_LOGIC;
  signal in31_28 : STD_LOGIC;
  signal in31_27 : STD_LOGIC;
  signal in31_26 : STD_LOGIC;
  signal in31_25 : STD_LOGIC;
  signal in31_24 : STD_LOGIC;
  signal in31_23 : STD_LOGIC;
  signal in31_22 : STD_LOGIC;
  signal in31_21 : STD_LOGIC;
  signal in31_20 : STD_LOGIC;
  signal in31_19 : STD_LOGIC;
  signal in31_18 : STD_LOGIC;
  signal in31_17 : STD_LOGIC;
  signal in31_16 : STD_LOGIC;
  signal in31_15 : STD_LOGIC;
  signal in31_14 : STD_LOGIC;
  signal in31_13 : STD_LOGIC;
  signal in31_12 : STD_LOGIC;
  signal in31_11 : STD_LOGIC;
  signal in31_10 : STD_LOGIC;
  signal in31_9 : STD_LOGIC;
  signal in31_8 : STD_LOGIC;
  signal in31_7 : STD_LOGIC;
  signal in31_6 : STD_LOGIC;
  signal in31_5 : STD_LOGIC;
  signal in31_4 : STD_LOGIC;
  signal in31_3 : STD_LOGIC;
  signal in31_2 : STD_LOGIC;
  signal in31_1 : STD_LOGIC;
  signal in31_0 : STD_LOGIC;
  signal in32_30 : STD_LOGIC;
  signal in32_29 : STD_LOGIC;
  signal in32_28 : STD_LOGIC;
  signal in32_27 : STD_LOGIC;
  signal in32_26 : STD_LOGIC;
  signal in32_25 : STD_LOGIC;
  signal in32_24 : STD_LOGIC;
  signal in32_23 : STD_LOGIC;
  signal in32_22 : STD_LOGIC;
  signal in32_21 : STD_LOGIC;
  signal in32_20 : STD_LOGIC;
  signal in32_19 : STD_LOGIC;
  signal in32_18 : STD_LOGIC;
  signal in32_17 : STD_LOGIC;
  signal in32_16 : STD_LOGIC;
  signal in32_15 : STD_LOGIC;
  signal in32_14 : STD_LOGIC;
  signal in32_13 : STD_LOGIC;
  signal in32_12 : STD_LOGIC;
  signal in32_11 : STD_LOGIC;
  signal in32_10 : STD_LOGIC;
  signal in32_9 : STD_LOGIC;
  signal in32_8 : STD_LOGIC;
  signal in32_7 : STD_LOGIC;
  signal in32_6 : STD_LOGIC;
  signal in32_5 : STD_LOGIC;
  signal in32_4 : STD_LOGIC;
  signal in32_3 : STD_LOGIC;
  signal in32_2 : STD_LOGIC;
  signal in32_1 : STD_LOGIC;
  signal in7_31 : STD_LOGIC;
  signal in7_30 : STD_LOGIC;
  signal in7_29 : STD_LOGIC;
  signal in7_28 : STD_LOGIC;
  signal in7_27 : STD_LOGIC;
  signal in7_26 : STD_LOGIC;
  signal in7_25 : STD_LOGIC;
  signal in7_24 : STD_LOGIC;
  signal in7_23 : STD_LOGIC;
  signal in7_22 : STD_LOGIC;
  signal in7_21 : STD_LOGIC;
  signal in7_20 : STD_LOGIC;
  signal in7_19 : STD_LOGIC;
  signal in7_18 : STD_LOGIC;
  signal in7_17 : STD_LOGIC;
  signal in7_16 : STD_LOGIC;
  signal in7_15 : STD_LOGIC;
  signal in7_14 : STD_LOGIC;
  signal in7_13 : STD_LOGIC;
  signal in7_12 : STD_LOGIC;
  signal in7_11 : STD_LOGIC;
  signal in7_10 : STD_LOGIC;
  signal in7_9 : STD_LOGIC;
  signal in7_8 : STD_LOGIC;
  signal in7_7 : STD_LOGIC;
  signal in7_6 : STD_LOGIC;
  signal in7_5 : STD_LOGIC;
  signal in7_4 : STD_LOGIC;
  signal in7_3 : STD_LOGIC;
  signal in7_2 : STD_LOGIC;
  signal in7_1 : STD_LOGIC;
  signal in7_0 : STD_LOGIC;
  signal msg_block_in_IBUF_0 : STD_LOGIC;
  signal msg_block_in_IBUF_1 : STD_LOGIC;
  signal msg_block_in_IBUF_2 : STD_LOGIC;
  signal msg_block_in_IBUF_3 : STD_LOGIC;
  signal msg_block_in_IBUF_4 : STD_LOGIC;
  signal msg_block_in_IBUF_5 : STD_LOGIC;
  signal msg_block_in_IBUF_6 : STD_LOGIC;
  signal msg_block_in_IBUF_7 : STD_LOGIC;
  signal msg_block_in_IBUF_8 : STD_LOGIC;
  signal msg_block_in_IBUF_9 : STD_LOGIC;
  signal msg_block_in_IBUF_10 : STD_LOGIC;
  signal msg_block_in_IBUF_11 : STD_LOGIC;
  signal msg_block_in_IBUF_12 : STD_LOGIC;
  signal msg_block_in_IBUF_13 : STD_LOGIC;
  signal msg_block_in_IBUF_14 : STD_LOGIC;
  signal msg_block_in_IBUF_15 : STD_LOGIC;
  signal msg_block_in_IBUF_16 : STD_LOGIC;
  signal msg_block_in_IBUF_17 : STD_LOGIC;
  signal msg_block_in_IBUF_18 : STD_LOGIC;
  signal msg_block_in_IBUF_19 : STD_LOGIC;
  signal msg_block_in_IBUF_20 : STD_LOGIC;
  signal msg_block_in_IBUF_21 : STD_LOGIC;
  signal msg_block_in_IBUF_22 : STD_LOGIC;
  signal msg_block_in_IBUF_23 : STD_LOGIC;
  signal msg_block_in_IBUF_24 : STD_LOGIC;
  signal msg_block_in_IBUF_25 : STD_LOGIC;
  signal msg_block_in_IBUF_26 : STD_LOGIC;
  signal msg_block_in_IBUF_27 : STD_LOGIC;
  signal msg_block_in_IBUF_28 : STD_LOGIC;
  signal msg_block_in_IBUF_29 : STD_LOGIC;
  signal msg_block_in_IBUF_30 : STD_LOGIC;
  signal msg_block_in_IBUF_31 : STD_LOGIC;
  signal msg_block_in_IBUF_32 : STD_LOGIC;
  signal msg_block_in_IBUF_33 : STD_LOGIC;
  signal msg_block_in_IBUF_34 : STD_LOGIC;
  signal msg_block_in_IBUF_35 : STD_LOGIC;
  signal msg_block_in_IBUF_36 : STD_LOGIC;
  signal msg_block_in_IBUF_37 : STD_LOGIC;
  signal msg_block_in_IBUF_38 : STD_LOGIC;
  signal msg_block_in_IBUF_39 : STD_LOGIC;
  signal msg_block_in_IBUF_40 : STD_LOGIC;
  signal msg_block_in_IBUF_41 : STD_LOGIC;
  signal msg_block_in_IBUF_42 : STD_LOGIC;
  signal msg_block_in_IBUF_43 : STD_LOGIC;
  signal msg_block_in_IBUF_44 : STD_LOGIC;
  signal msg_block_in_IBUF_45 : STD_LOGIC;
  signal msg_block_in_IBUF_46 : STD_LOGIC;
  signal msg_block_in_IBUF_47 : STD_LOGIC;
  signal msg_block_in_IBUF_48 : STD_LOGIC;
  signal msg_block_in_IBUF_49 : STD_LOGIC;
  signal msg_block_in_IBUF_50 : STD_LOGIC;
  signal msg_block_in_IBUF_51 : STD_LOGIC;
  signal msg_block_in_IBUF_52 : STD_LOGIC;
  signal msg_block_in_IBUF_53 : STD_LOGIC;
  signal msg_block_in_IBUF_54 : STD_LOGIC;
  signal msg_block_in_IBUF_55 : STD_LOGIC;
  signal msg_block_in_IBUF_56 : STD_LOGIC;
  signal msg_block_in_IBUF_57 : STD_LOGIC;
  signal msg_block_in_IBUF_58 : STD_LOGIC;
  signal msg_block_in_IBUF_59 : STD_LOGIC;
  signal msg_block_in_IBUF_60 : STD_LOGIC;
  signal msg_block_in_IBUF_61 : STD_LOGIC;
  signal msg_block_in_IBUF_62 : STD_LOGIC;
  signal msg_block_in_IBUF_63 : STD_LOGIC;
  signal msg_block_in_IBUF_64 : STD_LOGIC;
  signal msg_block_in_IBUF_65 : STD_LOGIC;
  signal msg_block_in_IBUF_66 : STD_LOGIC;
  signal msg_block_in_IBUF_67 : STD_LOGIC;
  signal msg_block_in_IBUF_68 : STD_LOGIC;
  signal msg_block_in_IBUF_69 : STD_LOGIC;
  signal msg_block_in_IBUF_70 : STD_LOGIC;
  signal msg_block_in_IBUF_71 : STD_LOGIC;
  signal msg_block_in_IBUF_72 : STD_LOGIC;
  signal msg_block_in_IBUF_73 : STD_LOGIC;
  signal msg_block_in_IBUF_74 : STD_LOGIC;
  signal msg_block_in_IBUF_75 : STD_LOGIC;
  signal msg_block_in_IBUF_76 : STD_LOGIC;
  signal msg_block_in_IBUF_77 : STD_LOGIC;
  signal msg_block_in_IBUF_78 : STD_LOGIC;
  signal msg_block_in_IBUF_79 : STD_LOGIC;
  signal msg_block_in_IBUF_80 : STD_LOGIC;
  signal msg_block_in_IBUF_81 : STD_LOGIC;
  signal msg_block_in_IBUF_82 : STD_LOGIC;
  signal msg_block_in_IBUF_83 : STD_LOGIC;
  signal msg_block_in_IBUF_84 : STD_LOGIC;
  signal msg_block_in_IBUF_85 : STD_LOGIC;
  signal msg_block_in_IBUF_86 : STD_LOGIC;
  signal msg_block_in_IBUF_87 : STD_LOGIC;
  signal msg_block_in_IBUF_88 : STD_LOGIC;
  signal msg_block_in_IBUF_89 : STD_LOGIC;
  signal msg_block_in_IBUF_90 : STD_LOGIC;
  signal msg_block_in_IBUF_91 : STD_LOGIC;
  signal msg_block_in_IBUF_92 : STD_LOGIC;
  signal msg_block_in_IBUF_93 : STD_LOGIC;
  signal msg_block_in_IBUF_94 : STD_LOGIC;
  signal msg_block_in_IBUF_95 : STD_LOGIC;
  signal msg_block_in_IBUF_96 : STD_LOGIC;
  signal msg_block_in_IBUF_97 : STD_LOGIC;
  signal msg_block_in_IBUF_98 : STD_LOGIC;
  signal msg_block_in_IBUF_99 : STD_LOGIC;
  signal msg_block_in_IBUF_100 : STD_LOGIC;
  signal msg_block_in_IBUF_101 : STD_LOGIC;
  signal msg_block_in_IBUF_102 : STD_LOGIC;
  signal msg_block_in_IBUF_103 : STD_LOGIC;
  signal msg_block_in_IBUF_104 : STD_LOGIC;
  signal msg_block_in_IBUF_105 : STD_LOGIC;
  signal msg_block_in_IBUF_106 : STD_LOGIC;
  signal msg_block_in_IBUF_107 : STD_LOGIC;
  signal msg_block_in_IBUF_108 : STD_LOGIC;
  signal msg_block_in_IBUF_109 : STD_LOGIC;
  signal msg_block_in_IBUF_110 : STD_LOGIC;
  signal msg_block_in_IBUF_111 : STD_LOGIC;
  signal msg_block_in_IBUF_112 : STD_LOGIC;
  signal msg_block_in_IBUF_113 : STD_LOGIC;
  signal msg_block_in_IBUF_114 : STD_LOGIC;
  signal msg_block_in_IBUF_115 : STD_LOGIC;
  signal msg_block_in_IBUF_116 : STD_LOGIC;
  signal msg_block_in_IBUF_117 : STD_LOGIC;
  signal msg_block_in_IBUF_118 : STD_LOGIC;
  signal msg_block_in_IBUF_119 : STD_LOGIC;
  signal msg_block_in_IBUF_120 : STD_LOGIC;
  signal msg_block_in_IBUF_121 : STD_LOGIC;
  signal msg_block_in_IBUF_122 : STD_LOGIC;
  signal msg_block_in_IBUF_123 : STD_LOGIC;
  signal msg_block_in_IBUF_124 : STD_LOGIC;
  signal msg_block_in_IBUF_125 : STD_LOGIC;
  signal msg_block_in_IBUF_126 : STD_LOGIC;
  signal msg_block_in_IBUF_127 : STD_LOGIC;
  signal msg_block_in_IBUF_128 : STD_LOGIC;
  signal msg_block_in_IBUF_129 : STD_LOGIC;
  signal msg_block_in_IBUF_130 : STD_LOGIC;
  signal msg_block_in_IBUF_131 : STD_LOGIC;
  signal msg_block_in_IBUF_132 : STD_LOGIC;
  signal msg_block_in_IBUF_133 : STD_LOGIC;
  signal msg_block_in_IBUF_134 : STD_LOGIC;
  signal msg_block_in_IBUF_135 : STD_LOGIC;
  signal msg_block_in_IBUF_136 : STD_LOGIC;
  signal msg_block_in_IBUF_137 : STD_LOGIC;
  signal msg_block_in_IBUF_138 : STD_LOGIC;
  signal msg_block_in_IBUF_139 : STD_LOGIC;
  signal msg_block_in_IBUF_140 : STD_LOGIC;
  signal msg_block_in_IBUF_141 : STD_LOGIC;
  signal msg_block_in_IBUF_142 : STD_LOGIC;
  signal msg_block_in_IBUF_143 : STD_LOGIC;
  signal msg_block_in_IBUF_144 : STD_LOGIC;
  signal msg_block_in_IBUF_145 : STD_LOGIC;
  signal msg_block_in_IBUF_146 : STD_LOGIC;
  signal msg_block_in_IBUF_147 : STD_LOGIC;
  signal msg_block_in_IBUF_148 : STD_LOGIC;
  signal msg_block_in_IBUF_149 : STD_LOGIC;
  signal msg_block_in_IBUF_150 : STD_LOGIC;
  signal msg_block_in_IBUF_151 : STD_LOGIC;
  signal msg_block_in_IBUF_152 : STD_LOGIC;
  signal msg_block_in_IBUF_153 : STD_LOGIC;
  signal msg_block_in_IBUF_154 : STD_LOGIC;
  signal msg_block_in_IBUF_155 : STD_LOGIC;
  signal msg_block_in_IBUF_156 : STD_LOGIC;
  signal msg_block_in_IBUF_157 : STD_LOGIC;
  signal msg_block_in_IBUF_158 : STD_LOGIC;
  signal msg_block_in_IBUF_159 : STD_LOGIC;
  signal msg_block_in_IBUF_160 : STD_LOGIC;
  signal msg_block_in_IBUF_161 : STD_LOGIC;
  signal msg_block_in_IBUF_162 : STD_LOGIC;
  signal msg_block_in_IBUF_163 : STD_LOGIC;
  signal msg_block_in_IBUF_164 : STD_LOGIC;
  signal msg_block_in_IBUF_165 : STD_LOGIC;
  signal msg_block_in_IBUF_166 : STD_LOGIC;
  signal msg_block_in_IBUF_167 : STD_LOGIC;
  signal msg_block_in_IBUF_168 : STD_LOGIC;
  signal msg_block_in_IBUF_169 : STD_LOGIC;
  signal msg_block_in_IBUF_170 : STD_LOGIC;
  signal msg_block_in_IBUF_171 : STD_LOGIC;
  signal msg_block_in_IBUF_172 : STD_LOGIC;
  signal msg_block_in_IBUF_173 : STD_LOGIC;
  signal msg_block_in_IBUF_174 : STD_LOGIC;
  signal msg_block_in_IBUF_175 : STD_LOGIC;
  signal msg_block_in_IBUF_176 : STD_LOGIC;
  signal msg_block_in_IBUF_177 : STD_LOGIC;
  signal msg_block_in_IBUF_178 : STD_LOGIC;
  signal msg_block_in_IBUF_179 : STD_LOGIC;
  signal msg_block_in_IBUF_180 : STD_LOGIC;
  signal msg_block_in_IBUF_181 : STD_LOGIC;
  signal msg_block_in_IBUF_182 : STD_LOGIC;
  signal msg_block_in_IBUF_183 : STD_LOGIC;
  signal msg_block_in_IBUF_184 : STD_LOGIC;
  signal msg_block_in_IBUF_185 : STD_LOGIC;
  signal msg_block_in_IBUF_186 : STD_LOGIC;
  signal msg_block_in_IBUF_187 : STD_LOGIC;
  signal msg_block_in_IBUF_188 : STD_LOGIC;
  signal msg_block_in_IBUF_189 : STD_LOGIC;
  signal msg_block_in_IBUF_190 : STD_LOGIC;
  signal msg_block_in_IBUF_191 : STD_LOGIC;
  signal msg_block_in_IBUF_192 : STD_LOGIC;
  signal msg_block_in_IBUF_193 : STD_LOGIC;
  signal msg_block_in_IBUF_194 : STD_LOGIC;
  signal msg_block_in_IBUF_195 : STD_LOGIC;
  signal msg_block_in_IBUF_196 : STD_LOGIC;
  signal msg_block_in_IBUF_197 : STD_LOGIC;
  signal msg_block_in_IBUF_198 : STD_LOGIC;
  signal msg_block_in_IBUF_199 : STD_LOGIC;
  signal msg_block_in_IBUF_200 : STD_LOGIC;
  signal msg_block_in_IBUF_201 : STD_LOGIC;
  signal msg_block_in_IBUF_202 : STD_LOGIC;
  signal msg_block_in_IBUF_203 : STD_LOGIC;
  signal msg_block_in_IBUF_204 : STD_LOGIC;
  signal msg_block_in_IBUF_205 : STD_LOGIC;
  signal msg_block_in_IBUF_206 : STD_LOGIC;
  signal msg_block_in_IBUF_207 : STD_LOGIC;
  signal msg_block_in_IBUF_208 : STD_LOGIC;
  signal msg_block_in_IBUF_209 : STD_LOGIC;
  signal msg_block_in_IBUF_210 : STD_LOGIC;
  signal msg_block_in_IBUF_211 : STD_LOGIC;
  signal msg_block_in_IBUF_212 : STD_LOGIC;
  signal msg_block_in_IBUF_213 : STD_LOGIC;
  signal msg_block_in_IBUF_214 : STD_LOGIC;
  signal msg_block_in_IBUF_215 : STD_LOGIC;
  signal msg_block_in_IBUF_216 : STD_LOGIC;
  signal msg_block_in_IBUF_217 : STD_LOGIC;
  signal msg_block_in_IBUF_218 : STD_LOGIC;
  signal msg_block_in_IBUF_219 : STD_LOGIC;
  signal msg_block_in_IBUF_220 : STD_LOGIC;
  signal msg_block_in_IBUF_221 : STD_LOGIC;
  signal msg_block_in_IBUF_222 : STD_LOGIC;
  signal msg_block_in_IBUF_223 : STD_LOGIC;
  signal msg_block_in_IBUF_224 : STD_LOGIC;
  signal msg_block_in_IBUF_225 : STD_LOGIC;
  signal msg_block_in_IBUF_226 : STD_LOGIC;
  signal msg_block_in_IBUF_227 : STD_LOGIC;
  signal msg_block_in_IBUF_228 : STD_LOGIC;
  signal msg_block_in_IBUF_229 : STD_LOGIC;
  signal msg_block_in_IBUF_230 : STD_LOGIC;
  signal msg_block_in_IBUF_231 : STD_LOGIC;
  signal msg_block_in_IBUF_232 : STD_LOGIC;
  signal msg_block_in_IBUF_233 : STD_LOGIC;
  signal msg_block_in_IBUF_234 : STD_LOGIC;
  signal msg_block_in_IBUF_235 : STD_LOGIC;
  signal msg_block_in_IBUF_236 : STD_LOGIC;
  signal msg_block_in_IBUF_237 : STD_LOGIC;
  signal msg_block_in_IBUF_238 : STD_LOGIC;
  signal msg_block_in_IBUF_239 : STD_LOGIC;
  signal msg_block_in_IBUF_240 : STD_LOGIC;
  signal msg_block_in_IBUF_241 : STD_LOGIC;
  signal msg_block_in_IBUF_242 : STD_LOGIC;
  signal msg_block_in_IBUF_243 : STD_LOGIC;
  signal msg_block_in_IBUF_244 : STD_LOGIC;
  signal msg_block_in_IBUF_245 : STD_LOGIC;
  signal msg_block_in_IBUF_246 : STD_LOGIC;
  signal msg_block_in_IBUF_247 : STD_LOGIC;
  signal msg_block_in_IBUF_248 : STD_LOGIC;
  signal msg_block_in_IBUF_249 : STD_LOGIC;
  signal msg_block_in_IBUF_250 : STD_LOGIC;
  signal msg_block_in_IBUF_251 : STD_LOGIC;
  signal msg_block_in_IBUF_252 : STD_LOGIC;
  signal msg_block_in_IBUF_253 : STD_LOGIC;
  signal msg_block_in_IBUF_254 : STD_LOGIC;
  signal msg_block_in_IBUF_255 : STD_LOGIC;
  signal msg_block_in_IBUF_256 : STD_LOGIC;
  signal msg_block_in_IBUF_257 : STD_LOGIC;
  signal msg_block_in_IBUF_258 : STD_LOGIC;
  signal msg_block_in_IBUF_259 : STD_LOGIC;
  signal msg_block_in_IBUF_260 : STD_LOGIC;
  signal msg_block_in_IBUF_261 : STD_LOGIC;
  signal msg_block_in_IBUF_262 : STD_LOGIC;
  signal msg_block_in_IBUF_263 : STD_LOGIC;
  signal msg_block_in_IBUF_264 : STD_LOGIC;
  signal msg_block_in_IBUF_265 : STD_LOGIC;
  signal msg_block_in_IBUF_266 : STD_LOGIC;
  signal msg_block_in_IBUF_267 : STD_LOGIC;
  signal msg_block_in_IBUF_268 : STD_LOGIC;
  signal msg_block_in_IBUF_269 : STD_LOGIC;
  signal msg_block_in_IBUF_270 : STD_LOGIC;
  signal msg_block_in_IBUF_271 : STD_LOGIC;
  signal msg_block_in_IBUF_272 : STD_LOGIC;
  signal msg_block_in_IBUF_273 : STD_LOGIC;
  signal msg_block_in_IBUF_274 : STD_LOGIC;
  signal msg_block_in_IBUF_275 : STD_LOGIC;
  signal msg_block_in_IBUF_276 : STD_LOGIC;
  signal msg_block_in_IBUF_277 : STD_LOGIC;
  signal msg_block_in_IBUF_278 : STD_LOGIC;
  signal msg_block_in_IBUF_279 : STD_LOGIC;
  signal msg_block_in_IBUF_280 : STD_LOGIC;
  signal msg_block_in_IBUF_281 : STD_LOGIC;
  signal msg_block_in_IBUF_282 : STD_LOGIC;
  signal msg_block_in_IBUF_283 : STD_LOGIC;
  signal msg_block_in_IBUF_284 : STD_LOGIC;
  signal msg_block_in_IBUF_285 : STD_LOGIC;
  signal msg_block_in_IBUF_286 : STD_LOGIC;
  signal msg_block_in_IBUF_287 : STD_LOGIC;
  signal msg_block_in_IBUF_288 : STD_LOGIC;
  signal msg_block_in_IBUF_289 : STD_LOGIC;
  signal msg_block_in_IBUF_290 : STD_LOGIC;
  signal msg_block_in_IBUF_291 : STD_LOGIC;
  signal msg_block_in_IBUF_292 : STD_LOGIC;
  signal msg_block_in_IBUF_293 : STD_LOGIC;
  signal msg_block_in_IBUF_294 : STD_LOGIC;
  signal msg_block_in_IBUF_295 : STD_LOGIC;
  signal msg_block_in_IBUF_296 : STD_LOGIC;
  signal msg_block_in_IBUF_297 : STD_LOGIC;
  signal msg_block_in_IBUF_298 : STD_LOGIC;
  signal msg_block_in_IBUF_299 : STD_LOGIC;
  signal msg_block_in_IBUF_300 : STD_LOGIC;
  signal msg_block_in_IBUF_301 : STD_LOGIC;
  signal msg_block_in_IBUF_302 : STD_LOGIC;
  signal msg_block_in_IBUF_303 : STD_LOGIC;
  signal msg_block_in_IBUF_304 : STD_LOGIC;
  signal msg_block_in_IBUF_305 : STD_LOGIC;
  signal msg_block_in_IBUF_306 : STD_LOGIC;
  signal msg_block_in_IBUF_307 : STD_LOGIC;
  signal msg_block_in_IBUF_308 : STD_LOGIC;
  signal msg_block_in_IBUF_309 : STD_LOGIC;
  signal msg_block_in_IBUF_310 : STD_LOGIC;
  signal msg_block_in_IBUF_311 : STD_LOGIC;
  signal msg_block_in_IBUF_312 : STD_LOGIC;
  signal msg_block_in_IBUF_313 : STD_LOGIC;
  signal msg_block_in_IBUF_314 : STD_LOGIC;
  signal msg_block_in_IBUF_315 : STD_LOGIC;
  signal msg_block_in_IBUF_316 : STD_LOGIC;
  signal msg_block_in_IBUF_317 : STD_LOGIC;
  signal msg_block_in_IBUF_318 : STD_LOGIC;
  signal msg_block_in_IBUF_319 : STD_LOGIC;
  signal msg_block_in_IBUF_320 : STD_LOGIC;
  signal msg_block_in_IBUF_321 : STD_LOGIC;
  signal msg_block_in_IBUF_322 : STD_LOGIC;
  signal msg_block_in_IBUF_323 : STD_LOGIC;
  signal msg_block_in_IBUF_324 : STD_LOGIC;
  signal msg_block_in_IBUF_325 : STD_LOGIC;
  signal msg_block_in_IBUF_326 : STD_LOGIC;
  signal msg_block_in_IBUF_327 : STD_LOGIC;
  signal msg_block_in_IBUF_328 : STD_LOGIC;
  signal msg_block_in_IBUF_329 : STD_LOGIC;
  signal msg_block_in_IBUF_330 : STD_LOGIC;
  signal msg_block_in_IBUF_331 : STD_LOGIC;
  signal msg_block_in_IBUF_332 : STD_LOGIC;
  signal msg_block_in_IBUF_333 : STD_LOGIC;
  signal msg_block_in_IBUF_334 : STD_LOGIC;
  signal msg_block_in_IBUF_335 : STD_LOGIC;
  signal msg_block_in_IBUF_336 : STD_LOGIC;
  signal msg_block_in_IBUF_337 : STD_LOGIC;
  signal msg_block_in_IBUF_338 : STD_LOGIC;
  signal msg_block_in_IBUF_339 : STD_LOGIC;
  signal msg_block_in_IBUF_340 : STD_LOGIC;
  signal msg_block_in_IBUF_341 : STD_LOGIC;
  signal msg_block_in_IBUF_342 : STD_LOGIC;
  signal msg_block_in_IBUF_343 : STD_LOGIC;
  signal msg_block_in_IBUF_344 : STD_LOGIC;
  signal msg_block_in_IBUF_345 : STD_LOGIC;
  signal msg_block_in_IBUF_346 : STD_LOGIC;
  signal msg_block_in_IBUF_347 : STD_LOGIC;
  signal msg_block_in_IBUF_348 : STD_LOGIC;
  signal msg_block_in_IBUF_349 : STD_LOGIC;
  signal msg_block_in_IBUF_350 : STD_LOGIC;
  signal msg_block_in_IBUF_351 : STD_LOGIC;
  signal msg_block_in_IBUF_352 : STD_LOGIC;
  signal msg_block_in_IBUF_353 : STD_LOGIC;
  signal msg_block_in_IBUF_354 : STD_LOGIC;
  signal msg_block_in_IBUF_355 : STD_LOGIC;
  signal msg_block_in_IBUF_356 : STD_LOGIC;
  signal msg_block_in_IBUF_357 : STD_LOGIC;
  signal msg_block_in_IBUF_358 : STD_LOGIC;
  signal msg_block_in_IBUF_359 : STD_LOGIC;
  signal msg_block_in_IBUF_360 : STD_LOGIC;
  signal msg_block_in_IBUF_361 : STD_LOGIC;
  signal msg_block_in_IBUF_362 : STD_LOGIC;
  signal msg_block_in_IBUF_363 : STD_LOGIC;
  signal msg_block_in_IBUF_364 : STD_LOGIC;
  signal msg_block_in_IBUF_365 : STD_LOGIC;
  signal msg_block_in_IBUF_366 : STD_LOGIC;
  signal msg_block_in_IBUF_367 : STD_LOGIC;
  signal msg_block_in_IBUF_368 : STD_LOGIC;
  signal msg_block_in_IBUF_369 : STD_LOGIC;
  signal msg_block_in_IBUF_370 : STD_LOGIC;
  signal msg_block_in_IBUF_371 : STD_LOGIC;
  signal msg_block_in_IBUF_372 : STD_LOGIC;
  signal msg_block_in_IBUF_373 : STD_LOGIC;
  signal msg_block_in_IBUF_374 : STD_LOGIC;
  signal msg_block_in_IBUF_375 : STD_LOGIC;
  signal msg_block_in_IBUF_376 : STD_LOGIC;
  signal msg_block_in_IBUF_377 : STD_LOGIC;
  signal msg_block_in_IBUF_378 : STD_LOGIC;
  signal msg_block_in_IBUF_379 : STD_LOGIC;
  signal msg_block_in_IBUF_380 : STD_LOGIC;
  signal msg_block_in_IBUF_381 : STD_LOGIC;
  signal msg_block_in_IBUF_382 : STD_LOGIC;
  signal msg_block_in_IBUF_383 : STD_LOGIC;
  signal msg_block_in_IBUF_384 : STD_LOGIC;
  signal msg_block_in_IBUF_385 : STD_LOGIC;
  signal msg_block_in_IBUF_386 : STD_LOGIC;
  signal msg_block_in_IBUF_387 : STD_LOGIC;
  signal msg_block_in_IBUF_388 : STD_LOGIC;
  signal msg_block_in_IBUF_389 : STD_LOGIC;
  signal msg_block_in_IBUF_390 : STD_LOGIC;
  signal msg_block_in_IBUF_391 : STD_LOGIC;
  signal msg_block_in_IBUF_392 : STD_LOGIC;
  signal msg_block_in_IBUF_393 : STD_LOGIC;
  signal msg_block_in_IBUF_394 : STD_LOGIC;
  signal msg_block_in_IBUF_395 : STD_LOGIC;
  signal msg_block_in_IBUF_396 : STD_LOGIC;
  signal msg_block_in_IBUF_397 : STD_LOGIC;
  signal msg_block_in_IBUF_398 : STD_LOGIC;
  signal msg_block_in_IBUF_399 : STD_LOGIC;
  signal msg_block_in_IBUF_400 : STD_LOGIC;
  signal msg_block_in_IBUF_401 : STD_LOGIC;
  signal msg_block_in_IBUF_402 : STD_LOGIC;
  signal msg_block_in_IBUF_403 : STD_LOGIC;
  signal msg_block_in_IBUF_404 : STD_LOGIC;
  signal msg_block_in_IBUF_405 : STD_LOGIC;
  signal msg_block_in_IBUF_406 : STD_LOGIC;
  signal msg_block_in_IBUF_407 : STD_LOGIC;
  signal msg_block_in_IBUF_408 : STD_LOGIC;
  signal msg_block_in_IBUF_409 : STD_LOGIC;
  signal msg_block_in_IBUF_410 : STD_LOGIC;
  signal msg_block_in_IBUF_411 : STD_LOGIC;
  signal msg_block_in_IBUF_412 : STD_LOGIC;
  signal msg_block_in_IBUF_413 : STD_LOGIC;
  signal msg_block_in_IBUF_414 : STD_LOGIC;
  signal msg_block_in_IBUF_415 : STD_LOGIC;
  signal msg_block_in_IBUF_416 : STD_LOGIC;
  signal msg_block_in_IBUF_417 : STD_LOGIC;
  signal msg_block_in_IBUF_418 : STD_LOGIC;
  signal msg_block_in_IBUF_419 : STD_LOGIC;
  signal msg_block_in_IBUF_420 : STD_LOGIC;
  signal msg_block_in_IBUF_421 : STD_LOGIC;
  signal msg_block_in_IBUF_422 : STD_LOGIC;
  signal msg_block_in_IBUF_423 : STD_LOGIC;
  signal msg_block_in_IBUF_424 : STD_LOGIC;
  signal msg_block_in_IBUF_425 : STD_LOGIC;
  signal msg_block_in_IBUF_426 : STD_LOGIC;
  signal msg_block_in_IBUF_427 : STD_LOGIC;
  signal msg_block_in_IBUF_428 : STD_LOGIC;
  signal msg_block_in_IBUF_429 : STD_LOGIC;
  signal msg_block_in_IBUF_430 : STD_LOGIC;
  signal msg_block_in_IBUF_431 : STD_LOGIC;
  signal msg_block_in_IBUF_432 : STD_LOGIC;
  signal msg_block_in_IBUF_433 : STD_LOGIC;
  signal msg_block_in_IBUF_434 : STD_LOGIC;
  signal msg_block_in_IBUF_435 : STD_LOGIC;
  signal msg_block_in_IBUF_436 : STD_LOGIC;
  signal msg_block_in_IBUF_437 : STD_LOGIC;
  signal msg_block_in_IBUF_438 : STD_LOGIC;
  signal msg_block_in_IBUF_439 : STD_LOGIC;
  signal msg_block_in_IBUF_440 : STD_LOGIC;
  signal msg_block_in_IBUF_441 : STD_LOGIC;
  signal msg_block_in_IBUF_442 : STD_LOGIC;
  signal msg_block_in_IBUF_443 : STD_LOGIC;
  signal msg_block_in_IBUF_444 : STD_LOGIC;
  signal msg_block_in_IBUF_445 : STD_LOGIC;
  signal msg_block_in_IBUF_446 : STD_LOGIC;
  signal msg_block_in_IBUF_447 : STD_LOGIC;
  signal msg_block_in_IBUF_448 : STD_LOGIC;
  signal msg_block_in_IBUF_449 : STD_LOGIC;
  signal msg_block_in_IBUF_450 : STD_LOGIC;
  signal msg_block_in_IBUF_451 : STD_LOGIC;
  signal msg_block_in_IBUF_452 : STD_LOGIC;
  signal msg_block_in_IBUF_453 : STD_LOGIC;
  signal msg_block_in_IBUF_454 : STD_LOGIC;
  signal msg_block_in_IBUF_455 : STD_LOGIC;
  signal msg_block_in_IBUF_456 : STD_LOGIC;
  signal msg_block_in_IBUF_457 : STD_LOGIC;
  signal msg_block_in_IBUF_458 : STD_LOGIC;
  signal msg_block_in_IBUF_459 : STD_LOGIC;
  signal msg_block_in_IBUF_460 : STD_LOGIC;
  signal msg_block_in_IBUF_461 : STD_LOGIC;
  signal msg_block_in_IBUF_462 : STD_LOGIC;
  signal msg_block_in_IBUF_463 : STD_LOGIC;
  signal msg_block_in_IBUF_464 : STD_LOGIC;
  signal msg_block_in_IBUF_465 : STD_LOGIC;
  signal msg_block_in_IBUF_466 : STD_LOGIC;
  signal msg_block_in_IBUF_467 : STD_LOGIC;
  signal msg_block_in_IBUF_468 : STD_LOGIC;
  signal msg_block_in_IBUF_469 : STD_LOGIC;
  signal msg_block_in_IBUF_470 : STD_LOGIC;
  signal msg_block_in_IBUF_471 : STD_LOGIC;
  signal msg_block_in_IBUF_472 : STD_LOGIC;
  signal msg_block_in_IBUF_473 : STD_LOGIC;
  signal msg_block_in_IBUF_474 : STD_LOGIC;
  signal msg_block_in_IBUF_475 : STD_LOGIC;
  signal msg_block_in_IBUF_476 : STD_LOGIC;
  signal msg_block_in_IBUF_477 : STD_LOGIC;
  signal msg_block_in_IBUF_478 : STD_LOGIC;
  signal msg_block_in_IBUF_479 : STD_LOGIC;
  signal msg_block_in_IBUF_480 : STD_LOGIC;
  signal msg_block_in_IBUF_481 : STD_LOGIC;
  signal msg_block_in_IBUF_482 : STD_LOGIC;
  signal msg_block_in_IBUF_483 : STD_LOGIC;
  signal msg_block_in_IBUF_484 : STD_LOGIC;
  signal msg_block_in_IBUF_485 : STD_LOGIC;
  signal msg_block_in_IBUF_486 : STD_LOGIC;
  signal msg_block_in_IBUF_487 : STD_LOGIC;
  signal msg_block_in_IBUF_488 : STD_LOGIC;
  signal msg_block_in_IBUF_489 : STD_LOGIC;
  signal msg_block_in_IBUF_490 : STD_LOGIC;
  signal msg_block_in_IBUF_491 : STD_LOGIC;
  signal msg_block_in_IBUF_492 : STD_LOGIC;
  signal msg_block_in_IBUF_493 : STD_LOGIC;
  signal msg_block_in_IBUF_494 : STD_LOGIC;
  signal msg_block_in_IBUF_495 : STD_LOGIC;
  signal msg_block_in_IBUF_496 : STD_LOGIC;
  signal msg_block_in_IBUF_497 : STD_LOGIC;
  signal msg_block_in_IBUF_498 : STD_LOGIC;
  signal msg_block_in_IBUF_499 : STD_LOGIC;
  signal msg_block_in_IBUF_500 : STD_LOGIC;
  signal msg_block_in_IBUF_501 : STD_LOGIC;
  signal msg_block_in_IBUF_502 : STD_LOGIC;
  signal msg_block_in_IBUF_503 : STD_LOGIC;
  signal msg_block_in_IBUF_504 : STD_LOGIC;
  signal msg_block_in_IBUF_505 : STD_LOGIC;
  signal msg_block_in_IBUF_506 : STD_LOGIC;
  signal msg_block_in_IBUF_507 : STD_LOGIC;
  signal msg_block_in_IBUF_508 : STD_LOGIC;
  signal msg_block_in_IBUF_509 : STD_LOGIC;
  signal msg_block_in_IBUF_510 : STD_LOGIC;
  signal msg_block_in_IBUF_511 : STD_LOGIC;
  signal M_0 : STD_LOGIC;
  signal M_reg_0_31 : STD_LOGIC;
  signal M_reg_0_30 : STD_LOGIC;
  signal M_reg_0_29 : STD_LOGIC;
  signal M_reg_0_28 : STD_LOGIC;
  signal M_reg_0_27 : STD_LOGIC;
  signal M_reg_0_26 : STD_LOGIC;
  signal M_reg_0_25 : STD_LOGIC;
  signal M_reg_0_24 : STD_LOGIC;
  signal M_reg_0_23 : STD_LOGIC;
  signal M_reg_0_22 : STD_LOGIC;
  signal M_reg_0_21 : STD_LOGIC;
  signal M_reg_0_20 : STD_LOGIC;
  signal M_reg_0_19 : STD_LOGIC;
  signal M_reg_0_18 : STD_LOGIC;
  signal M_reg_0_17 : STD_LOGIC;
  signal M_reg_0_16 : STD_LOGIC;
  signal M_reg_0_15 : STD_LOGIC;
  signal M_reg_0_14 : STD_LOGIC;
  signal M_reg_0_13 : STD_LOGIC;
  signal M_reg_0_12 : STD_LOGIC;
  signal M_reg_0_11 : STD_LOGIC;
  signal M_reg_0_10 : STD_LOGIC;
  signal M_reg_0_9 : STD_LOGIC;
  signal M_reg_0_8 : STD_LOGIC;
  signal M_reg_0_7 : STD_LOGIC;
  signal M_reg_0_6 : STD_LOGIC;
  signal M_reg_0_5 : STD_LOGIC;
  signal M_reg_0_4 : STD_LOGIC;
  signal M_reg_0_3 : STD_LOGIC;
  signal M_reg_0_2 : STD_LOGIC;
  signal M_reg_0_1 : STD_LOGIC;
  signal M_reg_0_0 : STD_LOGIC;
  signal M_reg_10_31 : STD_LOGIC;
  signal M_reg_10_30 : STD_LOGIC;
  signal M_reg_10_29 : STD_LOGIC;
  signal M_reg_10_28 : STD_LOGIC;
  signal M_reg_10_27 : STD_LOGIC;
  signal M_reg_10_26 : STD_LOGIC;
  signal M_reg_10_25 : STD_LOGIC;
  signal M_reg_10_24 : STD_LOGIC;
  signal M_reg_10_23 : STD_LOGIC;
  signal M_reg_10_22 : STD_LOGIC;
  signal M_reg_10_21 : STD_LOGIC;
  signal M_reg_10_20 : STD_LOGIC;
  signal M_reg_10_19 : STD_LOGIC;
  signal M_reg_10_18 : STD_LOGIC;
  signal M_reg_10_17 : STD_LOGIC;
  signal M_reg_10_16 : STD_LOGIC;
  signal M_reg_10_15 : STD_LOGIC;
  signal M_reg_10_14 : STD_LOGIC;
  signal M_reg_10_13 : STD_LOGIC;
  signal M_reg_10_12 : STD_LOGIC;
  signal M_reg_10_11 : STD_LOGIC;
  signal M_reg_10_10 : STD_LOGIC;
  signal M_reg_10_9 : STD_LOGIC;
  signal M_reg_10_8 : STD_LOGIC;
  signal M_reg_10_7 : STD_LOGIC;
  signal M_reg_10_6 : STD_LOGIC;
  signal M_reg_10_5 : STD_LOGIC;
  signal M_reg_10_4 : STD_LOGIC;
  signal M_reg_10_3 : STD_LOGIC;
  signal M_reg_10_2 : STD_LOGIC;
  signal M_reg_10_1 : STD_LOGIC;
  signal M_reg_10_0 : STD_LOGIC;
  signal M_reg_11_31 : STD_LOGIC;
  signal M_reg_11_30 : STD_LOGIC;
  signal M_reg_11_29 : STD_LOGIC;
  signal M_reg_11_28 : STD_LOGIC;
  signal M_reg_11_27 : STD_LOGIC;
  signal M_reg_11_26 : STD_LOGIC;
  signal M_reg_11_25 : STD_LOGIC;
  signal M_reg_11_24 : STD_LOGIC;
  signal M_reg_11_23 : STD_LOGIC;
  signal M_reg_11_22 : STD_LOGIC;
  signal M_reg_11_21 : STD_LOGIC;
  signal M_reg_11_20 : STD_LOGIC;
  signal M_reg_11_19 : STD_LOGIC;
  signal M_reg_11_18 : STD_LOGIC;
  signal M_reg_11_17 : STD_LOGIC;
  signal M_reg_11_16 : STD_LOGIC;
  signal M_reg_11_15 : STD_LOGIC;
  signal M_reg_11_14 : STD_LOGIC;
  signal M_reg_11_13 : STD_LOGIC;
  signal M_reg_11_12 : STD_LOGIC;
  signal M_reg_11_11 : STD_LOGIC;
  signal M_reg_11_10 : STD_LOGIC;
  signal M_reg_11_9 : STD_LOGIC;
  signal M_reg_11_8 : STD_LOGIC;
  signal M_reg_11_7 : STD_LOGIC;
  signal M_reg_11_6 : STD_LOGIC;
  signal M_reg_11_5 : STD_LOGIC;
  signal M_reg_11_4 : STD_LOGIC;
  signal M_reg_11_3 : STD_LOGIC;
  signal M_reg_11_2 : STD_LOGIC;
  signal M_reg_11_1 : STD_LOGIC;
  signal M_reg_11_0 : STD_LOGIC;
  signal M_reg_12_31 : STD_LOGIC;
  signal M_reg_12_30 : STD_LOGIC;
  signal M_reg_12_29 : STD_LOGIC;
  signal M_reg_12_28 : STD_LOGIC;
  signal M_reg_12_27 : STD_LOGIC;
  signal M_reg_12_26 : STD_LOGIC;
  signal M_reg_12_25 : STD_LOGIC;
  signal M_reg_12_24 : STD_LOGIC;
  signal M_reg_12_23 : STD_LOGIC;
  signal M_reg_12_22 : STD_LOGIC;
  signal M_reg_12_21 : STD_LOGIC;
  signal M_reg_12_20 : STD_LOGIC;
  signal M_reg_12_19 : STD_LOGIC;
  signal M_reg_12_18 : STD_LOGIC;
  signal M_reg_12_17 : STD_LOGIC;
  signal M_reg_12_16 : STD_LOGIC;
  signal M_reg_12_15 : STD_LOGIC;
  signal M_reg_12_14 : STD_LOGIC;
  signal M_reg_12_13 : STD_LOGIC;
  signal M_reg_12_12 : STD_LOGIC;
  signal M_reg_12_11 : STD_LOGIC;
  signal M_reg_12_10 : STD_LOGIC;
  signal M_reg_12_9 : STD_LOGIC;
  signal M_reg_12_8 : STD_LOGIC;
  signal M_reg_12_7 : STD_LOGIC;
  signal M_reg_12_6 : STD_LOGIC;
  signal M_reg_12_5 : STD_LOGIC;
  signal M_reg_12_4 : STD_LOGIC;
  signal M_reg_12_3 : STD_LOGIC;
  signal M_reg_12_2 : STD_LOGIC;
  signal M_reg_12_1 : STD_LOGIC;
  signal M_reg_12_0 : STD_LOGIC;
  signal M_reg_13_31 : STD_LOGIC;
  signal M_reg_13_30 : STD_LOGIC;
  signal M_reg_13_29 : STD_LOGIC;
  signal M_reg_13_28 : STD_LOGIC;
  signal M_reg_13_27 : STD_LOGIC;
  signal M_reg_13_26 : STD_LOGIC;
  signal M_reg_13_25 : STD_LOGIC;
  signal M_reg_13_24 : STD_LOGIC;
  signal M_reg_13_23 : STD_LOGIC;
  signal M_reg_13_22 : STD_LOGIC;
  signal M_reg_13_21 : STD_LOGIC;
  signal M_reg_13_20 : STD_LOGIC;
  signal M_reg_13_19 : STD_LOGIC;
  signal M_reg_13_18 : STD_LOGIC;
  signal M_reg_13_17 : STD_LOGIC;
  signal M_reg_13_16 : STD_LOGIC;
  signal M_reg_13_15 : STD_LOGIC;
  signal M_reg_13_14 : STD_LOGIC;
  signal M_reg_13_13 : STD_LOGIC;
  signal M_reg_13_12 : STD_LOGIC;
  signal M_reg_13_11 : STD_LOGIC;
  signal M_reg_13_10 : STD_LOGIC;
  signal M_reg_13_9 : STD_LOGIC;
  signal M_reg_13_8 : STD_LOGIC;
  signal M_reg_13_7 : STD_LOGIC;
  signal M_reg_13_6 : STD_LOGIC;
  signal M_reg_13_5 : STD_LOGIC;
  signal M_reg_13_4 : STD_LOGIC;
  signal M_reg_13_3 : STD_LOGIC;
  signal M_reg_13_2 : STD_LOGIC;
  signal M_reg_13_1 : STD_LOGIC;
  signal M_reg_13_0 : STD_LOGIC;
  signal M_reg_14_31 : STD_LOGIC;
  signal M_reg_14_30 : STD_LOGIC;
  signal M_reg_14_29 : STD_LOGIC;
  signal M_reg_14_28 : STD_LOGIC;
  signal M_reg_14_27 : STD_LOGIC;
  signal M_reg_14_26 : STD_LOGIC;
  signal M_reg_14_25 : STD_LOGIC;
  signal M_reg_14_24 : STD_LOGIC;
  signal M_reg_14_23 : STD_LOGIC;
  signal M_reg_14_22 : STD_LOGIC;
  signal M_reg_14_21 : STD_LOGIC;
  signal M_reg_14_20 : STD_LOGIC;
  signal M_reg_14_19 : STD_LOGIC;
  signal M_reg_14_18 : STD_LOGIC;
  signal M_reg_14_17 : STD_LOGIC;
  signal M_reg_14_16 : STD_LOGIC;
  signal M_reg_14_15 : STD_LOGIC;
  signal M_reg_14_14 : STD_LOGIC;
  signal M_reg_14_13 : STD_LOGIC;
  signal M_reg_14_12 : STD_LOGIC;
  signal M_reg_14_11 : STD_LOGIC;
  signal M_reg_14_10 : STD_LOGIC;
  signal M_reg_14_9 : STD_LOGIC;
  signal M_reg_14_8 : STD_LOGIC;
  signal M_reg_14_7 : STD_LOGIC;
  signal M_reg_14_6 : STD_LOGIC;
  signal M_reg_14_5 : STD_LOGIC;
  signal M_reg_14_4 : STD_LOGIC;
  signal M_reg_14_3 : STD_LOGIC;
  signal M_reg_14_2 : STD_LOGIC;
  signal M_reg_14_1 : STD_LOGIC;
  signal M_reg_14_0 : STD_LOGIC;
  signal M_reg_15_31 : STD_LOGIC;
  signal M_reg_15_30 : STD_LOGIC;
  signal M_reg_15_29 : STD_LOGIC;
  signal M_reg_15_28 : STD_LOGIC;
  signal M_reg_15_27 : STD_LOGIC;
  signal M_reg_15_26 : STD_LOGIC;
  signal M_reg_15_25 : STD_LOGIC;
  signal M_reg_15_24 : STD_LOGIC;
  signal M_reg_15_23 : STD_LOGIC;
  signal M_reg_15_22 : STD_LOGIC;
  signal M_reg_15_21 : STD_LOGIC;
  signal M_reg_15_20 : STD_LOGIC;
  signal M_reg_15_19 : STD_LOGIC;
  signal M_reg_15_18 : STD_LOGIC;
  signal M_reg_15_17 : STD_LOGIC;
  signal M_reg_15_16 : STD_LOGIC;
  signal M_reg_15_15 : STD_LOGIC;
  signal M_reg_15_14 : STD_LOGIC;
  signal M_reg_15_13 : STD_LOGIC;
  signal M_reg_15_12 : STD_LOGIC;
  signal M_reg_15_11 : STD_LOGIC;
  signal M_reg_15_10 : STD_LOGIC;
  signal M_reg_15_9 : STD_LOGIC;
  signal M_reg_15_8 : STD_LOGIC;
  signal M_reg_15_7 : STD_LOGIC;
  signal M_reg_15_6 : STD_LOGIC;
  signal M_reg_15_5 : STD_LOGIC;
  signal M_reg_15_4 : STD_LOGIC;
  signal M_reg_15_3 : STD_LOGIC;
  signal M_reg_15_2 : STD_LOGIC;
  signal M_reg_15_1 : STD_LOGIC;
  signal M_reg_15_0 : STD_LOGIC;
  signal M_reg_1_31 : STD_LOGIC;
  signal M_reg_1_30 : STD_LOGIC;
  signal M_reg_1_29 : STD_LOGIC;
  signal M_reg_1_28 : STD_LOGIC;
  signal M_reg_1_27 : STD_LOGIC;
  signal M_reg_1_26 : STD_LOGIC;
  signal M_reg_1_25 : STD_LOGIC;
  signal M_reg_1_24 : STD_LOGIC;
  signal M_reg_1_23 : STD_LOGIC;
  signal M_reg_1_22 : STD_LOGIC;
  signal M_reg_1_21 : STD_LOGIC;
  signal M_reg_1_20 : STD_LOGIC;
  signal M_reg_1_19 : STD_LOGIC;
  signal M_reg_1_18 : STD_LOGIC;
  signal M_reg_1_17 : STD_LOGIC;
  signal M_reg_1_16 : STD_LOGIC;
  signal M_reg_1_15 : STD_LOGIC;
  signal M_reg_1_14 : STD_LOGIC;
  signal M_reg_1_13 : STD_LOGIC;
  signal M_reg_1_12 : STD_LOGIC;
  signal M_reg_1_11 : STD_LOGIC;
  signal M_reg_1_10 : STD_LOGIC;
  signal M_reg_1_9 : STD_LOGIC;
  signal M_reg_1_8 : STD_LOGIC;
  signal M_reg_1_7 : STD_LOGIC;
  signal M_reg_1_6 : STD_LOGIC;
  signal M_reg_1_5 : STD_LOGIC;
  signal M_reg_1_4 : STD_LOGIC;
  signal M_reg_1_3 : STD_LOGIC;
  signal M_reg_1_2 : STD_LOGIC;
  signal M_reg_1_1 : STD_LOGIC;
  signal M_reg_1_0 : STD_LOGIC;
  signal M_reg_2_31 : STD_LOGIC;
  signal M_reg_2_30 : STD_LOGIC;
  signal M_reg_2_29 : STD_LOGIC;
  signal M_reg_2_28 : STD_LOGIC;
  signal M_reg_2_27 : STD_LOGIC;
  signal M_reg_2_26 : STD_LOGIC;
  signal M_reg_2_25 : STD_LOGIC;
  signal M_reg_2_24 : STD_LOGIC;
  signal M_reg_2_23 : STD_LOGIC;
  signal M_reg_2_22 : STD_LOGIC;
  signal M_reg_2_21 : STD_LOGIC;
  signal M_reg_2_20 : STD_LOGIC;
  signal M_reg_2_19 : STD_LOGIC;
  signal M_reg_2_18 : STD_LOGIC;
  signal M_reg_2_17 : STD_LOGIC;
  signal M_reg_2_16 : STD_LOGIC;
  signal M_reg_2_15 : STD_LOGIC;
  signal M_reg_2_14 : STD_LOGIC;
  signal M_reg_2_13 : STD_LOGIC;
  signal M_reg_2_12 : STD_LOGIC;
  signal M_reg_2_11 : STD_LOGIC;
  signal M_reg_2_10 : STD_LOGIC;
  signal M_reg_2_9 : STD_LOGIC;
  signal M_reg_2_8 : STD_LOGIC;
  signal M_reg_2_7 : STD_LOGIC;
  signal M_reg_2_6 : STD_LOGIC;
  signal M_reg_2_5 : STD_LOGIC;
  signal M_reg_2_4 : STD_LOGIC;
  signal M_reg_2_3 : STD_LOGIC;
  signal M_reg_2_2 : STD_LOGIC;
  signal M_reg_2_1 : STD_LOGIC;
  signal M_reg_2_0 : STD_LOGIC;
  signal M_reg_3_31 : STD_LOGIC;
  signal M_reg_3_30 : STD_LOGIC;
  signal M_reg_3_29 : STD_LOGIC;
  signal M_reg_3_28 : STD_LOGIC;
  signal M_reg_3_27 : STD_LOGIC;
  signal M_reg_3_26 : STD_LOGIC;
  signal M_reg_3_25 : STD_LOGIC;
  signal M_reg_3_24 : STD_LOGIC;
  signal M_reg_3_23 : STD_LOGIC;
  signal M_reg_3_22 : STD_LOGIC;
  signal M_reg_3_21 : STD_LOGIC;
  signal M_reg_3_20 : STD_LOGIC;
  signal M_reg_3_19 : STD_LOGIC;
  signal M_reg_3_18 : STD_LOGIC;
  signal M_reg_3_17 : STD_LOGIC;
  signal M_reg_3_16 : STD_LOGIC;
  signal M_reg_3_15 : STD_LOGIC;
  signal M_reg_3_14 : STD_LOGIC;
  signal M_reg_3_13 : STD_LOGIC;
  signal M_reg_3_12 : STD_LOGIC;
  signal M_reg_3_11 : STD_LOGIC;
  signal M_reg_3_10 : STD_LOGIC;
  signal M_reg_3_9 : STD_LOGIC;
  signal M_reg_3_8 : STD_LOGIC;
  signal M_reg_3_7 : STD_LOGIC;
  signal M_reg_3_6 : STD_LOGIC;
  signal M_reg_3_5 : STD_LOGIC;
  signal M_reg_3_4 : STD_LOGIC;
  signal M_reg_3_3 : STD_LOGIC;
  signal M_reg_3_2 : STD_LOGIC;
  signal M_reg_3_1 : STD_LOGIC;
  signal M_reg_3_0 : STD_LOGIC;
  signal M_reg_4_31 : STD_LOGIC;
  signal M_reg_4_30 : STD_LOGIC;
  signal M_reg_4_29 : STD_LOGIC;
  signal M_reg_4_28 : STD_LOGIC;
  signal M_reg_4_27 : STD_LOGIC;
  signal M_reg_4_26 : STD_LOGIC;
  signal M_reg_4_25 : STD_LOGIC;
  signal M_reg_4_24 : STD_LOGIC;
  signal M_reg_4_23 : STD_LOGIC;
  signal M_reg_4_22 : STD_LOGIC;
  signal M_reg_4_21 : STD_LOGIC;
  signal M_reg_4_20 : STD_LOGIC;
  signal M_reg_4_19 : STD_LOGIC;
  signal M_reg_4_18 : STD_LOGIC;
  signal M_reg_4_17 : STD_LOGIC;
  signal M_reg_4_16 : STD_LOGIC;
  signal M_reg_4_15 : STD_LOGIC;
  signal M_reg_4_14 : STD_LOGIC;
  signal M_reg_4_13 : STD_LOGIC;
  signal M_reg_4_12 : STD_LOGIC;
  signal M_reg_4_11 : STD_LOGIC;
  signal M_reg_4_10 : STD_LOGIC;
  signal M_reg_4_9 : STD_LOGIC;
  signal M_reg_4_8 : STD_LOGIC;
  signal M_reg_4_7 : STD_LOGIC;
  signal M_reg_4_6 : STD_LOGIC;
  signal M_reg_4_5 : STD_LOGIC;
  signal M_reg_4_4 : STD_LOGIC;
  signal M_reg_4_3 : STD_LOGIC;
  signal M_reg_4_2 : STD_LOGIC;
  signal M_reg_4_1 : STD_LOGIC;
  signal M_reg_4_0 : STD_LOGIC;
  signal M_reg_5_31 : STD_LOGIC;
  signal M_reg_5_30 : STD_LOGIC;
  signal M_reg_5_29 : STD_LOGIC;
  signal M_reg_5_28 : STD_LOGIC;
  signal M_reg_5_27 : STD_LOGIC;
  signal M_reg_5_26 : STD_LOGIC;
  signal M_reg_5_25 : STD_LOGIC;
  signal M_reg_5_24 : STD_LOGIC;
  signal M_reg_5_23 : STD_LOGIC;
  signal M_reg_5_22 : STD_LOGIC;
  signal M_reg_5_21 : STD_LOGIC;
  signal M_reg_5_20 : STD_LOGIC;
  signal M_reg_5_19 : STD_LOGIC;
  signal M_reg_5_18 : STD_LOGIC;
  signal M_reg_5_17 : STD_LOGIC;
  signal M_reg_5_16 : STD_LOGIC;
  signal M_reg_5_15 : STD_LOGIC;
  signal M_reg_5_14 : STD_LOGIC;
  signal M_reg_5_13 : STD_LOGIC;
  signal M_reg_5_12 : STD_LOGIC;
  signal M_reg_5_11 : STD_LOGIC;
  signal M_reg_5_10 : STD_LOGIC;
  signal M_reg_5_9 : STD_LOGIC;
  signal M_reg_5_8 : STD_LOGIC;
  signal M_reg_5_7 : STD_LOGIC;
  signal M_reg_5_6 : STD_LOGIC;
  signal M_reg_5_5 : STD_LOGIC;
  signal M_reg_5_4 : STD_LOGIC;
  signal M_reg_5_3 : STD_LOGIC;
  signal M_reg_5_2 : STD_LOGIC;
  signal M_reg_5_1 : STD_LOGIC;
  signal M_reg_5_0 : STD_LOGIC;
  signal M_reg_6_31 : STD_LOGIC;
  signal M_reg_6_30 : STD_LOGIC;
  signal M_reg_6_29 : STD_LOGIC;
  signal M_reg_6_28 : STD_LOGIC;
  signal M_reg_6_27 : STD_LOGIC;
  signal M_reg_6_26 : STD_LOGIC;
  signal M_reg_6_25 : STD_LOGIC;
  signal M_reg_6_24 : STD_LOGIC;
  signal M_reg_6_23 : STD_LOGIC;
  signal M_reg_6_22 : STD_LOGIC;
  signal M_reg_6_21 : STD_LOGIC;
  signal M_reg_6_20 : STD_LOGIC;
  signal M_reg_6_19 : STD_LOGIC;
  signal M_reg_6_18 : STD_LOGIC;
  signal M_reg_6_17 : STD_LOGIC;
  signal M_reg_6_16 : STD_LOGIC;
  signal M_reg_6_15 : STD_LOGIC;
  signal M_reg_6_14 : STD_LOGIC;
  signal M_reg_6_13 : STD_LOGIC;
  signal M_reg_6_12 : STD_LOGIC;
  signal M_reg_6_11 : STD_LOGIC;
  signal M_reg_6_10 : STD_LOGIC;
  signal M_reg_6_9 : STD_LOGIC;
  signal M_reg_6_8 : STD_LOGIC;
  signal M_reg_6_7 : STD_LOGIC;
  signal M_reg_6_6 : STD_LOGIC;
  signal M_reg_6_5 : STD_LOGIC;
  signal M_reg_6_4 : STD_LOGIC;
  signal M_reg_6_3 : STD_LOGIC;
  signal M_reg_6_2 : STD_LOGIC;
  signal M_reg_6_1 : STD_LOGIC;
  signal M_reg_6_0 : STD_LOGIC;
  signal M_reg_7_31 : STD_LOGIC;
  signal M_reg_7_30 : STD_LOGIC;
  signal M_reg_7_29 : STD_LOGIC;
  signal M_reg_7_28 : STD_LOGIC;
  signal M_reg_7_27 : STD_LOGIC;
  signal M_reg_7_26 : STD_LOGIC;
  signal M_reg_7_25 : STD_LOGIC;
  signal M_reg_7_24 : STD_LOGIC;
  signal M_reg_7_23 : STD_LOGIC;
  signal M_reg_7_22 : STD_LOGIC;
  signal M_reg_7_21 : STD_LOGIC;
  signal M_reg_7_20 : STD_LOGIC;
  signal M_reg_7_19 : STD_LOGIC;
  signal M_reg_7_18 : STD_LOGIC;
  signal M_reg_7_17 : STD_LOGIC;
  signal M_reg_7_16 : STD_LOGIC;
  signal M_reg_7_15 : STD_LOGIC;
  signal M_reg_7_14 : STD_LOGIC;
  signal M_reg_7_13 : STD_LOGIC;
  signal M_reg_7_12 : STD_LOGIC;
  signal M_reg_7_11 : STD_LOGIC;
  signal M_reg_7_10 : STD_LOGIC;
  signal M_reg_7_9 : STD_LOGIC;
  signal M_reg_7_8 : STD_LOGIC;
  signal M_reg_7_7 : STD_LOGIC;
  signal M_reg_7_6 : STD_LOGIC;
  signal M_reg_7_5 : STD_LOGIC;
  signal M_reg_7_4 : STD_LOGIC;
  signal M_reg_7_3 : STD_LOGIC;
  signal M_reg_7_2 : STD_LOGIC;
  signal M_reg_7_1 : STD_LOGIC;
  signal M_reg_7_0 : STD_LOGIC;
  signal M_reg_8_31 : STD_LOGIC;
  signal M_reg_8_30 : STD_LOGIC;
  signal M_reg_8_29 : STD_LOGIC;
  signal M_reg_8_28 : STD_LOGIC;
  signal M_reg_8_27 : STD_LOGIC;
  signal M_reg_8_26 : STD_LOGIC;
  signal M_reg_8_25 : STD_LOGIC;
  signal M_reg_8_24 : STD_LOGIC;
  signal M_reg_8_23 : STD_LOGIC;
  signal M_reg_8_22 : STD_LOGIC;
  signal M_reg_8_21 : STD_LOGIC;
  signal M_reg_8_20 : STD_LOGIC;
  signal M_reg_8_19 : STD_LOGIC;
  signal M_reg_8_18 : STD_LOGIC;
  signal M_reg_8_17 : STD_LOGIC;
  signal M_reg_8_16 : STD_LOGIC;
  signal M_reg_8_15 : STD_LOGIC;
  signal M_reg_8_14 : STD_LOGIC;
  signal M_reg_8_13 : STD_LOGIC;
  signal M_reg_8_12 : STD_LOGIC;
  signal M_reg_8_11 : STD_LOGIC;
  signal M_reg_8_10 : STD_LOGIC;
  signal M_reg_8_9 : STD_LOGIC;
  signal M_reg_8_8 : STD_LOGIC;
  signal M_reg_8_7 : STD_LOGIC;
  signal M_reg_8_6 : STD_LOGIC;
  signal M_reg_8_5 : STD_LOGIC;
  signal M_reg_8_4 : STD_LOGIC;
  signal M_reg_8_3 : STD_LOGIC;
  signal M_reg_8_2 : STD_LOGIC;
  signal M_reg_8_1 : STD_LOGIC;
  signal M_reg_8_0 : STD_LOGIC;
  signal M_reg_9_31 : STD_LOGIC;
  signal M_reg_9_30 : STD_LOGIC;
  signal M_reg_9_29 : STD_LOGIC;
  signal M_reg_9_28 : STD_LOGIC;
  signal M_reg_9_27 : STD_LOGIC;
  signal M_reg_9_26 : STD_LOGIC;
  signal M_reg_9_25 : STD_LOGIC;
  signal M_reg_9_24 : STD_LOGIC;
  signal M_reg_9_23 : STD_LOGIC;
  signal M_reg_9_22 : STD_LOGIC;
  signal M_reg_9_21 : STD_LOGIC;
  signal M_reg_9_20 : STD_LOGIC;
  signal M_reg_9_19 : STD_LOGIC;
  signal M_reg_9_18 : STD_LOGIC;
  signal M_reg_9_17 : STD_LOGIC;
  signal M_reg_9_16 : STD_LOGIC;
  signal M_reg_9_15 : STD_LOGIC;
  signal M_reg_9_14 : STD_LOGIC;
  signal M_reg_9_13 : STD_LOGIC;
  signal M_reg_9_12 : STD_LOGIC;
  signal M_reg_9_11 : STD_LOGIC;
  signal M_reg_9_10 : STD_LOGIC;
  signal M_reg_9_9 : STD_LOGIC;
  signal M_reg_9_8 : STD_LOGIC;
  signal M_reg_9_7 : STD_LOGIC;
  signal M_reg_9_6 : STD_LOGIC;
  signal M_reg_9_5 : STD_LOGIC;
  signal M_reg_9_4 : STD_LOGIC;
  signal M_reg_9_3 : STD_LOGIC;
  signal M_reg_9_2 : STD_LOGIC;
  signal M_reg_9_1 : STD_LOGIC;
  signal M_reg_9_0 : STD_LOGIC;
  signal NLW_a_reg_31_i_3_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_e_reg_31_i_2_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_HASH_02_COUNTER_reg_30_i_3_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_HASH_02_COUNTER_reg_30_i_3_CO_UNCONNECTED_2 : STD_LOGIC;
  signal NLW_HASH_02_COUNTER_reg_30_i_3_CO_UNCONNECTED_1 : STD_LOGIC;
  signal NLW_HASH_02_COUNTER_reg_30_i_3_O_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_HASH_02_COUNTER_reg_30_i_3_O_UNCONNECTED_2 : STD_LOGIC;
  signal NLW_HV_reg_0_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_HV_reg_1_30_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_HV_reg_2_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_HV_reg_3_30_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_HV_reg_4_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_HV_reg_5_30_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_HV_reg_6_31_i_3_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_HV_reg_7_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_T1_reg_31_i_10_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_T1_reg_31_i_2_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_T2_reg_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_16_31_i_2_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_17_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_18_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_19_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_20_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_21_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_22_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_23_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_24_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_25_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_26_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_27_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_28_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_29_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_30_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_31_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_32_31_i_2_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_33_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_34_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_35_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_36_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_37_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_38_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_39_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_40_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_41_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_42_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_43_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_44_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_45_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_46_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_47_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_48_31_i_2_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_49_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_50_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_51_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_52_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_53_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_54_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_55_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_56_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_57_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_58_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_59_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_60_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_61_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_62_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal NLW_W_reg_63_31_i_1_CO_UNCONNECTED_3 : STD_LOGIC;
  signal ROTR11_out_1 : STD_LOGIC;
  signal ROTR11_out_2 : STD_LOGIC;
  signal ROTR11_out_3 : STD_LOGIC;
  signal ROTR11_out_4 : STD_LOGIC;
  signal ROTR11_out_5 : STD_LOGIC;
  signal ROTR11_out_6 : STD_LOGIC;
  signal ROTR11_out_7 : STD_LOGIC;
  signal ROTR11_out_8 : STD_LOGIC;
  signal ROTR11_out_9 : STD_LOGIC;
  signal ROTR11_out_10 : STD_LOGIC;
  signal ROTR11_out_11 : STD_LOGIC;
  signal ROTR11_out_12 : STD_LOGIC;
  signal ROTR11_out_13 : STD_LOGIC;
  signal ROTR11_out_14 : STD_LOGIC;
  signal ROTR11_out_15 : STD_LOGIC;
  signal ROTR11_out_16 : STD_LOGIC;
  signal ROTR11_out_17 : STD_LOGIC;
  signal ROTR11_out_18 : STD_LOGIC;
  signal ROTR11_out_19 : STD_LOGIC;
  signal ROTR11_out_20 : STD_LOGIC;
  signal ROTR11_out_21 : STD_LOGIC;
  signal ROTR11_out_22 : STD_LOGIC;
  signal ROTR11_out_23 : STD_LOGIC;
  signal ROTR11_out_24 : STD_LOGIC;
  signal ROTR11_out_25 : STD_LOGIC;
  signal ROTR11_out_26 : STD_LOGIC;
  signal ROTR11_out_27 : STD_LOGIC;
  signal ROTR11_out_28 : STD_LOGIC;
  signal ROTR11_out_29 : STD_LOGIC;
  signal ROTR11_out_30 : STD_LOGIC;
  signal ROTR11_out_31 : STD_LOGIC;
  signal ROTR11_out_32 : STD_LOGIC;
  signal ROTR2_out_1 : STD_LOGIC;
  signal ROTR2_out_2 : STD_LOGIC;
  signal ROTR2_out_3 : STD_LOGIC;
  signal ROTR2_out_4 : STD_LOGIC;
  signal ROTR2_out_5 : STD_LOGIC;
  signal ROTR2_out_6 : STD_LOGIC;
  signal ROTR2_out_7 : STD_LOGIC;
  signal ROTR2_out_8 : STD_LOGIC;
  signal ROTR2_out_9 : STD_LOGIC;
  signal ROTR2_out_10 : STD_LOGIC;
  signal ROTR2_out_11 : STD_LOGIC;
  signal ROTR2_out_12 : STD_LOGIC;
  signal ROTR2_out_13 : STD_LOGIC;
  signal ROTR2_out_14 : STD_LOGIC;
  signal ROTR2_out_15 : STD_LOGIC;
  signal ROTR2_out_16 : STD_LOGIC;
  signal ROTR2_out_17 : STD_LOGIC;
  signal ROTR2_out_18 : STD_LOGIC;
  signal ROTR2_out_19 : STD_LOGIC;
  signal ROTR2_out_20 : STD_LOGIC;
  signal ROTR2_out_21 : STD_LOGIC;
  signal ROTR2_out_22 : STD_LOGIC;
  signal ROTR2_out_23 : STD_LOGIC;
  signal ROTR2_out_24 : STD_LOGIC;
  signal ROTR2_out_25 : STD_LOGIC;
  signal ROTR2_out_26 : STD_LOGIC;
  signal ROTR2_out_27 : STD_LOGIC;
  signal ROTR2_out_28 : STD_LOGIC;
  signal ROTR2_out_29 : STD_LOGIC;
  signal ROTR2_out_30 : STD_LOGIC;
  signal ROTR2_out_31 : STD_LOGIC;
  signal ROTR2_out_32 : STD_LOGIC;
  signal rst_IBUF : STD_LOGIC;
  signal SIGMA_LCASE_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_0_1 : STD_LOGIC;
  signal SIGMA_LCASE_0_0 : STD_LOGIC;
  signal SIGMA_LCASE_0103_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_0103_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_0103_out_0 : STD_LOGIC;
  signal SIGMA_LCASE_0111_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_0111_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_0111_out_0 : STD_LOGIC;
  signal SIGMA_LCASE_0119_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_0119_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_0119_out_0 : STD_LOGIC;
  signal SIGMA_LCASE_0127_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_0127_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_0127_out_0 : STD_LOGIC;
  signal SIGMA_LCASE_0135_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_0135_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_0135_out_0 : STD_LOGIC;
  signal SIGMA_LCASE_0143_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_0143_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_0143_out_0 : STD_LOGIC;
  signal SIGMA_LCASE_0151_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_0151_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_0151_out_0 : STD_LOGIC;
  signal SIGMA_LCASE_0159_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_0159_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_0159_out_0 : STD_LOGIC;
  signal SIGMA_LCASE_015_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_015_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_015_out_0 : STD_LOGIC;
  signal SIGMA_LCASE_0167_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_0167_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_0167_out_0 : STD_LOGIC;
  signal SIGMA_LCASE_0175_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_0175_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_0175_out_0 : STD_LOGIC;
  signal SIGMA_LCASE_0183_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_0183_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_0183_out_0 : STD_LOGIC;
  signal SIGMA_LCASE_0191_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_0191_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_0191_out_0 : STD_LOGIC;
  signal SIGMA_LCASE_0199_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_0199_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_0199_out_0 : STD_LOGIC;
  signal SIGMA_LCASE_0207_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_0207_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_0207_out_0 : STD_LOGIC;
  signal SIGMA_LCASE_0215_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_0215_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_0215_out_0 : STD_LOGIC;
  signal SIGMA_LCASE_0223_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_0223_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_0223_out_0 : STD_LOGIC;
  signal SIGMA_LCASE_0231_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_0231_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_0231_out_0 : STD_LOGIC;
  signal SIGMA_LCASE_0239_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_0239_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_0239_out_0 : STD_LOGIC;
  signal SIGMA_LCASE_023_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_023_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_023_out_0 : STD_LOGIC;
  signal SIGMA_LCASE_0247_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_0247_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_0247_out_0 : STD_LOGIC;
  signal SIGMA_LCASE_0255_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_0255_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_0255_out_0 : STD_LOGIC;
  signal SIGMA_LCASE_0263_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_0263_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_0263_out_0 : STD_LOGIC;
  signal SIGMA_LCASE_0271_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_0271_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_0279_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_0279_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_0287_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_0287_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_0295_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_0295_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_0303_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_0303_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_0311_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_0311_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_0319_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_0319_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_031_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_031_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_031_out_0 : STD_LOGIC;
  signal SIGMA_LCASE_0327_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_0327_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_0335_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_0335_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_0343_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_0343_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_0351_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_0351_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_0359_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_0359_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_0367_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_0367_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_0375_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_0375_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_0383_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_0383_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_039_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_039_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_039_out_0 : STD_LOGIC;
  signal SIGMA_LCASE_047_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_047_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_047_out_0 : STD_LOGIC;
  signal SIGMA_LCASE_055_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_055_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_055_out_0 : STD_LOGIC;
  signal SIGMA_LCASE_063_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_063_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_063_out_0 : STD_LOGIC;
  signal SIGMA_LCASE_071_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_071_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_071_out_0 : STD_LOGIC;
  signal SIGMA_LCASE_079_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_079_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_079_out_0 : STD_LOGIC;
  signal SIGMA_LCASE_087_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_087_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_087_out_0 : STD_LOGIC;
  signal SIGMA_LCASE_095_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_095_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_095_out_0 : STD_LOGIC;
  signal SIGMA_LCASE_1_1 : STD_LOGIC;
  signal SIGMA_LCASE_1107_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_1107_out_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_1107_out_0_2 : STD_LOGIC;
  signal SIGMA_LCASE_1115_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_1115_out_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_1115_out_0_2 : STD_LOGIC;
  signal SIGMA_LCASE_1123_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_1123_out_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_1123_out_0_2 : STD_LOGIC;
  signal SIGMA_LCASE_1131_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_1131_out_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_1131_out_0_2 : STD_LOGIC;
  signal SIGMA_LCASE_1139_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_1139_out_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_1139_out_0_2 : STD_LOGIC;
  signal SIGMA_LCASE_1147_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_1147_out_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_1147_out_0_2 : STD_LOGIC;
  signal SIGMA_LCASE_1155_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_1155_out_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_1155_out_0_2 : STD_LOGIC;
  signal SIGMA_LCASE_1163_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_1163_out_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_1163_out_0_2 : STD_LOGIC;
  signal SIGMA_LCASE_1171_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_1171_out_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_1171_out_0_2 : STD_LOGIC;
  signal SIGMA_LCASE_1179_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_1179_out_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_1179_out_0_2 : STD_LOGIC;
  signal SIGMA_LCASE_1187_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_1187_out_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_1187_out_0_2 : STD_LOGIC;
  signal SIGMA_LCASE_1195_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_1195_out_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_1195_out_0_2 : STD_LOGIC;
  signal SIGMA_LCASE_119_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_119_out_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_119_out_0_2 : STD_LOGIC;
  signal SIGMA_LCASE_1203_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_1203_out_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_1203_out_0_2 : STD_LOGIC;
  signal SIGMA_LCASE_1211_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_1211_out_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_1211_out_0_2 : STD_LOGIC;
  signal SIGMA_LCASE_1219_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_1219_out_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_1219_out_0_2 : STD_LOGIC;
  signal SIGMA_LCASE_1227_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_1227_out_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_1227_out_0_2 : STD_LOGIC;
  signal SIGMA_LCASE_1235_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_1235_out_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_1235_out_0_2 : STD_LOGIC;
  signal SIGMA_LCASE_1243_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_1243_out_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_1243_out_0_2 : STD_LOGIC;
  signal SIGMA_LCASE_1251_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_1251_out_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_1251_out_0_2 : STD_LOGIC;
  signal SIGMA_LCASE_1259_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_1259_out_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_1259_out_0_2 : STD_LOGIC;
  signal SIGMA_LCASE_1267_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_1267_out_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_1267_out_0_2 : STD_LOGIC;
  signal SIGMA_LCASE_1275_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_1275_out_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_1275_out_0_2 : STD_LOGIC;
  signal SIGMA_LCASE_127_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_127_out_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_127_out_0_2 : STD_LOGIC;
  signal SIGMA_LCASE_1283_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_1283_out_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_1283_out_0_2 : STD_LOGIC;
  signal SIGMA_LCASE_1291_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_1291_out_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_1291_out_0_2 : STD_LOGIC;
  signal SIGMA_LCASE_1299_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_1299_out_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_1299_out_0_2 : STD_LOGIC;
  signal SIGMA_LCASE_1307_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_1307_out_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_1307_out_0_2 : STD_LOGIC;
  signal SIGMA_LCASE_1315_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_1315_out_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_1315_out_0_2 : STD_LOGIC;
  signal SIGMA_LCASE_1323_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_1323_out_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_1323_out_0_2 : STD_LOGIC;
  signal SIGMA_LCASE_1331_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_1331_out_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_1331_out_0_2 : STD_LOGIC;
  signal SIGMA_LCASE_1339_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_1347_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_1355_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_135_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_135_out_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_135_out_0_2 : STD_LOGIC;
  signal SIGMA_LCASE_1363_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_1371_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_1379_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_1387_out_30 : STD_LOGIC;
  signal SIGMA_LCASE_143_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_143_out_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_143_out_0_2 : STD_LOGIC;
  signal SIGMA_LCASE_151_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_151_out_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_151_out_0_2 : STD_LOGIC;
  signal SIGMA_LCASE_159_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_159_out_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_159_out_0_2 : STD_LOGIC;
  signal SIGMA_LCASE_167_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_167_out_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_167_out_0_2 : STD_LOGIC;
  signal SIGMA_LCASE_175_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_175_out_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_175_out_0_2 : STD_LOGIC;
  signal SIGMA_LCASE_183_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_183_out_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_183_out_0_2 : STD_LOGIC;
  signal SIGMA_LCASE_191_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_191_out_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_191_out_0_2 : STD_LOGIC;
  signal SIGMA_LCASE_199_out_1 : STD_LOGIC;
  signal SIGMA_LCASE_199_out_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_199_out_0_2 : STD_LOGIC;
  signal SIGMA_LCASE_1_0_30 : STD_LOGIC;
  signal SIGMA_LCASE_1_0_2 : STD_LOGIC;
  signal SIGMA_UCASE_0_30 : STD_LOGIC;
  signal SIGMA_UCASE_0_29 : STD_LOGIC;
  signal SIGMA_UCASE_0_28 : STD_LOGIC;
  signal SIGMA_UCASE_0_27 : STD_LOGIC;
  signal SIGMA_UCASE_0_26 : STD_LOGIC;
  signal SIGMA_UCASE_0_25 : STD_LOGIC;
  signal SIGMA_UCASE_0_24 : STD_LOGIC;
  signal SIGMA_UCASE_0_23 : STD_LOGIC;
  signal SIGMA_UCASE_0_22 : STD_LOGIC;
  signal SIGMA_UCASE_0_21 : STD_LOGIC;
  signal SIGMA_UCASE_0_20 : STD_LOGIC;
  signal SIGMA_UCASE_0_19 : STD_LOGIC;
  signal SIGMA_UCASE_0_18 : STD_LOGIC;
  signal SIGMA_UCASE_0_17 : STD_LOGIC;
  signal SIGMA_UCASE_0_16 : STD_LOGIC;
  signal SIGMA_UCASE_0_15 : STD_LOGIC;
  signal SIGMA_UCASE_0_14 : STD_LOGIC;
  signal SIGMA_UCASE_0_13 : STD_LOGIC;
  signal SIGMA_UCASE_0_12 : STD_LOGIC;
  signal SIGMA_UCASE_0_11 : STD_LOGIC;
  signal SIGMA_UCASE_0_10 : STD_LOGIC;
  signal SIGMA_UCASE_0_9 : STD_LOGIC;
  signal SIGMA_UCASE_0_8 : STD_LOGIC;
  signal SIGMA_UCASE_0_7 : STD_LOGIC;
  signal SIGMA_UCASE_0_6 : STD_LOGIC;
  signal SIGMA_UCASE_0_5 : STD_LOGIC;
  signal SIGMA_UCASE_0_4 : STD_LOGIC;
  signal SIGMA_UCASE_0_3 : STD_LOGIC;
  signal SIGMA_UCASE_0_2 : STD_LOGIC;
  signal SIGMA_UCASE_0_1 : STD_LOGIC;
  signal SIGMA_UCASE_0_0 : STD_LOGIC;
  signal T100_in_31 : STD_LOGIC;
  signal T100_in_30 : STD_LOGIC;
  signal T100_in_29 : STD_LOGIC;
  signal T100_in_28 : STD_LOGIC;
  signal T100_in_27 : STD_LOGIC;
  signal T100_in_26 : STD_LOGIC;
  signal T100_in_25 : STD_LOGIC;
  signal T100_in_24 : STD_LOGIC;
  signal T100_in_23 : STD_LOGIC;
  signal T100_in_22 : STD_LOGIC;
  signal T100_in_21 : STD_LOGIC;
  signal T100_in_20 : STD_LOGIC;
  signal T100_in_19 : STD_LOGIC;
  signal T100_in_18 : STD_LOGIC;
  signal T100_in_17 : STD_LOGIC;
  signal T100_in_16 : STD_LOGIC;
  signal T100_in_15 : STD_LOGIC;
  signal T100_in_14 : STD_LOGIC;
  signal T100_in_13 : STD_LOGIC;
  signal T100_in_12 : STD_LOGIC;
  signal T100_in_11 : STD_LOGIC;
  signal T100_in_10 : STD_LOGIC;
  signal T100_in_9 : STD_LOGIC;
  signal T100_in_8 : STD_LOGIC;
  signal T100_in_7 : STD_LOGIC;
  signal T100_in_6 : STD_LOGIC;
  signal T100_in_5 : STD_LOGIC;
  signal T100_in_4 : STD_LOGIC;
  signal T100_in_3 : STD_LOGIC;
  signal T100_in_2 : STD_LOGIC;
  signal T100_in_1 : STD_LOGIC;
  signal T100_in_0 : STD_LOGIC;
  signal T1_11_i_100_n_0 : STD_LOGIC;
  signal T1_11_i_101_n_0 : STD_LOGIC;
  signal T1_11_i_102_n_0 : STD_LOGIC;
  signal T1_11_i_103_n_0 : STD_LOGIC;
  signal T1_11_i_104_n_0 : STD_LOGIC;
  signal T1_11_i_105_n_0 : STD_LOGIC;
  signal T1_11_i_106_n_0 : STD_LOGIC;
  signal T1_11_i_10_n_0 : STD_LOGIC;
  signal T1_11_i_11_n_0 : STD_LOGIC;
  signal T1_11_i_12_n_0 : STD_LOGIC;
  signal T1_11_i_14_n_0 : STD_LOGIC;
  signal T1_11_i_15_n_0 : STD_LOGIC;
  signal T1_11_i_16_n_0 : STD_LOGIC;
  signal T1_11_i_17_n_0 : STD_LOGIC;
  signal T1_11_i_18_n_0 : STD_LOGIC;
  signal T1_11_i_19_n_0 : STD_LOGIC;
  signal T1_11_i_20_n_0 : STD_LOGIC;
  signal T1_11_i_21_n_0 : STD_LOGIC;
  signal T1_11_i_22_n_0 : STD_LOGIC;
  signal T1_11_i_23_n_0 : STD_LOGIC;
  signal T1_11_i_24_n_0 : STD_LOGIC;
  signal T1_11_i_25_n_0 : STD_LOGIC;
  signal T1_11_i_26_n_0 : STD_LOGIC;
  signal T1_11_i_27_n_0 : STD_LOGIC;
  signal T1_11_i_28_n_0 : STD_LOGIC;
  signal T1_11_i_29_n_0 : STD_LOGIC;
  signal T1_11_i_2_n_0 : STD_LOGIC;
  signal T1_11_i_30_n_0 : STD_LOGIC;
  signal T1_11_i_31_n_0 : STD_LOGIC;
  signal T1_11_i_32_n_0 : STD_LOGIC;
  signal T1_11_i_33_n_0 : STD_LOGIC;
  signal T1_11_i_34_n_0 : STD_LOGIC;
  signal T1_11_i_35_n_0 : STD_LOGIC;
  signal T1_11_i_36_n_0 : STD_LOGIC;
  signal T1_11_i_37_n_0 : STD_LOGIC;
  signal T1_11_i_38_n_0 : STD_LOGIC;
  signal T1_11_i_39_n_0 : STD_LOGIC;
  signal T1_11_i_3_n_0 : STD_LOGIC;
  signal T1_11_i_40_n_0 : STD_LOGIC;
  signal T1_11_i_41_n_0 : STD_LOGIC;
  signal T1_11_i_42_n_0 : STD_LOGIC;
  signal T1_11_i_43_n_0 : STD_LOGIC;
  signal T1_11_i_44_n_0 : STD_LOGIC;
  signal T1_11_i_45_n_0 : STD_LOGIC;
  signal T1_11_i_46_n_0 : STD_LOGIC;
  signal T1_11_i_47_n_0 : STD_LOGIC;
  signal T1_11_i_48_n_0 : STD_LOGIC;
  signal T1_11_i_49_n_0 : STD_LOGIC;
  signal T1_11_i_4_n_0 : STD_LOGIC;
  signal T1_11_i_50_n_0 : STD_LOGIC;
  signal T1_11_i_51_n_0 : STD_LOGIC;
  signal T1_11_i_52_n_0 : STD_LOGIC;
  signal T1_11_i_53_n_0 : STD_LOGIC;
  signal T1_11_i_54_n_0 : STD_LOGIC;
  signal T1_11_i_55_n_0 : STD_LOGIC;
  signal T1_11_i_56_n_0 : STD_LOGIC;
  signal T1_11_i_57_n_0 : STD_LOGIC;
  signal T1_11_i_58_n_0 : STD_LOGIC;
  signal T1_11_i_59_n_0 : STD_LOGIC;
  signal T1_11_i_5_n_0 : STD_LOGIC;
  signal T1_11_i_60_n_0 : STD_LOGIC;
  signal T1_11_i_61_n_0 : STD_LOGIC;
  signal T1_11_i_62_n_0 : STD_LOGIC;
  signal T1_11_i_63_n_0 : STD_LOGIC;
  signal T1_11_i_64_n_0 : STD_LOGIC;
  signal T1_11_i_65_n_0 : STD_LOGIC;
  signal T1_11_i_66_n_0 : STD_LOGIC;
  signal T1_11_i_67_n_0 : STD_LOGIC;
  signal T1_11_i_68_n_0 : STD_LOGIC;
  signal T1_11_i_69_n_0 : STD_LOGIC;
  signal T1_11_i_6_n_0 : STD_LOGIC;
  signal T1_11_i_70_n_0 : STD_LOGIC;
  signal T1_11_i_71_n_0 : STD_LOGIC;
  signal T1_11_i_72_n_0 : STD_LOGIC;
  signal T1_11_i_73_n_0 : STD_LOGIC;
  signal T1_11_i_74_n_0 : STD_LOGIC;
  signal T1_11_i_75_n_0 : STD_LOGIC;
  signal T1_11_i_76_n_0 : STD_LOGIC;
  signal T1_11_i_77_n_0 : STD_LOGIC;
  signal T1_11_i_78_n_0 : STD_LOGIC;
  signal T1_11_i_79_n_0 : STD_LOGIC;
  signal T1_11_i_7_n_0 : STD_LOGIC;
  signal T1_11_i_80_n_0 : STD_LOGIC;
  signal T1_11_i_81_n_0 : STD_LOGIC;
  signal T1_11_i_82_n_0 : STD_LOGIC;
  signal T1_11_i_83_n_0 : STD_LOGIC;
  signal T1_11_i_84_n_0 : STD_LOGIC;
  signal T1_11_i_85_n_0 : STD_LOGIC;
  signal T1_11_i_86_n_0 : STD_LOGIC;
  signal T1_11_i_87_n_0 : STD_LOGIC;
  signal T1_11_i_88_n_0 : STD_LOGIC;
  signal T1_11_i_89_n_0 : STD_LOGIC;
  signal T1_11_i_8_n_0 : STD_LOGIC;
  signal T1_11_i_90_n_0 : STD_LOGIC;
  signal T1_11_i_91_n_0 : STD_LOGIC;
  signal T1_11_i_92_n_0 : STD_LOGIC;
  signal T1_11_i_93_n_0 : STD_LOGIC;
  signal T1_11_i_94_n_0 : STD_LOGIC;
  signal T1_11_i_95_n_0 : STD_LOGIC;
  signal T1_11_i_96_n_0 : STD_LOGIC;
  signal T1_11_i_97_n_0 : STD_LOGIC;
  signal T1_11_i_98_n_0 : STD_LOGIC;
  signal T1_11_i_99_n_0 : STD_LOGIC;
  signal T1_11_i_9_n_0 : STD_LOGIC;
  signal T1_15_i_100_n_0 : STD_LOGIC;
  signal T1_15_i_101_n_0 : STD_LOGIC;
  signal T1_15_i_102_n_0 : STD_LOGIC;
  signal T1_15_i_103_n_0 : STD_LOGIC;
  signal T1_15_i_104_n_0 : STD_LOGIC;
  signal T1_15_i_105_n_0 : STD_LOGIC;
  signal T1_15_i_106_n_0 : STD_LOGIC;
  signal T1_15_i_107_n_0 : STD_LOGIC;
  signal T1_15_i_108_n_0 : STD_LOGIC;
  signal T1_15_i_109_n_0 : STD_LOGIC;
  signal T1_15_i_10_n_0 : STD_LOGIC;
  signal T1_15_i_110_n_0 : STD_LOGIC;
  signal T1_15_i_111_n_0 : STD_LOGIC;
  signal T1_15_i_112_n_0 : STD_LOGIC;
  signal T1_15_i_11_n_0 : STD_LOGIC;
  signal T1_15_i_12_n_0 : STD_LOGIC;
  signal T1_15_i_14_n_0 : STD_LOGIC;
  signal T1_15_i_15_n_0 : STD_LOGIC;
  signal T1_15_i_16_n_0 : STD_LOGIC;
  signal T1_15_i_17_n_0 : STD_LOGIC;
  signal T1_15_i_18_n_0 : STD_LOGIC;
  signal T1_15_i_19_n_0 : STD_LOGIC;
  signal T1_15_i_20_n_0 : STD_LOGIC;
  signal T1_15_i_21_n_0 : STD_LOGIC;
  signal T1_15_i_22_n_0 : STD_LOGIC;
  signal T1_15_i_23_n_0 : STD_LOGIC;
  signal T1_15_i_24_n_0 : STD_LOGIC;
  signal T1_15_i_25_n_0 : STD_LOGIC;
  signal T1_15_i_26_n_0 : STD_LOGIC;
  signal T1_15_i_27_n_0 : STD_LOGIC;
  signal T1_15_i_28_n_0 : STD_LOGIC;
  signal T1_15_i_2_n_0 : STD_LOGIC;
  signal T1_15_i_30_n_0 : STD_LOGIC;
  signal T1_15_i_31_n_0 : STD_LOGIC;
  signal T1_15_i_32_n_0 : STD_LOGIC;
  signal T1_15_i_34_n_0 : STD_LOGIC;
  signal T1_15_i_35_n_0 : STD_LOGIC;
  signal T1_15_i_36_n_0 : STD_LOGIC;
  signal T1_15_i_38_n_0 : STD_LOGIC;
  signal T1_15_i_39_n_0 : STD_LOGIC;
  signal T1_15_i_3_n_0 : STD_LOGIC;
  signal T1_15_i_40_n_0 : STD_LOGIC;
  signal T1_15_i_41_n_0 : STD_LOGIC;
  signal T1_15_i_42_n_0 : STD_LOGIC;
  signal T1_15_i_43_n_0 : STD_LOGIC;
  signal T1_15_i_44_n_0 : STD_LOGIC;
  signal T1_15_i_45_n_0 : STD_LOGIC;
  signal T1_15_i_46_n_0 : STD_LOGIC;
  signal T1_15_i_47_n_0 : STD_LOGIC;
  signal T1_15_i_48_n_0 : STD_LOGIC;
  signal T1_15_i_49_n_0 : STD_LOGIC;
  signal T1_15_i_4_n_0 : STD_LOGIC;
  signal T1_15_i_50_n_0 : STD_LOGIC;
  signal T1_15_i_53_n_0 : STD_LOGIC;
  signal T1_15_i_54_n_0 : STD_LOGIC;
  signal T1_15_i_55_n_0 : STD_LOGIC;
  signal T1_15_i_56_n_0 : STD_LOGIC;
  signal T1_15_i_57_n_0 : STD_LOGIC;
  signal T1_15_i_58_n_0 : STD_LOGIC;
  signal T1_15_i_59_n_0 : STD_LOGIC;
  signal T1_15_i_5_n_0 : STD_LOGIC;
  signal T1_15_i_60_n_0 : STD_LOGIC;
  signal T1_15_i_61_n_0 : STD_LOGIC;
  signal T1_15_i_62_n_0 : STD_LOGIC;
  signal T1_15_i_63_n_0 : STD_LOGIC;
  signal T1_15_i_64_n_0 : STD_LOGIC;
  signal T1_15_i_67_n_0 : STD_LOGIC;
  signal T1_15_i_68_n_0 : STD_LOGIC;
  signal T1_15_i_69_n_0 : STD_LOGIC;
  signal T1_15_i_6_n_0 : STD_LOGIC;
  signal T1_15_i_70_n_0 : STD_LOGIC;
  signal T1_15_i_71_n_0 : STD_LOGIC;
  signal T1_15_i_72_n_0 : STD_LOGIC;
  signal T1_15_i_73_n_0 : STD_LOGIC;
  signal T1_15_i_74_n_0 : STD_LOGIC;
  signal T1_15_i_75_n_0 : STD_LOGIC;
  signal T1_15_i_76_n_0 : STD_LOGIC;
  signal T1_15_i_77_n_0 : STD_LOGIC;
  signal T1_15_i_78_n_0 : STD_LOGIC;
  signal T1_15_i_7_n_0 : STD_LOGIC;
  signal T1_15_i_81_n_0 : STD_LOGIC;
  signal T1_15_i_82_n_0 : STD_LOGIC;
  signal T1_15_i_83_n_0 : STD_LOGIC;
  signal T1_15_i_84_n_0 : STD_LOGIC;
  signal T1_15_i_85_n_0 : STD_LOGIC;
  signal T1_15_i_86_n_0 : STD_LOGIC;
  signal T1_15_i_87_n_0 : STD_LOGIC;
  signal T1_15_i_88_n_0 : STD_LOGIC;
  signal T1_15_i_89_n_0 : STD_LOGIC;
  signal T1_15_i_8_n_0 : STD_LOGIC;
  signal T1_15_i_90_n_0 : STD_LOGIC;
  signal T1_15_i_91_n_0 : STD_LOGIC;
  signal T1_15_i_92_n_0 : STD_LOGIC;
  signal T1_15_i_93_n_0 : STD_LOGIC;
  signal T1_15_i_94_n_0 : STD_LOGIC;
  signal T1_15_i_95_n_0 : STD_LOGIC;
  signal T1_15_i_96_n_0 : STD_LOGIC;
  signal T1_15_i_97_n_0 : STD_LOGIC;
  signal T1_15_i_98_n_0 : STD_LOGIC;
  signal T1_15_i_99_n_0 : STD_LOGIC;
  signal T1_15_i_9_n_0 : STD_LOGIC;
  signal T1_19_i_101_n_0 : STD_LOGIC;
  signal T1_19_i_102_n_0 : STD_LOGIC;
  signal T1_19_i_103_n_0 : STD_LOGIC;
  signal T1_19_i_104_n_0 : STD_LOGIC;
  signal T1_19_i_105_n_0 : STD_LOGIC;
  signal T1_19_i_106_n_0 : STD_LOGIC;
  signal T1_19_i_107_n_0 : STD_LOGIC;
  signal T1_19_i_108_n_0 : STD_LOGIC;
  signal T1_19_i_10_n_0 : STD_LOGIC;
  signal T1_19_i_11_n_0 : STD_LOGIC;
  signal T1_19_i_12_n_0 : STD_LOGIC;
  signal T1_19_i_14_n_0 : STD_LOGIC;
  signal T1_19_i_15_n_0 : STD_LOGIC;
  signal T1_19_i_16_n_0 : STD_LOGIC;
  signal T1_19_i_17_n_0 : STD_LOGIC;
  signal T1_19_i_18_n_0 : STD_LOGIC;
  signal T1_19_i_19_n_0 : STD_LOGIC;
  signal T1_19_i_20_n_0 : STD_LOGIC;
  signal T1_19_i_21_n_0 : STD_LOGIC;
  signal T1_19_i_22_n_0 : STD_LOGIC;
  signal T1_19_i_23_n_0 : STD_LOGIC;
  signal T1_19_i_24_n_0 : STD_LOGIC;
  signal T1_19_i_25_n_0 : STD_LOGIC;
  signal T1_19_i_26_n_0 : STD_LOGIC;
  signal T1_19_i_27_n_0 : STD_LOGIC;
  signal T1_19_i_28_n_0 : STD_LOGIC;
  signal T1_19_i_29_n_0 : STD_LOGIC;
  signal T1_19_i_2_n_0 : STD_LOGIC;
  signal T1_19_i_30_n_0 : STD_LOGIC;
  signal T1_19_i_31_n_0 : STD_LOGIC;
  signal T1_19_i_32_n_0 : STD_LOGIC;
  signal T1_19_i_33_n_0 : STD_LOGIC;
  signal T1_19_i_34_n_0 : STD_LOGIC;
  signal T1_19_i_35_n_0 : STD_LOGIC;
  signal T1_19_i_36_n_0 : STD_LOGIC;
  signal T1_19_i_37_n_0 : STD_LOGIC;
  signal T1_19_i_38_n_0 : STD_LOGIC;
  signal T1_19_i_39_n_0 : STD_LOGIC;
  signal T1_19_i_3_n_0 : STD_LOGIC;
  signal T1_19_i_40_n_0 : STD_LOGIC;
  signal T1_19_i_42_n_0 : STD_LOGIC;
  signal T1_19_i_43_n_0 : STD_LOGIC;
  signal T1_19_i_44_n_0 : STD_LOGIC;
  signal T1_19_i_45_n_0 : STD_LOGIC;
  signal T1_19_i_46_n_0 : STD_LOGIC;
  signal T1_19_i_47_n_0 : STD_LOGIC;
  signal T1_19_i_48_n_0 : STD_LOGIC;
  signal T1_19_i_49_n_0 : STD_LOGIC;
  signal T1_19_i_4_n_0 : STD_LOGIC;
  signal T1_19_i_50_n_0 : STD_LOGIC;
  signal T1_19_i_51_n_0 : STD_LOGIC;
  signal T1_19_i_52_n_0 : STD_LOGIC;
  signal T1_19_i_53_n_0 : STD_LOGIC;
  signal T1_19_i_54_n_0 : STD_LOGIC;
  signal T1_19_i_55_n_0 : STD_LOGIC;
  signal T1_19_i_56_n_0 : STD_LOGIC;
  signal T1_19_i_57_n_0 : STD_LOGIC;
  signal T1_19_i_58_n_0 : STD_LOGIC;
  signal T1_19_i_59_n_0 : STD_LOGIC;
  signal T1_19_i_5_n_0 : STD_LOGIC;
  signal T1_19_i_60_n_0 : STD_LOGIC;
  signal T1_19_i_61_n_0 : STD_LOGIC;
  signal T1_19_i_62_n_0 : STD_LOGIC;
  signal T1_19_i_63_n_0 : STD_LOGIC;
  signal T1_19_i_64_n_0 : STD_LOGIC;
  signal T1_19_i_65_n_0 : STD_LOGIC;
  signal T1_19_i_66_n_0 : STD_LOGIC;
  signal T1_19_i_67_n_0 : STD_LOGIC;
  signal T1_19_i_68_n_0 : STD_LOGIC;
  signal T1_19_i_69_n_0 : STD_LOGIC;
  signal T1_19_i_6_n_0 : STD_LOGIC;
  signal T1_19_i_70_n_0 : STD_LOGIC;
  signal T1_19_i_71_n_0 : STD_LOGIC;
  signal T1_19_i_72_n_0 : STD_LOGIC;
  signal T1_19_i_73_n_0 : STD_LOGIC;
  signal T1_19_i_74_n_0 : STD_LOGIC;
  signal T1_19_i_75_n_0 : STD_LOGIC;
  signal T1_19_i_76_n_0 : STD_LOGIC;
  signal T1_19_i_77_n_0 : STD_LOGIC;
  signal T1_19_i_78_n_0 : STD_LOGIC;
  signal T1_19_i_79_n_0 : STD_LOGIC;
  signal T1_19_i_7_n_0 : STD_LOGIC;
  signal T1_19_i_80_n_0 : STD_LOGIC;
  signal T1_19_i_81_n_0 : STD_LOGIC;
  signal T1_19_i_82_n_0 : STD_LOGIC;
  signal T1_19_i_83_n_0 : STD_LOGIC;
  signal T1_19_i_84_n_0 : STD_LOGIC;
  signal T1_19_i_85_n_0 : STD_LOGIC;
  signal T1_19_i_86_n_0 : STD_LOGIC;
  signal T1_19_i_87_n_0 : STD_LOGIC;
  signal T1_19_i_88_n_0 : STD_LOGIC;
  signal T1_19_i_89_n_0 : STD_LOGIC;
  signal T1_19_i_8_n_0 : STD_LOGIC;
  signal T1_19_i_90_n_0 : STD_LOGIC;
  signal T1_19_i_91_n_0 : STD_LOGIC;
  signal T1_19_i_92_n_0 : STD_LOGIC;
  signal T1_19_i_93_n_0 : STD_LOGIC;
  signal T1_19_i_94_n_0 : STD_LOGIC;
  signal T1_19_i_95_n_0 : STD_LOGIC;
  signal T1_19_i_96_n_0 : STD_LOGIC;
  signal T1_19_i_97_n_0 : STD_LOGIC;
  signal T1_19_i_98_n_0 : STD_LOGIC;
  signal T1_19_i_9_n_0 : STD_LOGIC;
  signal T1_23_i_100_n_0 : STD_LOGIC;
  signal T1_23_i_101_n_0 : STD_LOGIC;
  signal T1_23_i_102_n_0 : STD_LOGIC;
  signal T1_23_i_103_n_0 : STD_LOGIC;
  signal T1_23_i_104_n_0 : STD_LOGIC;
  signal T1_23_i_105_n_0 : STD_LOGIC;
  signal T1_23_i_106_n_0 : STD_LOGIC;
  signal T1_23_i_107_n_0 : STD_LOGIC;
  signal T1_23_i_108_n_0 : STD_LOGIC;
  signal T1_23_i_10_n_0 : STD_LOGIC;
  signal T1_23_i_11_n_0 : STD_LOGIC;
  signal T1_23_i_12_n_0 : STD_LOGIC;
  signal T1_23_i_14_n_0 : STD_LOGIC;
  signal T1_23_i_15_n_0 : STD_LOGIC;
  signal T1_23_i_16_n_0 : STD_LOGIC;
  signal T1_23_i_17_n_0 : STD_LOGIC;
  signal T1_23_i_18_n_0 : STD_LOGIC;
  signal T1_23_i_19_n_0 : STD_LOGIC;
  signal T1_23_i_20_n_0 : STD_LOGIC;
  signal T1_23_i_21_n_0 : STD_LOGIC;
  signal T1_23_i_22_n_0 : STD_LOGIC;
  signal T1_23_i_23_n_0 : STD_LOGIC;
  signal T1_23_i_24_n_0 : STD_LOGIC;
  signal T1_23_i_25_n_0 : STD_LOGIC;
  signal T1_23_i_26_n_0 : STD_LOGIC;
  signal T1_23_i_27_n_0 : STD_LOGIC;
  signal T1_23_i_28_n_0 : STD_LOGIC;
  signal T1_23_i_29_n_0 : STD_LOGIC;
  signal T1_23_i_2_n_0 : STD_LOGIC;
  signal T1_23_i_30_n_0 : STD_LOGIC;
  signal T1_23_i_31_n_0 : STD_LOGIC;
  signal T1_23_i_32_n_0 : STD_LOGIC;
  signal T1_23_i_33_n_0 : STD_LOGIC;
  signal T1_23_i_34_n_0 : STD_LOGIC;
  signal T1_23_i_35_n_0 : STD_LOGIC;
  signal T1_23_i_36_n_0 : STD_LOGIC;
  signal T1_23_i_37_n_0 : STD_LOGIC;
  signal T1_23_i_38_n_0 : STD_LOGIC;
  signal T1_23_i_39_n_0 : STD_LOGIC;
  signal T1_23_i_3_n_0 : STD_LOGIC;
  signal T1_23_i_41_n_0 : STD_LOGIC;
  signal T1_23_i_42_n_0 : STD_LOGIC;
  signal T1_23_i_43_n_0 : STD_LOGIC;
  signal T1_23_i_44_n_0 : STD_LOGIC;
  signal T1_23_i_45_n_0 : STD_LOGIC;
  signal T1_23_i_46_n_0 : STD_LOGIC;
  signal T1_23_i_47_n_0 : STD_LOGIC;
  signal T1_23_i_48_n_0 : STD_LOGIC;
  signal T1_23_i_49_n_0 : STD_LOGIC;
  signal T1_23_i_4_n_0 : STD_LOGIC;
  signal T1_23_i_50_n_0 : STD_LOGIC;
  signal T1_23_i_51_n_0 : STD_LOGIC;
  signal T1_23_i_52_n_0 : STD_LOGIC;
  signal T1_23_i_53_n_0 : STD_LOGIC;
  signal T1_23_i_54_n_0 : STD_LOGIC;
  signal T1_23_i_55_n_0 : STD_LOGIC;
  signal T1_23_i_56_n_0 : STD_LOGIC;
  signal T1_23_i_57_n_0 : STD_LOGIC;
  signal T1_23_i_58_n_0 : STD_LOGIC;
  signal T1_23_i_59_n_0 : STD_LOGIC;
  signal T1_23_i_5_n_0 : STD_LOGIC;
  signal T1_23_i_60_n_0 : STD_LOGIC;
  signal T1_23_i_61_n_0 : STD_LOGIC;
  signal T1_23_i_62_n_0 : STD_LOGIC;
  signal T1_23_i_63_n_0 : STD_LOGIC;
  signal T1_23_i_64_n_0 : STD_LOGIC;
  signal T1_23_i_65_n_0 : STD_LOGIC;
  signal T1_23_i_66_n_0 : STD_LOGIC;
  signal T1_23_i_67_n_0 : STD_LOGIC;
  signal T1_23_i_68_n_0 : STD_LOGIC;
  signal T1_23_i_69_n_0 : STD_LOGIC;
  signal T1_23_i_6_n_0 : STD_LOGIC;
  signal T1_23_i_70_n_0 : STD_LOGIC;
  signal T1_23_i_71_n_0 : STD_LOGIC;
  signal T1_23_i_72_n_0 : STD_LOGIC;
  signal T1_23_i_73_n_0 : STD_LOGIC;
  signal T1_23_i_74_n_0 : STD_LOGIC;
  signal T1_23_i_75_n_0 : STD_LOGIC;
  signal T1_23_i_76_n_0 : STD_LOGIC;
  signal T1_23_i_77_n_0 : STD_LOGIC;
  signal T1_23_i_78_n_0 : STD_LOGIC;
  signal T1_23_i_79_n_0 : STD_LOGIC;
  signal T1_23_i_7_n_0 : STD_LOGIC;
  signal T1_23_i_80_n_0 : STD_LOGIC;
  signal T1_23_i_81_n_0 : STD_LOGIC;
  signal T1_23_i_82_n_0 : STD_LOGIC;
  signal T1_23_i_83_n_0 : STD_LOGIC;
  signal T1_23_i_84_n_0 : STD_LOGIC;
  signal T1_23_i_85_n_0 : STD_LOGIC;
  signal T1_23_i_86_n_0 : STD_LOGIC;
  signal T1_23_i_87_n_0 : STD_LOGIC;
  signal T1_23_i_88_n_0 : STD_LOGIC;
  signal T1_23_i_89_n_0 : STD_LOGIC;
  signal T1_23_i_8_n_0 : STD_LOGIC;
  signal T1_23_i_90_n_0 : STD_LOGIC;
  signal T1_23_i_91_n_0 : STD_LOGIC;
  signal T1_23_i_92_n_0 : STD_LOGIC;
  signal T1_23_i_93_n_0 : STD_LOGIC;
  signal T1_23_i_94_n_0 : STD_LOGIC;
  signal T1_23_i_97_n_0 : STD_LOGIC;
  signal T1_23_i_98_n_0 : STD_LOGIC;
  signal T1_23_i_99_n_0 : STD_LOGIC;
  signal T1_23_i_9_n_0 : STD_LOGIC;
  signal T1_27_i_100_n_0 : STD_LOGIC;
  signal T1_27_i_101_n_0 : STD_LOGIC;
  signal T1_27_i_102_n_0 : STD_LOGIC;
  signal T1_27_i_103_n_0 : STD_LOGIC;
  signal T1_27_i_104_n_0 : STD_LOGIC;
  signal T1_27_i_105_n_0 : STD_LOGIC;
  signal T1_27_i_106_n_0 : STD_LOGIC;
  signal T1_27_i_107_n_0 : STD_LOGIC;
  signal T1_27_i_108_n_0 : STD_LOGIC;
  signal T1_27_i_10_n_0 : STD_LOGIC;
  signal T1_27_i_11_n_0 : STD_LOGIC;
  signal T1_27_i_12_n_0 : STD_LOGIC;
  signal T1_27_i_14_n_0 : STD_LOGIC;
  signal T1_27_i_15_n_0 : STD_LOGIC;
  signal T1_27_i_16_n_0 : STD_LOGIC;
  signal T1_27_i_17_n_0 : STD_LOGIC;
  signal T1_27_i_18_n_0 : STD_LOGIC;
  signal T1_27_i_19_n_0 : STD_LOGIC;
  signal T1_27_i_20_n_0 : STD_LOGIC;
  signal T1_27_i_21_n_0 : STD_LOGIC;
  signal T1_27_i_22_n_0 : STD_LOGIC;
  signal T1_27_i_23_n_0 : STD_LOGIC;
  signal T1_27_i_24_n_0 : STD_LOGIC;
  signal T1_27_i_25_n_0 : STD_LOGIC;
  signal T1_27_i_26_n_0 : STD_LOGIC;
  signal T1_27_i_27_n_0 : STD_LOGIC;
  signal T1_27_i_29_n_0 : STD_LOGIC;
  signal T1_27_i_2_n_0 : STD_LOGIC;
  signal T1_27_i_30_n_0 : STD_LOGIC;
  signal T1_27_i_31_n_0 : STD_LOGIC;
  signal T1_27_i_32_n_0 : STD_LOGIC;
  signal T1_27_i_33_n_0 : STD_LOGIC;
  signal T1_27_i_34_n_0 : STD_LOGIC;
  signal T1_27_i_35_n_0 : STD_LOGIC;
  signal T1_27_i_36_n_0 : STD_LOGIC;
  signal T1_27_i_37_n_0 : STD_LOGIC;
  signal T1_27_i_38_n_0 : STD_LOGIC;
  signal T1_27_i_39_n_0 : STD_LOGIC;
  signal T1_27_i_3_n_0 : STD_LOGIC;
  signal T1_27_i_40_n_0 : STD_LOGIC;
  signal T1_27_i_41_n_0 : STD_LOGIC;
  signal T1_27_i_42_n_0 : STD_LOGIC;
  signal T1_27_i_43_n_0 : STD_LOGIC;
  signal T1_27_i_44_n_0 : STD_LOGIC;
  signal T1_27_i_45_n_0 : STD_LOGIC;
  signal T1_27_i_46_n_0 : STD_LOGIC;
  signal T1_27_i_49_n_0 : STD_LOGIC;
  signal T1_27_i_4_n_0 : STD_LOGIC;
  signal T1_27_i_50_n_0 : STD_LOGIC;
  signal T1_27_i_51_n_0 : STD_LOGIC;
  signal T1_27_i_52_n_0 : STD_LOGIC;
  signal T1_27_i_53_n_0 : STD_LOGIC;
  signal T1_27_i_54_n_0 : STD_LOGIC;
  signal T1_27_i_55_n_0 : STD_LOGIC;
  signal T1_27_i_56_n_0 : STD_LOGIC;
  signal T1_27_i_57_n_0 : STD_LOGIC;
  signal T1_27_i_58_n_0 : STD_LOGIC;
  signal T1_27_i_59_n_0 : STD_LOGIC;
  signal T1_27_i_5_n_0 : STD_LOGIC;
  signal T1_27_i_60_n_0 : STD_LOGIC;
  signal T1_27_i_61_n_0 : STD_LOGIC;
  signal T1_27_i_62_n_0 : STD_LOGIC;
  signal T1_27_i_63_n_0 : STD_LOGIC;
  signal T1_27_i_64_n_0 : STD_LOGIC;
  signal T1_27_i_65_n_0 : STD_LOGIC;
  signal T1_27_i_66_n_0 : STD_LOGIC;
  signal T1_27_i_67_n_0 : STD_LOGIC;
  signal T1_27_i_68_n_0 : STD_LOGIC;
  signal T1_27_i_69_n_0 : STD_LOGIC;
  signal T1_27_i_6_n_0 : STD_LOGIC;
  signal T1_27_i_70_n_0 : STD_LOGIC;
  signal T1_27_i_71_n_0 : STD_LOGIC;
  signal T1_27_i_72_n_0 : STD_LOGIC;
  signal T1_27_i_73_n_0 : STD_LOGIC;
  signal T1_27_i_74_n_0 : STD_LOGIC;
  signal T1_27_i_75_n_0 : STD_LOGIC;
  signal T1_27_i_76_n_0 : STD_LOGIC;
  signal T1_27_i_77_n_0 : STD_LOGIC;
  signal T1_27_i_78_n_0 : STD_LOGIC;
  signal T1_27_i_79_n_0 : STD_LOGIC;
  signal T1_27_i_7_n_0 : STD_LOGIC;
  signal T1_27_i_80_n_0 : STD_LOGIC;
  signal T1_27_i_81_n_0 : STD_LOGIC;
  signal T1_27_i_82_n_0 : STD_LOGIC;
  signal T1_27_i_83_n_0 : STD_LOGIC;
  signal T1_27_i_84_n_0 : STD_LOGIC;
  signal T1_27_i_85_n_0 : STD_LOGIC;
  signal T1_27_i_86_n_0 : STD_LOGIC;
  signal T1_27_i_87_n_0 : STD_LOGIC;
  signal T1_27_i_88_n_0 : STD_LOGIC;
  signal T1_27_i_89_n_0 : STD_LOGIC;
  signal T1_27_i_8_n_0 : STD_LOGIC;
  signal T1_27_i_90_n_0 : STD_LOGIC;
  signal T1_27_i_91_n_0 : STD_LOGIC;
  signal T1_27_i_92_n_0 : STD_LOGIC;
  signal T1_27_i_93_n_0 : STD_LOGIC;
  signal T1_27_i_94_n_0 : STD_LOGIC;
  signal T1_27_i_95_n_0 : STD_LOGIC;
  signal T1_27_i_96_n_0 : STD_LOGIC;
  signal T1_27_i_97_n_0 : STD_LOGIC;
  signal T1_27_i_98_n_0 : STD_LOGIC;
  signal T1_27_i_99_n_0 : STD_LOGIC;
  signal T1_27_i_9_n_0 : STD_LOGIC;
  signal T1_31_i_100_n_0 : STD_LOGIC;
  signal T1_31_i_101_n_0 : STD_LOGIC;
  signal T1_31_i_102_n_0 : STD_LOGIC;
  signal T1_31_i_103_n_0 : STD_LOGIC;
  signal T1_31_i_104_n_0 : STD_LOGIC;
  signal T1_31_i_105_n_0 : STD_LOGIC;
  signal T1_31_i_106_n_0 : STD_LOGIC;
  signal T1_31_i_107_n_0 : STD_LOGIC;
  signal T1_31_i_108_n_0 : STD_LOGIC;
  signal T1_31_i_109_n_0 : STD_LOGIC;
  signal T1_31_i_112_n_0 : STD_LOGIC;
  signal T1_31_i_113_n_0 : STD_LOGIC;
  signal T1_31_i_114_n_0 : STD_LOGIC;
  signal T1_31_i_115_n_0 : STD_LOGIC;
  signal T1_31_i_116_n_0 : STD_LOGIC;
  signal T1_31_i_117_n_0 : STD_LOGIC;
  signal T1_31_i_118_n_0 : STD_LOGIC;
  signal T1_31_i_119_n_0 : STD_LOGIC;
  signal T1_31_i_11_n_0 : STD_LOGIC;
  signal T1_31_i_128_n_0 : STD_LOGIC;
  signal T1_31_i_129_n_0 : STD_LOGIC;
  signal T1_31_i_12_n_0 : STD_LOGIC;
  signal T1_31_i_130_n_0 : STD_LOGIC;
  signal T1_31_i_131_n_0 : STD_LOGIC;
  signal T1_31_i_132_n_0 : STD_LOGIC;
  signal T1_31_i_133_n_0 : STD_LOGIC;
  signal T1_31_i_134_n_0 : STD_LOGIC;
  signal T1_31_i_135_n_0 : STD_LOGIC;
  signal T1_31_i_138_n_0 : STD_LOGIC;
  signal T1_31_i_139_n_0 : STD_LOGIC;
  signal T1_31_i_140_n_0 : STD_LOGIC;
  signal T1_31_i_141_n_0 : STD_LOGIC;
  signal T1_31_i_142_n_0 : STD_LOGIC;
  signal T1_31_i_143_n_0 : STD_LOGIC;
  signal T1_31_i_144_n_0 : STD_LOGIC;
  signal T1_31_i_145_n_0 : STD_LOGIC;
  signal T1_31_i_146_n_0 : STD_LOGIC;
  signal T1_31_i_147_n_0 : STD_LOGIC;
  signal T1_31_i_148_n_0 : STD_LOGIC;
  signal T1_31_i_149_n_0 : STD_LOGIC;
  signal T1_31_i_14_n_0 : STD_LOGIC;
  signal T1_31_i_152_n_0 : STD_LOGIC;
  signal T1_31_i_153_n_0 : STD_LOGIC;
  signal T1_31_i_154_n_0 : STD_LOGIC;
  signal T1_31_i_155_n_0 : STD_LOGIC;
  signal T1_31_i_156_n_0 : STD_LOGIC;
  signal T1_31_i_157_n_0 : STD_LOGIC;
  signal T1_31_i_158_n_0 : STD_LOGIC;
  signal T1_31_i_159_n_0 : STD_LOGIC;
  signal T1_31_i_15_n_0 : STD_LOGIC;
  signal T1_31_i_160_n_0 : STD_LOGIC;
  signal T1_31_i_161_n_0 : STD_LOGIC;
  signal T1_31_i_162_n_0 : STD_LOGIC;
  signal T1_31_i_163_n_0 : STD_LOGIC;
  signal T1_31_i_164_n_0 : STD_LOGIC;
  signal T1_31_i_165_n_0 : STD_LOGIC;
  signal T1_31_i_166_n_0 : STD_LOGIC;
  signal T1_31_i_167_n_0 : STD_LOGIC;
  signal T1_31_i_168_n_0 : STD_LOGIC;
  signal T1_31_i_169_n_0 : STD_LOGIC;
  signal T1_31_i_16_n_0 : STD_LOGIC;
  signal T1_31_i_170_n_0 : STD_LOGIC;
  signal T1_31_i_171_n_0 : STD_LOGIC;
  signal T1_31_i_172_n_0 : STD_LOGIC;
  signal T1_31_i_173_n_0 : STD_LOGIC;
  signal T1_31_i_174_n_0 : STD_LOGIC;
  signal T1_31_i_175_n_0 : STD_LOGIC;
  signal T1_31_i_176_n_0 : STD_LOGIC;
  signal T1_31_i_177_n_0 : STD_LOGIC;
  signal T1_31_i_178_n_0 : STD_LOGIC;
  signal T1_31_i_179_n_0 : STD_LOGIC;
  signal T1_31_i_17_n_0 : STD_LOGIC;
  signal T1_31_i_180_n_0 : STD_LOGIC;
  signal T1_31_i_181_n_0 : STD_LOGIC;
  signal T1_31_i_182_n_0 : STD_LOGIC;
  signal T1_31_i_183_n_0 : STD_LOGIC;
  signal T1_31_i_184_n_0 : STD_LOGIC;
  signal T1_31_i_185_n_0 : STD_LOGIC;
  signal T1_31_i_186_n_0 : STD_LOGIC;
  signal T1_31_i_187_n_0 : STD_LOGIC;
  signal T1_31_i_188_n_0 : STD_LOGIC;
  signal T1_31_i_189_n_0 : STD_LOGIC;
  signal T1_31_i_18_n_0 : STD_LOGIC;
  signal T1_31_i_190_n_0 : STD_LOGIC;
  signal T1_31_i_191_n_0 : STD_LOGIC;
  signal T1_31_i_192_n_0 : STD_LOGIC;
  signal T1_31_i_193_n_0 : STD_LOGIC;
  signal T1_31_i_194_n_0 : STD_LOGIC;
  signal T1_31_i_195_n_0 : STD_LOGIC;
  signal T1_31_i_196_n_0 : STD_LOGIC;
  signal T1_31_i_197_n_0 : STD_LOGIC;
  signal T1_31_i_198_n_0 : STD_LOGIC;
  signal T1_31_i_199_n_0 : STD_LOGIC;
  signal T1_31_i_19_n_0 : STD_LOGIC;
  signal T1_31_i_1_n_0 : STD_LOGIC;
  signal T1_31_i_200_n_0 : STD_LOGIC;
  signal T1_31_i_201_n_0 : STD_LOGIC;
  signal T1_31_i_202_n_0 : STD_LOGIC;
  signal T1_31_i_203_n_0 : STD_LOGIC;
  signal T1_31_i_204_n_0 : STD_LOGIC;
  signal T1_31_i_205_n_0 : STD_LOGIC;
  signal T1_31_i_206_n_0 : STD_LOGIC;
  signal T1_31_i_207_n_0 : STD_LOGIC;
  signal T1_31_i_208_n_0 : STD_LOGIC;
  signal T1_31_i_209_n_0 : STD_LOGIC;
  signal T1_31_i_20_n_0 : STD_LOGIC;
  signal T1_31_i_210_n_0 : STD_LOGIC;
  signal T1_31_i_211_n_0 : STD_LOGIC;
  signal T1_31_i_212_n_0 : STD_LOGIC;
  signal T1_31_i_213_n_0 : STD_LOGIC;
  signal T1_31_i_214_n_0 : STD_LOGIC;
  signal T1_31_i_215_n_0 : STD_LOGIC;
  signal T1_31_i_216_n_0 : STD_LOGIC;
  signal T1_31_i_217_n_0 : STD_LOGIC;
  signal T1_31_i_218_n_0 : STD_LOGIC;
  signal T1_31_i_219_n_0 : STD_LOGIC;
  signal T1_31_i_21_n_0 : STD_LOGIC;
  signal T1_31_i_220_n_0 : STD_LOGIC;
  signal T1_31_i_221_n_0 : STD_LOGIC;
  signal T1_31_i_222_n_0 : STD_LOGIC;
  signal T1_31_i_223_n_0 : STD_LOGIC;
  signal T1_31_i_224_n_0 : STD_LOGIC;
  signal T1_31_i_225_n_0 : STD_LOGIC;
  signal T1_31_i_226_n_0 : STD_LOGIC;
  signal T1_31_i_227_n_0 : STD_LOGIC;
  signal T1_31_i_228_n_0 : STD_LOGIC;
  signal T1_31_i_229_n_0 : STD_LOGIC;
  signal T1_31_i_22_n_0 : STD_LOGIC;
  signal T1_31_i_230_n_0 : STD_LOGIC;
  signal T1_31_i_231_n_0 : STD_LOGIC;
  signal T1_31_i_232_n_0 : STD_LOGIC;
  signal T1_31_i_233_n_0 : STD_LOGIC;
  signal T1_31_i_234_n_0 : STD_LOGIC;
  signal T1_31_i_235_n_0 : STD_LOGIC;
  signal T1_31_i_236_n_0 : STD_LOGIC;
  signal T1_31_i_237_n_0 : STD_LOGIC;
  signal T1_31_i_238_n_0 : STD_LOGIC;
  signal T1_31_i_239_n_0 : STD_LOGIC;
  signal T1_31_i_23_n_0 : STD_LOGIC;
  signal T1_31_i_24_n_0 : STD_LOGIC;
  signal T1_31_i_25_n_0 : STD_LOGIC;
  signal T1_31_i_26_n_0 : STD_LOGIC;
  signal T1_31_i_27_n_0 : STD_LOGIC;
  signal T1_31_i_28_n_0 : STD_LOGIC;
  signal T1_31_i_29_n_0 : STD_LOGIC;
  signal T1_31_i_30_n_0 : STD_LOGIC;
  signal T1_31_i_31_n_0 : STD_LOGIC;
  signal T1_31_i_32_n_0 : STD_LOGIC;
  signal T1_31_i_33_n_0 : STD_LOGIC;
  signal T1_31_i_34_n_0 : STD_LOGIC;
  signal T1_31_i_35_n_0 : STD_LOGIC;
  signal T1_31_i_36_n_0 : STD_LOGIC;
  signal T1_31_i_38_n_0 : STD_LOGIC;
  signal T1_31_i_39_n_0 : STD_LOGIC;
  signal T1_31_i_3_n_0 : STD_LOGIC;
  signal T1_31_i_40_n_0 : STD_LOGIC;
  signal T1_31_i_41_n_0 : STD_LOGIC;
  signal T1_31_i_42_n_0 : STD_LOGIC;
  signal T1_31_i_43_n_0 : STD_LOGIC;
  signal T1_31_i_44_n_0 : STD_LOGIC;
  signal T1_31_i_45_n_0 : STD_LOGIC;
  signal T1_31_i_46_n_0 : STD_LOGIC;
  signal T1_31_i_48_n_0 : STD_LOGIC;
  signal T1_31_i_49_n_0 : STD_LOGIC;
  signal T1_31_i_4_n_0 : STD_LOGIC;
  signal T1_31_i_50_n_0 : STD_LOGIC;
  signal T1_31_i_52_n_0 : STD_LOGIC;
  signal T1_31_i_53_n_0 : STD_LOGIC;
  signal T1_31_i_5_n_0 : STD_LOGIC;
  signal T1_31_i_60_n_0 : STD_LOGIC;
  signal T1_31_i_62_n_0 : STD_LOGIC;
  signal T1_31_i_63_n_0 : STD_LOGIC;
  signal T1_31_i_64_n_0 : STD_LOGIC;
  signal T1_31_i_66_n_0 : STD_LOGIC;
  signal T1_31_i_67_n_0 : STD_LOGIC;
  signal T1_31_i_68_n_0 : STD_LOGIC;
  signal T1_31_i_69_n_0 : STD_LOGIC;
  signal T1_31_i_6_n_0 : STD_LOGIC;
  signal T1_31_i_70_n_0 : STD_LOGIC;
  signal T1_31_i_71_n_0 : STD_LOGIC;
  signal T1_31_i_72_n_0 : STD_LOGIC;
  signal T1_31_i_73_n_0 : STD_LOGIC;
  signal T1_31_i_74_n_0 : STD_LOGIC;
  signal T1_31_i_75_n_0 : STD_LOGIC;
  signal T1_31_i_76_n_0 : STD_LOGIC;
  signal T1_31_i_77_n_0 : STD_LOGIC;
  signal T1_31_i_78_n_0 : STD_LOGIC;
  signal T1_31_i_79_n_0 : STD_LOGIC;
  signal T1_31_i_7_n_0 : STD_LOGIC;
  signal T1_31_i_80_n_0 : STD_LOGIC;
  signal T1_31_i_81_n_0 : STD_LOGIC;
  signal T1_31_i_82_n_0 : STD_LOGIC;
  signal T1_31_i_83_n_0 : STD_LOGIC;
  signal T1_31_i_84_n_0 : STD_LOGIC;
  signal T1_31_i_85_n_0 : STD_LOGIC;
  signal T1_31_i_86_n_0 : STD_LOGIC;
  signal T1_31_i_87_n_0 : STD_LOGIC;
  signal T1_31_i_88_n_0 : STD_LOGIC;
  signal T1_31_i_89_n_0 : STD_LOGIC;
  signal T1_31_i_8_n_0 : STD_LOGIC;
  signal T1_31_i_90_n_0 : STD_LOGIC;
  signal T1_31_i_91_n_0 : STD_LOGIC;
  signal T1_31_i_92_n_0 : STD_LOGIC;
  signal T1_31_i_93_n_0 : STD_LOGIC;
  signal T1_31_i_94_n_0 : STD_LOGIC;
  signal T1_31_i_95_n_0 : STD_LOGIC;
  signal T1_31_i_98_n_0 : STD_LOGIC;
  signal T1_31_i_99_n_0 : STD_LOGIC;
  signal T1_31_i_9_n_0 : STD_LOGIC;
  signal T1_3_i_10_n_0 : STD_LOGIC;
  signal T1_3_i_11_n_0 : STD_LOGIC;
  signal T1_3_i_2_n_0 : STD_LOGIC;
  signal T1_3_i_3_n_0 : STD_LOGIC;
  signal T1_3_i_4_n_0 : STD_LOGIC;
  signal T1_3_i_5_n_0 : STD_LOGIC;
  signal T1_3_i_6_n_0 : STD_LOGIC;
  signal T1_3_i_7_n_0 : STD_LOGIC;
  signal T1_3_i_8_n_0 : STD_LOGIC;
  signal T1_3_i_9_n_0 : STD_LOGIC;
  signal T1_7_i_10_n_0 : STD_LOGIC;
  signal T1_7_i_11_n_0 : STD_LOGIC;
  signal T1_7_i_12_n_0 : STD_LOGIC;
  signal T1_7_i_14_n_0 : STD_LOGIC;
  signal T1_7_i_15_n_0 : STD_LOGIC;
  signal T1_7_i_16_n_0 : STD_LOGIC;
  signal T1_7_i_17_n_0 : STD_LOGIC;
  signal T1_7_i_18_n_0 : STD_LOGIC;
  signal T1_7_i_19_n_0 : STD_LOGIC;
  signal T1_7_i_20_n_0 : STD_LOGIC;
  signal T1_7_i_21_n_0 : STD_LOGIC;
  signal T1_7_i_22_n_0 : STD_LOGIC;
  signal T1_7_i_23_n_0 : STD_LOGIC;
  signal T1_7_i_24_n_0 : STD_LOGIC;
  signal T1_7_i_25_n_0 : STD_LOGIC;
  signal T1_7_i_26_n_0 : STD_LOGIC;
  signal T1_7_i_27_n_0 : STD_LOGIC;
  signal T1_7_i_28_n_0 : STD_LOGIC;
  signal T1_7_i_29_n_0 : STD_LOGIC;
  signal T1_7_i_2_n_0 : STD_LOGIC;
  signal T1_7_i_30_n_0 : STD_LOGIC;
  signal T1_7_i_31_n_0 : STD_LOGIC;
  signal T1_7_i_32_n_0 : STD_LOGIC;
  signal T1_7_i_33_n_0 : STD_LOGIC;
  signal T1_7_i_34_n_0 : STD_LOGIC;
  signal T1_7_i_35_n_0 : STD_LOGIC;
  signal T1_7_i_36_n_0 : STD_LOGIC;
  signal T1_7_i_37_n_0 : STD_LOGIC;
  signal T1_7_i_38_n_0 : STD_LOGIC;
  signal T1_7_i_39_n_0 : STD_LOGIC;
  signal T1_7_i_3_n_0 : STD_LOGIC;
  signal T1_7_i_40_n_0 : STD_LOGIC;
  signal T1_7_i_41_n_0 : STD_LOGIC;
  signal T1_7_i_42_n_0 : STD_LOGIC;
  signal T1_7_i_43_n_0 : STD_LOGIC;
  signal T1_7_i_44_n_0 : STD_LOGIC;
  signal T1_7_i_45_n_0 : STD_LOGIC;
  signal T1_7_i_46_n_0 : STD_LOGIC;
  signal T1_7_i_47_n_0 : STD_LOGIC;
  signal T1_7_i_48_n_0 : STD_LOGIC;
  signal T1_7_i_49_n_0 : STD_LOGIC;
  signal T1_7_i_4_n_0 : STD_LOGIC;
  signal T1_7_i_50_n_0 : STD_LOGIC;
  signal T1_7_i_51_n_0 : STD_LOGIC;
  signal T1_7_i_52_n_0 : STD_LOGIC;
  signal T1_7_i_53_n_0 : STD_LOGIC;
  signal T1_7_i_54_n_0 : STD_LOGIC;
  signal T1_7_i_55_n_0 : STD_LOGIC;
  signal T1_7_i_56_n_0 : STD_LOGIC;
  signal T1_7_i_57_n_0 : STD_LOGIC;
  signal T1_7_i_58_n_0 : STD_LOGIC;
  signal T1_7_i_59_n_0 : STD_LOGIC;
  signal T1_7_i_5_n_0 : STD_LOGIC;
  signal T1_7_i_60_n_0 : STD_LOGIC;
  signal T1_7_i_61_n_0 : STD_LOGIC;
  signal T1_7_i_62_n_0 : STD_LOGIC;
  signal T1_7_i_63_n_0 : STD_LOGIC;
  signal T1_7_i_64_n_0 : STD_LOGIC;
  signal T1_7_i_65_n_0 : STD_LOGIC;
  signal T1_7_i_66_n_0 : STD_LOGIC;
  signal T1_7_i_67_n_0 : STD_LOGIC;
  signal T1_7_i_68_n_0 : STD_LOGIC;
  signal T1_7_i_69_n_0 : STD_LOGIC;
  signal T1_7_i_6_n_0 : STD_LOGIC;
  signal T1_7_i_70_n_0 : STD_LOGIC;
  signal T1_7_i_71_n_0 : STD_LOGIC;
  signal T1_7_i_72_n_0 : STD_LOGIC;
  signal T1_7_i_73_n_0 : STD_LOGIC;
  signal T1_7_i_74_n_0 : STD_LOGIC;
  signal T1_7_i_75_n_0 : STD_LOGIC;
  signal T1_7_i_76_n_0 : STD_LOGIC;
  signal T1_7_i_77_n_0 : STD_LOGIC;
  signal T1_7_i_78_n_0 : STD_LOGIC;
  signal T1_7_i_79_n_0 : STD_LOGIC;
  signal T1_7_i_7_n_0 : STD_LOGIC;
  signal T1_7_i_80_n_0 : STD_LOGIC;
  signal T1_7_i_81_n_0 : STD_LOGIC;
  signal T1_7_i_82_n_0 : STD_LOGIC;
  signal T1_7_i_83_n_0 : STD_LOGIC;
  signal T1_7_i_84_n_0 : STD_LOGIC;
  signal T1_7_i_8_n_0 : STD_LOGIC;
  signal T1_7_i_9_n_0 : STD_LOGIC;
  signal T1_reg_11_i_13_n_0 : STD_LOGIC;
  signal T1_reg_11_i_13_n_1 : STD_LOGIC;
  signal T1_reg_11_i_13_n_2 : STD_LOGIC;
  signal T1_reg_11_i_13_n_3 : STD_LOGIC;
  signal T1_reg_11_i_13_n_4 : STD_LOGIC;
  signal T1_reg_11_i_13_n_5 : STD_LOGIC;
  signal T1_reg_11_i_13_n_6 : STD_LOGIC;
  signal T1_reg_11_i_13_n_7 : STD_LOGIC;
  signal T1_reg_11_i_1_n_0 : STD_LOGIC;
  signal T1_reg_11_i_1_n_1 : STD_LOGIC;
  signal T1_reg_11_i_1_n_2 : STD_LOGIC;
  signal T1_reg_11_i_1_n_3 : STD_LOGIC;
  signal T1_reg_15_i_13_n_0 : STD_LOGIC;
  signal T1_reg_15_i_13_n_1 : STD_LOGIC;
  signal T1_reg_15_i_13_n_2 : STD_LOGIC;
  signal T1_reg_15_i_13_n_3 : STD_LOGIC;
  signal T1_reg_15_i_13_n_4 : STD_LOGIC;
  signal T1_reg_15_i_13_n_5 : STD_LOGIC;
  signal T1_reg_15_i_13_n_6 : STD_LOGIC;
  signal T1_reg_15_i_13_n_7 : STD_LOGIC;
  signal T1_reg_15_i_1_n_0 : STD_LOGIC;
  signal T1_reg_15_i_1_n_1 : STD_LOGIC;
  signal T1_reg_15_i_1_n_2 : STD_LOGIC;
  signal T1_reg_15_i_1_n_3 : STD_LOGIC;
  signal T1_reg_15_i_29_n_0 : STD_LOGIC;
  signal T1_reg_15_i_33_n_0 : STD_LOGIC;
  signal T1_reg_15_i_37_n_0 : STD_LOGIC;
  signal T1_reg_15_i_51_n_0 : STD_LOGIC;
  signal T1_reg_15_i_52_n_0 : STD_LOGIC;
  signal T1_reg_15_i_65_n_0 : STD_LOGIC;
  signal T1_reg_15_i_66_n_0 : STD_LOGIC;
  signal T1_reg_15_i_79_n_0 : STD_LOGIC;
  signal T1_reg_15_i_80_n_0 : STD_LOGIC;
  signal T1_reg_19_i_100_n_0 : STD_LOGIC;
  signal T1_reg_19_i_13_n_0 : STD_LOGIC;
  signal T1_reg_19_i_13_n_1 : STD_LOGIC;
  signal T1_reg_19_i_13_n_2 : STD_LOGIC;
  signal T1_reg_19_i_13_n_3 : STD_LOGIC;
  signal T1_reg_19_i_13_n_4 : STD_LOGIC;
  signal T1_reg_19_i_13_n_5 : STD_LOGIC;
  signal T1_reg_19_i_13_n_6 : STD_LOGIC;
  signal T1_reg_19_i_13_n_7 : STD_LOGIC;
  signal T1_reg_19_i_1_n_0 : STD_LOGIC;
  signal T1_reg_19_i_1_n_1 : STD_LOGIC;
  signal T1_reg_19_i_1_n_2 : STD_LOGIC;
  signal T1_reg_19_i_1_n_3 : STD_LOGIC;
  signal T1_reg_19_i_41_n_0 : STD_LOGIC;
  signal T1_reg_19_i_99_n_0 : STD_LOGIC;
  signal T1_reg_23_i_13_n_0 : STD_LOGIC;
  signal T1_reg_23_i_13_n_1 : STD_LOGIC;
  signal T1_reg_23_i_13_n_2 : STD_LOGIC;
  signal T1_reg_23_i_13_n_3 : STD_LOGIC;
  signal T1_reg_23_i_13_n_4 : STD_LOGIC;
  signal T1_reg_23_i_13_n_5 : STD_LOGIC;
  signal T1_reg_23_i_13_n_6 : STD_LOGIC;
  signal T1_reg_23_i_13_n_7 : STD_LOGIC;
  signal T1_reg_23_i_1_n_0 : STD_LOGIC;
  signal T1_reg_23_i_1_n_1 : STD_LOGIC;
  signal T1_reg_23_i_1_n_2 : STD_LOGIC;
  signal T1_reg_23_i_1_n_3 : STD_LOGIC;
  signal T1_reg_23_i_40_n_0 : STD_LOGIC;
  signal T1_reg_23_i_95_n_0 : STD_LOGIC;
  signal T1_reg_23_i_96_n_0 : STD_LOGIC;
  signal T1_reg_27_i_13_n_0 : STD_LOGIC;
  signal T1_reg_27_i_13_n_1 : STD_LOGIC;
  signal T1_reg_27_i_13_n_2 : STD_LOGIC;
  signal T1_reg_27_i_13_n_3 : STD_LOGIC;
  signal T1_reg_27_i_13_n_4 : STD_LOGIC;
  signal T1_reg_27_i_13_n_5 : STD_LOGIC;
  signal T1_reg_27_i_13_n_6 : STD_LOGIC;
  signal T1_reg_27_i_13_n_7 : STD_LOGIC;
  signal T1_reg_27_i_1_n_0 : STD_LOGIC;
  signal T1_reg_27_i_1_n_1 : STD_LOGIC;
  signal T1_reg_27_i_1_n_2 : STD_LOGIC;
  signal T1_reg_27_i_1_n_3 : STD_LOGIC;
  signal T1_reg_27_i_28_n_0 : STD_LOGIC;
  signal T1_reg_27_i_47_n_0 : STD_LOGIC;
  signal T1_reg_27_i_48_n_0 : STD_LOGIC;
  signal T1_reg_31_i_10_n_1 : STD_LOGIC;
  signal T1_reg_31_i_10_n_2 : STD_LOGIC;
  signal T1_reg_31_i_10_n_3 : STD_LOGIC;
  signal T1_reg_31_i_10_n_4 : STD_LOGIC;
  signal T1_reg_31_i_10_n_5 : STD_LOGIC;
  signal T1_reg_31_i_10_n_6 : STD_LOGIC;
  signal T1_reg_31_i_10_n_7 : STD_LOGIC;
  signal T1_reg_31_i_110_n_0 : STD_LOGIC;
  signal T1_reg_31_i_111_n_0 : STD_LOGIC;
  signal T1_reg_31_i_120_n_0 : STD_LOGIC;
  signal T1_reg_31_i_121_n_0 : STD_LOGIC;
  signal T1_reg_31_i_122_n_0 : STD_LOGIC;
  signal T1_reg_31_i_123_n_0 : STD_LOGIC;
  signal T1_reg_31_i_124_n_0 : STD_LOGIC;
  signal T1_reg_31_i_125_n_0 : STD_LOGIC;
  signal T1_reg_31_i_126_n_0 : STD_LOGIC;
  signal T1_reg_31_i_127_n_0 : STD_LOGIC;
  signal T1_reg_31_i_136_n_0 : STD_LOGIC;
  signal T1_reg_31_i_137_n_0 : STD_LOGIC;
  signal T1_reg_31_i_13_n_0 : STD_LOGIC;
  signal T1_reg_31_i_13_n_1 : STD_LOGIC;
  signal T1_reg_31_i_13_n_2 : STD_LOGIC;
  signal T1_reg_31_i_13_n_3 : STD_LOGIC;
  signal T1_reg_31_i_13_n_4 : STD_LOGIC;
  signal T1_reg_31_i_13_n_5 : STD_LOGIC;
  signal T1_reg_31_i_13_n_6 : STD_LOGIC;
  signal T1_reg_31_i_13_n_7 : STD_LOGIC;
  signal T1_reg_31_i_150_n_0 : STD_LOGIC;
  signal T1_reg_31_i_151_n_0 : STD_LOGIC;
  signal T1_reg_31_i_2_n_1 : STD_LOGIC;
  signal T1_reg_31_i_2_n_2 : STD_LOGIC;
  signal T1_reg_31_i_2_n_3 : STD_LOGIC;
  signal T1_reg_31_i_37_n_0 : STD_LOGIC;
  signal T1_reg_31_i_47_n_0 : STD_LOGIC;
  signal T1_reg_31_i_51_n_0 : STD_LOGIC;
  signal T1_reg_31_i_54_n_0 : STD_LOGIC;
  signal T1_reg_31_i_55_n_0 : STD_LOGIC;
  signal T1_reg_31_i_56_n_0 : STD_LOGIC;
  signal T1_reg_31_i_57_n_0 : STD_LOGIC;
  signal T1_reg_31_i_58_n_0 : STD_LOGIC;
  signal T1_reg_31_i_59_n_0 : STD_LOGIC;
  signal T1_reg_31_i_61_n_0 : STD_LOGIC;
  signal T1_reg_31_i_65_n_0 : STD_LOGIC;
  signal T1_reg_31_i_96_n_0 : STD_LOGIC;
  signal T1_reg_31_i_97_n_0 : STD_LOGIC;
  signal T1_reg_3_i_1_n_0 : STD_LOGIC;
  signal T1_reg_3_i_1_n_1 : STD_LOGIC;
  signal T1_reg_3_i_1_n_2 : STD_LOGIC;
  signal T1_reg_3_i_1_n_3 : STD_LOGIC;
  signal T1_reg_7_i_13_n_0 : STD_LOGIC;
  signal T1_reg_7_i_13_n_1 : STD_LOGIC;
  signal T1_reg_7_i_13_n_2 : STD_LOGIC;
  signal T1_reg_7_i_13_n_3 : STD_LOGIC;
  signal T1_reg_7_i_13_n_4 : STD_LOGIC;
  signal T1_reg_7_i_13_n_5 : STD_LOGIC;
  signal T1_reg_7_i_13_n_6 : STD_LOGIC;
  signal T1_reg_7_i_13_n_7 : STD_LOGIC;
  signal T1_reg_7_i_1_n_0 : STD_LOGIC;
  signal T1_reg_7_i_1_n_1 : STD_LOGIC;
  signal T1_reg_7_i_1_n_2 : STD_LOGIC;
  signal T1_reg_7_i_1_n_3 : STD_LOGIC;
  signal T1_0_31 : STD_LOGIC;
  signal T1_0_30 : STD_LOGIC;
  signal T1_0_29 : STD_LOGIC;
  signal T1_0_28 : STD_LOGIC;
  signal T1_0_27 : STD_LOGIC;
  signal T1_0_26 : STD_LOGIC;
  signal T1_0_25 : STD_LOGIC;
  signal T1_0_24 : STD_LOGIC;
  signal T1_0_23 : STD_LOGIC;
  signal T1_0_22 : STD_LOGIC;
  signal T1_0_21 : STD_LOGIC;
  signal T1_0_20 : STD_LOGIC;
  signal T1_0_19 : STD_LOGIC;
  signal T1_0_18 : STD_LOGIC;
  signal T1_0_17 : STD_LOGIC;
  signal T1_0_16 : STD_LOGIC;
  signal T1_0_15 : STD_LOGIC;
  signal T1_0_14 : STD_LOGIC;
  signal T1_0_13 : STD_LOGIC;
  signal T1_0_12 : STD_LOGIC;
  signal T1_0_11 : STD_LOGIC;
  signal T1_0_10 : STD_LOGIC;
  signal T1_0_9 : STD_LOGIC;
  signal T1_0_8 : STD_LOGIC;
  signal T1_0_7 : STD_LOGIC;
  signal T1_0_6 : STD_LOGIC;
  signal T1_0_5 : STD_LOGIC;
  signal T1_0_4 : STD_LOGIC;
  signal T1_0_3 : STD_LOGIC;
  signal T1_0_2 : STD_LOGIC;
  signal T1_0_1 : STD_LOGIC;
  signal T1_0_0 : STD_LOGIC;
  signal T2_31 : STD_LOGIC;
  signal T2_30 : STD_LOGIC;
  signal T2_29 : STD_LOGIC;
  signal T2_28 : STD_LOGIC;
  signal T2_27 : STD_LOGIC;
  signal T2_26 : STD_LOGIC;
  signal T2_25 : STD_LOGIC;
  signal T2_24 : STD_LOGIC;
  signal T2_23 : STD_LOGIC;
  signal T2_22 : STD_LOGIC;
  signal T2_21 : STD_LOGIC;
  signal T2_20 : STD_LOGIC;
  signal T2_19 : STD_LOGIC;
  signal T2_18 : STD_LOGIC;
  signal T2_17 : STD_LOGIC;
  signal T2_16 : STD_LOGIC;
  signal T2_15 : STD_LOGIC;
  signal T2_14 : STD_LOGIC;
  signal T2_13 : STD_LOGIC;
  signal T2_12 : STD_LOGIC;
  signal T2_11 : STD_LOGIC;
  signal T2_10 : STD_LOGIC;
  signal T2_9 : STD_LOGIC;
  signal T2_8 : STD_LOGIC;
  signal T2_7 : STD_LOGIC;
  signal T2_6 : STD_LOGIC;
  signal T2_5 : STD_LOGIC;
  signal T2_4 : STD_LOGIC;
  signal T2_3 : STD_LOGIC;
  signal T2_2 : STD_LOGIC;
  signal T2_1 : STD_LOGIC;
  signal T2_0 : STD_LOGIC;
  signal T20_31 : STD_LOGIC;
  signal T20_30 : STD_LOGIC;
  signal T20_29 : STD_LOGIC;
  signal T20_28 : STD_LOGIC;
  signal T20_27 : STD_LOGIC;
  signal T20_26 : STD_LOGIC;
  signal T20_25 : STD_LOGIC;
  signal T20_24 : STD_LOGIC;
  signal T20_23 : STD_LOGIC;
  signal T20_22 : STD_LOGIC;
  signal T20_21 : STD_LOGIC;
  signal T20_20 : STD_LOGIC;
  signal T20_19 : STD_LOGIC;
  signal T20_18 : STD_LOGIC;
  signal T20_17 : STD_LOGIC;
  signal T20_16 : STD_LOGIC;
  signal T20_15 : STD_LOGIC;
  signal T20_14 : STD_LOGIC;
  signal T20_13 : STD_LOGIC;
  signal T20_12 : STD_LOGIC;
  signal T20_11 : STD_LOGIC;
  signal T20_10 : STD_LOGIC;
  signal T20_9 : STD_LOGIC;
  signal T20_8 : STD_LOGIC;
  signal T20_7 : STD_LOGIC;
  signal T20_6 : STD_LOGIC;
  signal T20_5 : STD_LOGIC;
  signal T20_4 : STD_LOGIC;
  signal T20_3 : STD_LOGIC;
  signal T20_2 : STD_LOGIC;
  signal T20_1 : STD_LOGIC;
  signal T20_0 : STD_LOGIC;
  signal T2_11_i_6_n_0 : STD_LOGIC;
  signal T2_11_i_7_n_0 : STD_LOGIC;
  signal T2_11_i_8_n_0 : STD_LOGIC;
  signal T2_11_i_9_n_0 : STD_LOGIC;
  signal T2_15_i_6_n_0 : STD_LOGIC;
  signal T2_15_i_7_n_0 : STD_LOGIC;
  signal T2_15_i_8_n_0 : STD_LOGIC;
  signal T2_15_i_9_n_0 : STD_LOGIC;
  signal T2_19_i_6_n_0 : STD_LOGIC;
  signal T2_19_i_7_n_0 : STD_LOGIC;
  signal T2_19_i_8_n_0 : STD_LOGIC;
  signal T2_19_i_9_n_0 : STD_LOGIC;
  signal T2_23_i_6_n_0 : STD_LOGIC;
  signal T2_23_i_7_n_0 : STD_LOGIC;
  signal T2_23_i_8_n_0 : STD_LOGIC;
  signal T2_23_i_9_n_0 : STD_LOGIC;
  signal T2_27_i_6_n_0 : STD_LOGIC;
  signal T2_27_i_7_n_0 : STD_LOGIC;
  signal T2_27_i_8_n_0 : STD_LOGIC;
  signal T2_27_i_9_n_0 : STD_LOGIC;
  signal T2_31_i_5_n_0 : STD_LOGIC;
  signal T2_31_i_6_n_0 : STD_LOGIC;
  signal T2_31_i_7_n_0 : STD_LOGIC;
  signal T2_31_i_8_n_0 : STD_LOGIC;
  signal T2_3_i_6_n_0 : STD_LOGIC;
  signal T2_3_i_7_n_0 : STD_LOGIC;
  signal T2_3_i_8_n_0 : STD_LOGIC;
  signal T2_3_i_9_n_0 : STD_LOGIC;
  signal T2_7_i_6_n_0 : STD_LOGIC;
  signal T2_7_i_7_n_0 : STD_LOGIC;
  signal T2_7_i_8_n_0 : STD_LOGIC;
  signal T2_7_i_9_n_0 : STD_LOGIC;
  signal T2_reg_11_i_1_n_0 : STD_LOGIC;
  signal T2_reg_11_i_1_n_1 : STD_LOGIC;
  signal T2_reg_11_i_1_n_2 : STD_LOGIC;
  signal T2_reg_11_i_1_n_3 : STD_LOGIC;
  signal T2_reg_15_i_1_n_0 : STD_LOGIC;
  signal T2_reg_15_i_1_n_1 : STD_LOGIC;
  signal T2_reg_15_i_1_n_2 : STD_LOGIC;
  signal T2_reg_15_i_1_n_3 : STD_LOGIC;
  signal T2_reg_19_i_1_n_0 : STD_LOGIC;
  signal T2_reg_19_i_1_n_1 : STD_LOGIC;
  signal T2_reg_19_i_1_n_2 : STD_LOGIC;
  signal T2_reg_19_i_1_n_3 : STD_LOGIC;
  signal T2_reg_23_i_1_n_0 : STD_LOGIC;
  signal T2_reg_23_i_1_n_1 : STD_LOGIC;
  signal T2_reg_23_i_1_n_2 : STD_LOGIC;
  signal T2_reg_23_i_1_n_3 : STD_LOGIC;
  signal T2_reg_27_i_1_n_0 : STD_LOGIC;
  signal T2_reg_27_i_1_n_1 : STD_LOGIC;
  signal T2_reg_27_i_1_n_2 : STD_LOGIC;
  signal T2_reg_27_i_1_n_3 : STD_LOGIC;
  signal T2_reg_31_i_1_n_1 : STD_LOGIC;
  signal T2_reg_31_i_1_n_2 : STD_LOGIC;
  signal T2_reg_31_i_1_n_3 : STD_LOGIC;
  signal T2_reg_3_i_1_n_0 : STD_LOGIC;
  signal T2_reg_3_i_1_n_1 : STD_LOGIC;
  signal T2_reg_3_i_1_n_2 : STD_LOGIC;
  signal T2_reg_3_i_1_n_3 : STD_LOGIC;
  signal T2_reg_7_i_1_n_0 : STD_LOGIC;
  signal T2_reg_7_i_1_n_1 : STD_LOGIC;
  signal T2_reg_7_i_1_n_2 : STD_LOGIC;
  signal T2_reg_7_i_1_n_3 : STD_LOGIC;
  signal W_0 : STD_LOGIC;
  signal W_16 : STD_LOGIC;
  signal W_16_11_i_10_n_0 : STD_LOGIC;
  signal W_16_11_i_11_n_0 : STD_LOGIC;
  signal W_16_11_i_12_n_0 : STD_LOGIC;
  signal W_16_11_i_13_n_0 : STD_LOGIC;
  signal W_16_11_i_14_n_0 : STD_LOGIC;
  signal W_16_11_i_15_n_0 : STD_LOGIC;
  signal W_16_11_i_16_n_0 : STD_LOGIC;
  signal W_16_11_i_17_n_0 : STD_LOGIC;
  signal W_16_11_i_2_n_0 : STD_LOGIC;
  signal W_16_11_i_3_n_0 : STD_LOGIC;
  signal W_16_11_i_4_n_0 : STD_LOGIC;
  signal W_16_11_i_5_n_0 : STD_LOGIC;
  signal W_16_11_i_6_n_0 : STD_LOGIC;
  signal W_16_11_i_7_n_0 : STD_LOGIC;
  signal W_16_11_i_8_n_0 : STD_LOGIC;
  signal W_16_11_i_9_n_0 : STD_LOGIC;
  signal W_16_15_i_10_n_0 : STD_LOGIC;
  signal W_16_15_i_11_n_0 : STD_LOGIC;
  signal W_16_15_i_12_n_0 : STD_LOGIC;
  signal W_16_15_i_13_n_0 : STD_LOGIC;
  signal W_16_15_i_14_n_0 : STD_LOGIC;
  signal W_16_15_i_15_n_0 : STD_LOGIC;
  signal W_16_15_i_16_n_0 : STD_LOGIC;
  signal W_16_15_i_17_n_0 : STD_LOGIC;
  signal W_16_15_i_2_n_0 : STD_LOGIC;
  signal W_16_15_i_3_n_0 : STD_LOGIC;
  signal W_16_15_i_4_n_0 : STD_LOGIC;
  signal W_16_15_i_5_n_0 : STD_LOGIC;
  signal W_16_15_i_6_n_0 : STD_LOGIC;
  signal W_16_15_i_7_n_0 : STD_LOGIC;
  signal W_16_15_i_8_n_0 : STD_LOGIC;
  signal W_16_15_i_9_n_0 : STD_LOGIC;
  signal W_16_19_i_10_n_0 : STD_LOGIC;
  signal W_16_19_i_11_n_0 : STD_LOGIC;
  signal W_16_19_i_12_n_0 : STD_LOGIC;
  signal W_16_19_i_13_n_0 : STD_LOGIC;
  signal W_16_19_i_14_n_0 : STD_LOGIC;
  signal W_16_19_i_15_n_0 : STD_LOGIC;
  signal W_16_19_i_16_n_0 : STD_LOGIC;
  signal W_16_19_i_17_n_0 : STD_LOGIC;
  signal W_16_19_i_2_n_0 : STD_LOGIC;
  signal W_16_19_i_3_n_0 : STD_LOGIC;
  signal W_16_19_i_4_n_0 : STD_LOGIC;
  signal W_16_19_i_5_n_0 : STD_LOGIC;
  signal W_16_19_i_6_n_0 : STD_LOGIC;
  signal W_16_19_i_7_n_0 : STD_LOGIC;
  signal W_16_19_i_8_n_0 : STD_LOGIC;
  signal W_16_19_i_9_n_0 : STD_LOGIC;
  signal W_16_23_i_10_n_0 : STD_LOGIC;
  signal W_16_23_i_11_n_0 : STD_LOGIC;
  signal W_16_23_i_12_n_0 : STD_LOGIC;
  signal W_16_23_i_13_n_0 : STD_LOGIC;
  signal W_16_23_i_14_n_0 : STD_LOGIC;
  signal W_16_23_i_15_n_0 : STD_LOGIC;
  signal W_16_23_i_16_n_0 : STD_LOGIC;
  signal W_16_23_i_17_n_0 : STD_LOGIC;
  signal W_16_23_i_2_n_0 : STD_LOGIC;
  signal W_16_23_i_3_n_0 : STD_LOGIC;
  signal W_16_23_i_4_n_0 : STD_LOGIC;
  signal W_16_23_i_5_n_0 : STD_LOGIC;
  signal W_16_23_i_6_n_0 : STD_LOGIC;
  signal W_16_23_i_7_n_0 : STD_LOGIC;
  signal W_16_23_i_8_n_0 : STD_LOGIC;
  signal W_16_23_i_9_n_0 : STD_LOGIC;
  signal W_16_27_i_10_n_0 : STD_LOGIC;
  signal W_16_27_i_11_n_0 : STD_LOGIC;
  signal W_16_27_i_12_n_0 : STD_LOGIC;
  signal W_16_27_i_13_n_0 : STD_LOGIC;
  signal W_16_27_i_14_n_0 : STD_LOGIC;
  signal W_16_27_i_15_n_0 : STD_LOGIC;
  signal W_16_27_i_16_n_0 : STD_LOGIC;
  signal W_16_27_i_17_n_0 : STD_LOGIC;
  signal W_16_27_i_2_n_0 : STD_LOGIC;
  signal W_16_27_i_3_n_0 : STD_LOGIC;
  signal W_16_27_i_4_n_0 : STD_LOGIC;
  signal W_16_27_i_5_n_0 : STD_LOGIC;
  signal W_16_27_i_6_n_0 : STD_LOGIC;
  signal W_16_27_i_7_n_0 : STD_LOGIC;
  signal W_16_27_i_8_n_0 : STD_LOGIC;
  signal W_16_27_i_9_n_0 : STD_LOGIC;
  signal W_16_31_i_10_n_0 : STD_LOGIC;
  signal W_16_31_i_11_n_0 : STD_LOGIC;
  signal W_16_31_i_12_n_0 : STD_LOGIC;
  signal W_16_31_i_13_n_0 : STD_LOGIC;
  signal W_16_31_i_14_n_0 : STD_LOGIC;
  signal W_16_31_i_15_n_0 : STD_LOGIC;
  signal W_16_31_i_16_n_0 : STD_LOGIC;
  signal W_16_31_i_18_n_0 : STD_LOGIC;
  signal W_16_31_i_20_n_0 : STD_LOGIC;
  signal W_16_31_i_3_n_0 : STD_LOGIC;
  signal W_16_31_i_4_n_0 : STD_LOGIC;
  signal W_16_31_i_5_n_0 : STD_LOGIC;
  signal W_16_31_i_6_n_0 : STD_LOGIC;
  signal W_16_31_i_7_n_0 : STD_LOGIC;
  signal W_16_31_i_8_n_0 : STD_LOGIC;
  signal W_16_31_i_9_n_0 : STD_LOGIC;
  signal W_16_3_i_10_n_0 : STD_LOGIC;
  signal W_16_3_i_11_n_0 : STD_LOGIC;
  signal W_16_3_i_13_n_0 : STD_LOGIC;
  signal W_16_3_i_2_n_0 : STD_LOGIC;
  signal W_16_3_i_3_n_0 : STD_LOGIC;
  signal W_16_3_i_4_n_0 : STD_LOGIC;
  signal W_16_3_i_5_n_0 : STD_LOGIC;
  signal W_16_3_i_6_n_0 : STD_LOGIC;
  signal W_16_3_i_7_n_0 : STD_LOGIC;
  signal W_16_3_i_8_n_0 : STD_LOGIC;
  signal W_16_3_i_9_n_0 : STD_LOGIC;
  signal W_16_7_i_10_n_0 : STD_LOGIC;
  signal W_16_7_i_11_n_0 : STD_LOGIC;
  signal W_16_7_i_12_n_0 : STD_LOGIC;
  signal W_16_7_i_13_n_0 : STD_LOGIC;
  signal W_16_7_i_14_n_0 : STD_LOGIC;
  signal W_16_7_i_15_n_0 : STD_LOGIC;
  signal W_16_7_i_16_n_0 : STD_LOGIC;
  signal W_16_7_i_17_n_0 : STD_LOGIC;
  signal W_16_7_i_2_n_0 : STD_LOGIC;
  signal W_16_7_i_3_n_0 : STD_LOGIC;
  signal W_16_7_i_4_n_0 : STD_LOGIC;
  signal W_16_7_i_5_n_0 : STD_LOGIC;
  signal W_16_7_i_6_n_0 : STD_LOGIC;
  signal W_16_7_i_7_n_0 : STD_LOGIC;
  signal W_16_7_i_8_n_0 : STD_LOGIC;
  signal W_16_7_i_9_n_0 : STD_LOGIC;
  signal W_17_11_i_10_n_0 : STD_LOGIC;
  signal W_17_11_i_11_n_0 : STD_LOGIC;
  signal W_17_11_i_12_n_0 : STD_LOGIC;
  signal W_17_11_i_13_n_0 : STD_LOGIC;
  signal W_17_11_i_14_n_0 : STD_LOGIC;
  signal W_17_11_i_15_n_0 : STD_LOGIC;
  signal W_17_11_i_16_n_0 : STD_LOGIC;
  signal W_17_11_i_17_n_0 : STD_LOGIC;
  signal W_17_11_i_2_n_0 : STD_LOGIC;
  signal W_17_11_i_3_n_0 : STD_LOGIC;
  signal W_17_11_i_4_n_0 : STD_LOGIC;
  signal W_17_11_i_5_n_0 : STD_LOGIC;
  signal W_17_11_i_6_n_0 : STD_LOGIC;
  signal W_17_11_i_7_n_0 : STD_LOGIC;
  signal W_17_11_i_8_n_0 : STD_LOGIC;
  signal W_17_11_i_9_n_0 : STD_LOGIC;
  signal W_17_15_i_10_n_0 : STD_LOGIC;
  signal W_17_15_i_11_n_0 : STD_LOGIC;
  signal W_17_15_i_12_n_0 : STD_LOGIC;
  signal W_17_15_i_13_n_0 : STD_LOGIC;
  signal W_17_15_i_14_n_0 : STD_LOGIC;
  signal W_17_15_i_15_n_0 : STD_LOGIC;
  signal W_17_15_i_16_n_0 : STD_LOGIC;
  signal W_17_15_i_17_n_0 : STD_LOGIC;
  signal W_17_15_i_2_n_0 : STD_LOGIC;
  signal W_17_15_i_3_n_0 : STD_LOGIC;
  signal W_17_15_i_4_n_0 : STD_LOGIC;
  signal W_17_15_i_5_n_0 : STD_LOGIC;
  signal W_17_15_i_6_n_0 : STD_LOGIC;
  signal W_17_15_i_7_n_0 : STD_LOGIC;
  signal W_17_15_i_8_n_0 : STD_LOGIC;
  signal W_17_15_i_9_n_0 : STD_LOGIC;
  signal W_17_19_i_10_n_0 : STD_LOGIC;
  signal W_17_19_i_11_n_0 : STD_LOGIC;
  signal W_17_19_i_12_n_0 : STD_LOGIC;
  signal W_17_19_i_13_n_0 : STD_LOGIC;
  signal W_17_19_i_14_n_0 : STD_LOGIC;
  signal W_17_19_i_15_n_0 : STD_LOGIC;
  signal W_17_19_i_16_n_0 : STD_LOGIC;
  signal W_17_19_i_17_n_0 : STD_LOGIC;
  signal W_17_19_i_2_n_0 : STD_LOGIC;
  signal W_17_19_i_3_n_0 : STD_LOGIC;
  signal W_17_19_i_4_n_0 : STD_LOGIC;
  signal W_17_19_i_5_n_0 : STD_LOGIC;
  signal W_17_19_i_6_n_0 : STD_LOGIC;
  signal W_17_19_i_7_n_0 : STD_LOGIC;
  signal W_17_19_i_8_n_0 : STD_LOGIC;
  signal W_17_19_i_9_n_0 : STD_LOGIC;
  signal W_17_23_i_10_n_0 : STD_LOGIC;
  signal W_17_23_i_11_n_0 : STD_LOGIC;
  signal W_17_23_i_12_n_0 : STD_LOGIC;
  signal W_17_23_i_13_n_0 : STD_LOGIC;
  signal W_17_23_i_14_n_0 : STD_LOGIC;
  signal W_17_23_i_15_n_0 : STD_LOGIC;
  signal W_17_23_i_16_n_0 : STD_LOGIC;
  signal W_17_23_i_17_n_0 : STD_LOGIC;
  signal W_17_23_i_2_n_0 : STD_LOGIC;
  signal W_17_23_i_3_n_0 : STD_LOGIC;
  signal W_17_23_i_4_n_0 : STD_LOGIC;
  signal W_17_23_i_5_n_0 : STD_LOGIC;
  signal W_17_23_i_6_n_0 : STD_LOGIC;
  signal W_17_23_i_7_n_0 : STD_LOGIC;
  signal W_17_23_i_8_n_0 : STD_LOGIC;
  signal W_17_23_i_9_n_0 : STD_LOGIC;
  signal W_17_27_i_10_n_0 : STD_LOGIC;
  signal W_17_27_i_11_n_0 : STD_LOGIC;
  signal W_17_27_i_12_n_0 : STD_LOGIC;
  signal W_17_27_i_13_n_0 : STD_LOGIC;
  signal W_17_27_i_14_n_0 : STD_LOGIC;
  signal W_17_27_i_15_n_0 : STD_LOGIC;
  signal W_17_27_i_16_n_0 : STD_LOGIC;
  signal W_17_27_i_17_n_0 : STD_LOGIC;
  signal W_17_27_i_2_n_0 : STD_LOGIC;
  signal W_17_27_i_3_n_0 : STD_LOGIC;
  signal W_17_27_i_4_n_0 : STD_LOGIC;
  signal W_17_27_i_5_n_0 : STD_LOGIC;
  signal W_17_27_i_6_n_0 : STD_LOGIC;
  signal W_17_27_i_7_n_0 : STD_LOGIC;
  signal W_17_27_i_8_n_0 : STD_LOGIC;
  signal W_17_27_i_9_n_0 : STD_LOGIC;
  signal W_17_31_i_10_n_0 : STD_LOGIC;
  signal W_17_31_i_11_n_0 : STD_LOGIC;
  signal W_17_31_i_12_n_0 : STD_LOGIC;
  signal W_17_31_i_13_n_0 : STD_LOGIC;
  signal W_17_31_i_14_n_0 : STD_LOGIC;
  signal W_17_31_i_15_n_0 : STD_LOGIC;
  signal W_17_31_i_17_n_0 : STD_LOGIC;
  signal W_17_31_i_19_n_0 : STD_LOGIC;
  signal W_17_31_i_2_n_0 : STD_LOGIC;
  signal W_17_31_i_3_n_0 : STD_LOGIC;
  signal W_17_31_i_4_n_0 : STD_LOGIC;
  signal W_17_31_i_5_n_0 : STD_LOGIC;
  signal W_17_31_i_6_n_0 : STD_LOGIC;
  signal W_17_31_i_7_n_0 : STD_LOGIC;
  signal W_17_31_i_8_n_0 : STD_LOGIC;
  signal W_17_31_i_9_n_0 : STD_LOGIC;
  signal W_17_3_i_10_n_0 : STD_LOGIC;
  signal W_17_3_i_11_n_0 : STD_LOGIC;
  signal W_17_3_i_13_n_0 : STD_LOGIC;
  signal W_17_3_i_2_n_0 : STD_LOGIC;
  signal W_17_3_i_3_n_0 : STD_LOGIC;
  signal W_17_3_i_4_n_0 : STD_LOGIC;
  signal W_17_3_i_5_n_0 : STD_LOGIC;
  signal W_17_3_i_6_n_0 : STD_LOGIC;
  signal W_17_3_i_7_n_0 : STD_LOGIC;
  signal W_17_3_i_8_n_0 : STD_LOGIC;
  signal W_17_3_i_9_n_0 : STD_LOGIC;
  signal W_17_7_i_10_n_0 : STD_LOGIC;
  signal W_17_7_i_11_n_0 : STD_LOGIC;
  signal W_17_7_i_12_n_0 : STD_LOGIC;
  signal W_17_7_i_13_n_0 : STD_LOGIC;
  signal W_17_7_i_14_n_0 : STD_LOGIC;
  signal W_17_7_i_15_n_0 : STD_LOGIC;
  signal W_17_7_i_16_n_0 : STD_LOGIC;
  signal W_17_7_i_17_n_0 : STD_LOGIC;
  signal W_17_7_i_2_n_0 : STD_LOGIC;
  signal W_17_7_i_3_n_0 : STD_LOGIC;
  signal W_17_7_i_4_n_0 : STD_LOGIC;
  signal W_17_7_i_5_n_0 : STD_LOGIC;
  signal W_17_7_i_6_n_0 : STD_LOGIC;
  signal W_17_7_i_7_n_0 : STD_LOGIC;
  signal W_17_7_i_8_n_0 : STD_LOGIC;
  signal W_17_7_i_9_n_0 : STD_LOGIC;
  signal W_18_11_i_10_n_0 : STD_LOGIC;
  signal W_18_11_i_11_n_0 : STD_LOGIC;
  signal W_18_11_i_12_n_0 : STD_LOGIC;
  signal W_18_11_i_13_n_0 : STD_LOGIC;
  signal W_18_11_i_14_n_0 : STD_LOGIC;
  signal W_18_11_i_15_n_0 : STD_LOGIC;
  signal W_18_11_i_16_n_0 : STD_LOGIC;
  signal W_18_11_i_17_n_0 : STD_LOGIC;
  signal W_18_11_i_2_n_0 : STD_LOGIC;
  signal W_18_11_i_3_n_0 : STD_LOGIC;
  signal W_18_11_i_4_n_0 : STD_LOGIC;
  signal W_18_11_i_5_n_0 : STD_LOGIC;
  signal W_18_11_i_6_n_0 : STD_LOGIC;
  signal W_18_11_i_7_n_0 : STD_LOGIC;
  signal W_18_11_i_8_n_0 : STD_LOGIC;
  signal W_18_11_i_9_n_0 : STD_LOGIC;
  signal W_18_15_i_10_n_0 : STD_LOGIC;
  signal W_18_15_i_11_n_0 : STD_LOGIC;
  signal W_18_15_i_12_n_0 : STD_LOGIC;
  signal W_18_15_i_13_n_0 : STD_LOGIC;
  signal W_18_15_i_14_n_0 : STD_LOGIC;
  signal W_18_15_i_15_n_0 : STD_LOGIC;
  signal W_18_15_i_16_n_0 : STD_LOGIC;
  signal W_18_15_i_17_n_0 : STD_LOGIC;
  signal W_18_15_i_2_n_0 : STD_LOGIC;
  signal W_18_15_i_3_n_0 : STD_LOGIC;
  signal W_18_15_i_4_n_0 : STD_LOGIC;
  signal W_18_15_i_5_n_0 : STD_LOGIC;
  signal W_18_15_i_6_n_0 : STD_LOGIC;
  signal W_18_15_i_7_n_0 : STD_LOGIC;
  signal W_18_15_i_8_n_0 : STD_LOGIC;
  signal W_18_15_i_9_n_0 : STD_LOGIC;
  signal W_18_19_i_10_n_0 : STD_LOGIC;
  signal W_18_19_i_11_n_0 : STD_LOGIC;
  signal W_18_19_i_12_n_0 : STD_LOGIC;
  signal W_18_19_i_13_n_0 : STD_LOGIC;
  signal W_18_19_i_14_n_0 : STD_LOGIC;
  signal W_18_19_i_15_n_0 : STD_LOGIC;
  signal W_18_19_i_16_n_0 : STD_LOGIC;
  signal W_18_19_i_17_n_0 : STD_LOGIC;
  signal W_18_19_i_2_n_0 : STD_LOGIC;
  signal W_18_19_i_3_n_0 : STD_LOGIC;
  signal W_18_19_i_4_n_0 : STD_LOGIC;
  signal W_18_19_i_5_n_0 : STD_LOGIC;
  signal W_18_19_i_6_n_0 : STD_LOGIC;
  signal W_18_19_i_7_n_0 : STD_LOGIC;
  signal W_18_19_i_8_n_0 : STD_LOGIC;
  signal W_18_19_i_9_n_0 : STD_LOGIC;
  signal W_18_23_i_10_n_0 : STD_LOGIC;
  signal W_18_23_i_11_n_0 : STD_LOGIC;
  signal W_18_23_i_12_n_0 : STD_LOGIC;
  signal W_18_23_i_13_n_0 : STD_LOGIC;
  signal W_18_23_i_14_n_0 : STD_LOGIC;
  signal W_18_23_i_15_n_0 : STD_LOGIC;
  signal W_18_23_i_16_n_0 : STD_LOGIC;
  signal W_18_23_i_17_n_0 : STD_LOGIC;
  signal W_18_23_i_2_n_0 : STD_LOGIC;
  signal W_18_23_i_3_n_0 : STD_LOGIC;
  signal W_18_23_i_4_n_0 : STD_LOGIC;
  signal W_18_23_i_5_n_0 : STD_LOGIC;
  signal W_18_23_i_6_n_0 : STD_LOGIC;
  signal W_18_23_i_7_n_0 : STD_LOGIC;
  signal W_18_23_i_8_n_0 : STD_LOGIC;
  signal W_18_23_i_9_n_0 : STD_LOGIC;
  signal W_18_27_i_10_n_0 : STD_LOGIC;
  signal W_18_27_i_11_n_0 : STD_LOGIC;
  signal W_18_27_i_12_n_0 : STD_LOGIC;
  signal W_18_27_i_13_n_0 : STD_LOGIC;
  signal W_18_27_i_14_n_0 : STD_LOGIC;
  signal W_18_27_i_15_n_0 : STD_LOGIC;
  signal W_18_27_i_16_n_0 : STD_LOGIC;
  signal W_18_27_i_17_n_0 : STD_LOGIC;
  signal W_18_27_i_2_n_0 : STD_LOGIC;
  signal W_18_27_i_3_n_0 : STD_LOGIC;
  signal W_18_27_i_4_n_0 : STD_LOGIC;
  signal W_18_27_i_5_n_0 : STD_LOGIC;
  signal W_18_27_i_6_n_0 : STD_LOGIC;
  signal W_18_27_i_7_n_0 : STD_LOGIC;
  signal W_18_27_i_8_n_0 : STD_LOGIC;
  signal W_18_27_i_9_n_0 : STD_LOGIC;
  signal W_18_31_i_10_n_0 : STD_LOGIC;
  signal W_18_31_i_11_n_0 : STD_LOGIC;
  signal W_18_31_i_12_n_0 : STD_LOGIC;
  signal W_18_31_i_13_n_0 : STD_LOGIC;
  signal W_18_31_i_14_n_0 : STD_LOGIC;
  signal W_18_31_i_15_n_0 : STD_LOGIC;
  signal W_18_31_i_17_n_0 : STD_LOGIC;
  signal W_18_31_i_19_n_0 : STD_LOGIC;
  signal W_18_31_i_2_n_0 : STD_LOGIC;
  signal W_18_31_i_3_n_0 : STD_LOGIC;
  signal W_18_31_i_4_n_0 : STD_LOGIC;
  signal W_18_31_i_5_n_0 : STD_LOGIC;
  signal W_18_31_i_6_n_0 : STD_LOGIC;
  signal W_18_31_i_7_n_0 : STD_LOGIC;
  signal W_18_31_i_8_n_0 : STD_LOGIC;
  signal W_18_31_i_9_n_0 : STD_LOGIC;
  signal W_18_3_i_10_n_0 : STD_LOGIC;
  signal W_18_3_i_11_n_0 : STD_LOGIC;
  signal W_18_3_i_13_n_0 : STD_LOGIC;
  signal W_18_3_i_2_n_0 : STD_LOGIC;
  signal W_18_3_i_3_n_0 : STD_LOGIC;
  signal W_18_3_i_4_n_0 : STD_LOGIC;
  signal W_18_3_i_5_n_0 : STD_LOGIC;
  signal W_18_3_i_6_n_0 : STD_LOGIC;
  signal W_18_3_i_7_n_0 : STD_LOGIC;
  signal W_18_3_i_8_n_0 : STD_LOGIC;
  signal W_18_3_i_9_n_0 : STD_LOGIC;
  signal W_18_7_i_10_n_0 : STD_LOGIC;
  signal W_18_7_i_11_n_0 : STD_LOGIC;
  signal W_18_7_i_12_n_0 : STD_LOGIC;
  signal W_18_7_i_13_n_0 : STD_LOGIC;
  signal W_18_7_i_14_n_0 : STD_LOGIC;
  signal W_18_7_i_15_n_0 : STD_LOGIC;
  signal W_18_7_i_16_n_0 : STD_LOGIC;
  signal W_18_7_i_17_n_0 : STD_LOGIC;
  signal W_18_7_i_2_n_0 : STD_LOGIC;
  signal W_18_7_i_3_n_0 : STD_LOGIC;
  signal W_18_7_i_4_n_0 : STD_LOGIC;
  signal W_18_7_i_5_n_0 : STD_LOGIC;
  signal W_18_7_i_6_n_0 : STD_LOGIC;
  signal W_18_7_i_7_n_0 : STD_LOGIC;
  signal W_18_7_i_8_n_0 : STD_LOGIC;
  signal W_18_7_i_9_n_0 : STD_LOGIC;
  signal W_19_11_i_10_n_0 : STD_LOGIC;
  signal W_19_11_i_11_n_0 : STD_LOGIC;
  signal W_19_11_i_12_n_0 : STD_LOGIC;
  signal W_19_11_i_13_n_0 : STD_LOGIC;
  signal W_19_11_i_14_n_0 : STD_LOGIC;
  signal W_19_11_i_15_n_0 : STD_LOGIC;
  signal W_19_11_i_16_n_0 : STD_LOGIC;
  signal W_19_11_i_17_n_0 : STD_LOGIC;
  signal W_19_11_i_2_n_0 : STD_LOGIC;
  signal W_19_11_i_3_n_0 : STD_LOGIC;
  signal W_19_11_i_4_n_0 : STD_LOGIC;
  signal W_19_11_i_5_n_0 : STD_LOGIC;
  signal W_19_11_i_6_n_0 : STD_LOGIC;
  signal W_19_11_i_7_n_0 : STD_LOGIC;
  signal W_19_11_i_8_n_0 : STD_LOGIC;
  signal W_19_11_i_9_n_0 : STD_LOGIC;
  signal W_19_15_i_10_n_0 : STD_LOGIC;
  signal W_19_15_i_11_n_0 : STD_LOGIC;
  signal W_19_15_i_12_n_0 : STD_LOGIC;
  signal W_19_15_i_13_n_0 : STD_LOGIC;
  signal W_19_15_i_14_n_0 : STD_LOGIC;
  signal W_19_15_i_15_n_0 : STD_LOGIC;
  signal W_19_15_i_16_n_0 : STD_LOGIC;
  signal W_19_15_i_17_n_0 : STD_LOGIC;
  signal W_19_15_i_2_n_0 : STD_LOGIC;
  signal W_19_15_i_3_n_0 : STD_LOGIC;
  signal W_19_15_i_4_n_0 : STD_LOGIC;
  signal W_19_15_i_5_n_0 : STD_LOGIC;
  signal W_19_15_i_6_n_0 : STD_LOGIC;
  signal W_19_15_i_7_n_0 : STD_LOGIC;
  signal W_19_15_i_8_n_0 : STD_LOGIC;
  signal W_19_15_i_9_n_0 : STD_LOGIC;
  signal W_19_19_i_10_n_0 : STD_LOGIC;
  signal W_19_19_i_11_n_0 : STD_LOGIC;
  signal W_19_19_i_12_n_0 : STD_LOGIC;
  signal W_19_19_i_13_n_0 : STD_LOGIC;
  signal W_19_19_i_14_n_0 : STD_LOGIC;
  signal W_19_19_i_15_n_0 : STD_LOGIC;
  signal W_19_19_i_16_n_0 : STD_LOGIC;
  signal W_19_19_i_17_n_0 : STD_LOGIC;
  signal W_19_19_i_2_n_0 : STD_LOGIC;
  signal W_19_19_i_3_n_0 : STD_LOGIC;
  signal W_19_19_i_4_n_0 : STD_LOGIC;
  signal W_19_19_i_5_n_0 : STD_LOGIC;
  signal W_19_19_i_6_n_0 : STD_LOGIC;
  signal W_19_19_i_7_n_0 : STD_LOGIC;
  signal W_19_19_i_8_n_0 : STD_LOGIC;
  signal W_19_19_i_9_n_0 : STD_LOGIC;
  signal W_19_23_i_10_n_0 : STD_LOGIC;
  signal W_19_23_i_11_n_0 : STD_LOGIC;
  signal W_19_23_i_12_n_0 : STD_LOGIC;
  signal W_19_23_i_13_n_0 : STD_LOGIC;
  signal W_19_23_i_14_n_0 : STD_LOGIC;
  signal W_19_23_i_15_n_0 : STD_LOGIC;
  signal W_19_23_i_16_n_0 : STD_LOGIC;
  signal W_19_23_i_17_n_0 : STD_LOGIC;
  signal W_19_23_i_2_n_0 : STD_LOGIC;
  signal W_19_23_i_3_n_0 : STD_LOGIC;
  signal W_19_23_i_4_n_0 : STD_LOGIC;
  signal W_19_23_i_5_n_0 : STD_LOGIC;
  signal W_19_23_i_6_n_0 : STD_LOGIC;
  signal W_19_23_i_7_n_0 : STD_LOGIC;
  signal W_19_23_i_8_n_0 : STD_LOGIC;
  signal W_19_23_i_9_n_0 : STD_LOGIC;
  signal W_19_27_i_10_n_0 : STD_LOGIC;
  signal W_19_27_i_11_n_0 : STD_LOGIC;
  signal W_19_27_i_12_n_0 : STD_LOGIC;
  signal W_19_27_i_13_n_0 : STD_LOGIC;
  signal W_19_27_i_14_n_0 : STD_LOGIC;
  signal W_19_27_i_15_n_0 : STD_LOGIC;
  signal W_19_27_i_16_n_0 : STD_LOGIC;
  signal W_19_27_i_17_n_0 : STD_LOGIC;
  signal W_19_27_i_2_n_0 : STD_LOGIC;
  signal W_19_27_i_3_n_0 : STD_LOGIC;
  signal W_19_27_i_4_n_0 : STD_LOGIC;
  signal W_19_27_i_5_n_0 : STD_LOGIC;
  signal W_19_27_i_6_n_0 : STD_LOGIC;
  signal W_19_27_i_7_n_0 : STD_LOGIC;
  signal W_19_27_i_8_n_0 : STD_LOGIC;
  signal W_19_27_i_9_n_0 : STD_LOGIC;
  signal W_19_31_i_10_n_0 : STD_LOGIC;
  signal W_19_31_i_11_n_0 : STD_LOGIC;
  signal W_19_31_i_12_n_0 : STD_LOGIC;
  signal W_19_31_i_13_n_0 : STD_LOGIC;
  signal W_19_31_i_14_n_0 : STD_LOGIC;
  signal W_19_31_i_15_n_0 : STD_LOGIC;
  signal W_19_31_i_17_n_0 : STD_LOGIC;
  signal W_19_31_i_19_n_0 : STD_LOGIC;
  signal W_19_31_i_2_n_0 : STD_LOGIC;
  signal W_19_31_i_3_n_0 : STD_LOGIC;
  signal W_19_31_i_4_n_0 : STD_LOGIC;
  signal W_19_31_i_5_n_0 : STD_LOGIC;
  signal W_19_31_i_6_n_0 : STD_LOGIC;
  signal W_19_31_i_7_n_0 : STD_LOGIC;
  signal W_19_31_i_8_n_0 : STD_LOGIC;
  signal W_19_31_i_9_n_0 : STD_LOGIC;
  signal W_19_3_i_10_n_0 : STD_LOGIC;
  signal W_19_3_i_11_n_0 : STD_LOGIC;
  signal W_19_3_i_13_n_0 : STD_LOGIC;
  signal W_19_3_i_2_n_0 : STD_LOGIC;
  signal W_19_3_i_3_n_0 : STD_LOGIC;
  signal W_19_3_i_4_n_0 : STD_LOGIC;
  signal W_19_3_i_5_n_0 : STD_LOGIC;
  signal W_19_3_i_6_n_0 : STD_LOGIC;
  signal W_19_3_i_7_n_0 : STD_LOGIC;
  signal W_19_3_i_8_n_0 : STD_LOGIC;
  signal W_19_3_i_9_n_0 : STD_LOGIC;
  signal W_19_7_i_10_n_0 : STD_LOGIC;
  signal W_19_7_i_11_n_0 : STD_LOGIC;
  signal W_19_7_i_12_n_0 : STD_LOGIC;
  signal W_19_7_i_13_n_0 : STD_LOGIC;
  signal W_19_7_i_14_n_0 : STD_LOGIC;
  signal W_19_7_i_15_n_0 : STD_LOGIC;
  signal W_19_7_i_16_n_0 : STD_LOGIC;
  signal W_19_7_i_17_n_0 : STD_LOGIC;
  signal W_19_7_i_2_n_0 : STD_LOGIC;
  signal W_19_7_i_3_n_0 : STD_LOGIC;
  signal W_19_7_i_4_n_0 : STD_LOGIC;
  signal W_19_7_i_5_n_0 : STD_LOGIC;
  signal W_19_7_i_6_n_0 : STD_LOGIC;
  signal W_19_7_i_7_n_0 : STD_LOGIC;
  signal W_19_7_i_8_n_0 : STD_LOGIC;
  signal W_19_7_i_9_n_0 : STD_LOGIC;
  signal W_20_11_i_10_n_0 : STD_LOGIC;
  signal W_20_11_i_11_n_0 : STD_LOGIC;
  signal W_20_11_i_12_n_0 : STD_LOGIC;
  signal W_20_11_i_13_n_0 : STD_LOGIC;
  signal W_20_11_i_14_n_0 : STD_LOGIC;
  signal W_20_11_i_15_n_0 : STD_LOGIC;
  signal W_20_11_i_16_n_0 : STD_LOGIC;
  signal W_20_11_i_17_n_0 : STD_LOGIC;
  signal W_20_11_i_2_n_0 : STD_LOGIC;
  signal W_20_11_i_3_n_0 : STD_LOGIC;
  signal W_20_11_i_4_n_0 : STD_LOGIC;
  signal W_20_11_i_5_n_0 : STD_LOGIC;
  signal W_20_11_i_6_n_0 : STD_LOGIC;
  signal W_20_11_i_7_n_0 : STD_LOGIC;
  signal W_20_11_i_8_n_0 : STD_LOGIC;
  signal W_20_11_i_9_n_0 : STD_LOGIC;
  signal W_20_15_i_10_n_0 : STD_LOGIC;
  signal W_20_15_i_11_n_0 : STD_LOGIC;
  signal W_20_15_i_12_n_0 : STD_LOGIC;
  signal W_20_15_i_13_n_0 : STD_LOGIC;
  signal W_20_15_i_14_n_0 : STD_LOGIC;
  signal W_20_15_i_15_n_0 : STD_LOGIC;
  signal W_20_15_i_16_n_0 : STD_LOGIC;
  signal W_20_15_i_17_n_0 : STD_LOGIC;
  signal W_20_15_i_2_n_0 : STD_LOGIC;
  signal W_20_15_i_3_n_0 : STD_LOGIC;
  signal W_20_15_i_4_n_0 : STD_LOGIC;
  signal W_20_15_i_5_n_0 : STD_LOGIC;
  signal W_20_15_i_6_n_0 : STD_LOGIC;
  signal W_20_15_i_7_n_0 : STD_LOGIC;
  signal W_20_15_i_8_n_0 : STD_LOGIC;
  signal W_20_15_i_9_n_0 : STD_LOGIC;
  signal W_20_19_i_10_n_0 : STD_LOGIC;
  signal W_20_19_i_11_n_0 : STD_LOGIC;
  signal W_20_19_i_12_n_0 : STD_LOGIC;
  signal W_20_19_i_13_n_0 : STD_LOGIC;
  signal W_20_19_i_14_n_0 : STD_LOGIC;
  signal W_20_19_i_15_n_0 : STD_LOGIC;
  signal W_20_19_i_16_n_0 : STD_LOGIC;
  signal W_20_19_i_17_n_0 : STD_LOGIC;
  signal W_20_19_i_2_n_0 : STD_LOGIC;
  signal W_20_19_i_3_n_0 : STD_LOGIC;
  signal W_20_19_i_4_n_0 : STD_LOGIC;
  signal W_20_19_i_5_n_0 : STD_LOGIC;
  signal W_20_19_i_6_n_0 : STD_LOGIC;
  signal W_20_19_i_7_n_0 : STD_LOGIC;
  signal W_20_19_i_8_n_0 : STD_LOGIC;
  signal W_20_19_i_9_n_0 : STD_LOGIC;
  signal W_20_23_i_10_n_0 : STD_LOGIC;
  signal W_20_23_i_11_n_0 : STD_LOGIC;
  signal W_20_23_i_12_n_0 : STD_LOGIC;
  signal W_20_23_i_13_n_0 : STD_LOGIC;
  signal W_20_23_i_14_n_0 : STD_LOGIC;
  signal W_20_23_i_15_n_0 : STD_LOGIC;
  signal W_20_23_i_16_n_0 : STD_LOGIC;
  signal W_20_23_i_17_n_0 : STD_LOGIC;
  signal W_20_23_i_2_n_0 : STD_LOGIC;
  signal W_20_23_i_3_n_0 : STD_LOGIC;
  signal W_20_23_i_4_n_0 : STD_LOGIC;
  signal W_20_23_i_5_n_0 : STD_LOGIC;
  signal W_20_23_i_6_n_0 : STD_LOGIC;
  signal W_20_23_i_7_n_0 : STD_LOGIC;
  signal W_20_23_i_8_n_0 : STD_LOGIC;
  signal W_20_23_i_9_n_0 : STD_LOGIC;
  signal W_20_27_i_10_n_0 : STD_LOGIC;
  signal W_20_27_i_11_n_0 : STD_LOGIC;
  signal W_20_27_i_12_n_0 : STD_LOGIC;
  signal W_20_27_i_13_n_0 : STD_LOGIC;
  signal W_20_27_i_14_n_0 : STD_LOGIC;
  signal W_20_27_i_15_n_0 : STD_LOGIC;
  signal W_20_27_i_16_n_0 : STD_LOGIC;
  signal W_20_27_i_17_n_0 : STD_LOGIC;
  signal W_20_27_i_2_n_0 : STD_LOGIC;
  signal W_20_27_i_3_n_0 : STD_LOGIC;
  signal W_20_27_i_4_n_0 : STD_LOGIC;
  signal W_20_27_i_5_n_0 : STD_LOGIC;
  signal W_20_27_i_6_n_0 : STD_LOGIC;
  signal W_20_27_i_7_n_0 : STD_LOGIC;
  signal W_20_27_i_8_n_0 : STD_LOGIC;
  signal W_20_27_i_9_n_0 : STD_LOGIC;
  signal W_20_31_i_10_n_0 : STD_LOGIC;
  signal W_20_31_i_11_n_0 : STD_LOGIC;
  signal W_20_31_i_12_n_0 : STD_LOGIC;
  signal W_20_31_i_13_n_0 : STD_LOGIC;
  signal W_20_31_i_14_n_0 : STD_LOGIC;
  signal W_20_31_i_15_n_0 : STD_LOGIC;
  signal W_20_31_i_17_n_0 : STD_LOGIC;
  signal W_20_31_i_19_n_0 : STD_LOGIC;
  signal W_20_31_i_2_n_0 : STD_LOGIC;
  signal W_20_31_i_3_n_0 : STD_LOGIC;
  signal W_20_31_i_4_n_0 : STD_LOGIC;
  signal W_20_31_i_5_n_0 : STD_LOGIC;
  signal W_20_31_i_6_n_0 : STD_LOGIC;
  signal W_20_31_i_7_n_0 : STD_LOGIC;
  signal W_20_31_i_8_n_0 : STD_LOGIC;
  signal W_20_31_i_9_n_0 : STD_LOGIC;
  signal W_20_3_i_10_n_0 : STD_LOGIC;
  signal W_20_3_i_11_n_0 : STD_LOGIC;
  signal W_20_3_i_13_n_0 : STD_LOGIC;
  signal W_20_3_i_2_n_0 : STD_LOGIC;
  signal W_20_3_i_3_n_0 : STD_LOGIC;
  signal W_20_3_i_4_n_0 : STD_LOGIC;
  signal W_20_3_i_5_n_0 : STD_LOGIC;
  signal W_20_3_i_6_n_0 : STD_LOGIC;
  signal W_20_3_i_7_n_0 : STD_LOGIC;
  signal W_20_3_i_8_n_0 : STD_LOGIC;
  signal W_20_3_i_9_n_0 : STD_LOGIC;
  signal W_20_7_i_10_n_0 : STD_LOGIC;
  signal W_20_7_i_11_n_0 : STD_LOGIC;
  signal W_20_7_i_12_n_0 : STD_LOGIC;
  signal W_20_7_i_13_n_0 : STD_LOGIC;
  signal W_20_7_i_14_n_0 : STD_LOGIC;
  signal W_20_7_i_15_n_0 : STD_LOGIC;
  signal W_20_7_i_16_n_0 : STD_LOGIC;
  signal W_20_7_i_17_n_0 : STD_LOGIC;
  signal W_20_7_i_2_n_0 : STD_LOGIC;
  signal W_20_7_i_3_n_0 : STD_LOGIC;
  signal W_20_7_i_4_n_0 : STD_LOGIC;
  signal W_20_7_i_5_n_0 : STD_LOGIC;
  signal W_20_7_i_6_n_0 : STD_LOGIC;
  signal W_20_7_i_7_n_0 : STD_LOGIC;
  signal W_20_7_i_8_n_0 : STD_LOGIC;
  signal W_20_7_i_9_n_0 : STD_LOGIC;
  signal W_21_11_i_10_n_0 : STD_LOGIC;
  signal W_21_11_i_11_n_0 : STD_LOGIC;
  signal W_21_11_i_12_n_0 : STD_LOGIC;
  signal W_21_11_i_13_n_0 : STD_LOGIC;
  signal W_21_11_i_14_n_0 : STD_LOGIC;
  signal W_21_11_i_15_n_0 : STD_LOGIC;
  signal W_21_11_i_16_n_0 : STD_LOGIC;
  signal W_21_11_i_17_n_0 : STD_LOGIC;
  signal W_21_11_i_2_n_0 : STD_LOGIC;
  signal W_21_11_i_3_n_0 : STD_LOGIC;
  signal W_21_11_i_4_n_0 : STD_LOGIC;
  signal W_21_11_i_5_n_0 : STD_LOGIC;
  signal W_21_11_i_6_n_0 : STD_LOGIC;
  signal W_21_11_i_7_n_0 : STD_LOGIC;
  signal W_21_11_i_8_n_0 : STD_LOGIC;
  signal W_21_11_i_9_n_0 : STD_LOGIC;
  signal W_21_15_i_10_n_0 : STD_LOGIC;
  signal W_21_15_i_11_n_0 : STD_LOGIC;
  signal W_21_15_i_12_n_0 : STD_LOGIC;
  signal W_21_15_i_13_n_0 : STD_LOGIC;
  signal W_21_15_i_14_n_0 : STD_LOGIC;
  signal W_21_15_i_15_n_0 : STD_LOGIC;
  signal W_21_15_i_16_n_0 : STD_LOGIC;
  signal W_21_15_i_17_n_0 : STD_LOGIC;
  signal W_21_15_i_2_n_0 : STD_LOGIC;
  signal W_21_15_i_3_n_0 : STD_LOGIC;
  signal W_21_15_i_4_n_0 : STD_LOGIC;
  signal W_21_15_i_5_n_0 : STD_LOGIC;
  signal W_21_15_i_6_n_0 : STD_LOGIC;
  signal W_21_15_i_7_n_0 : STD_LOGIC;
  signal W_21_15_i_8_n_0 : STD_LOGIC;
  signal W_21_15_i_9_n_0 : STD_LOGIC;
  signal W_21_19_i_10_n_0 : STD_LOGIC;
  signal W_21_19_i_11_n_0 : STD_LOGIC;
  signal W_21_19_i_12_n_0 : STD_LOGIC;
  signal W_21_19_i_13_n_0 : STD_LOGIC;
  signal W_21_19_i_14_n_0 : STD_LOGIC;
  signal W_21_19_i_15_n_0 : STD_LOGIC;
  signal W_21_19_i_16_n_0 : STD_LOGIC;
  signal W_21_19_i_17_n_0 : STD_LOGIC;
  signal W_21_19_i_2_n_0 : STD_LOGIC;
  signal W_21_19_i_3_n_0 : STD_LOGIC;
  signal W_21_19_i_4_n_0 : STD_LOGIC;
  signal W_21_19_i_5_n_0 : STD_LOGIC;
  signal W_21_19_i_6_n_0 : STD_LOGIC;
  signal W_21_19_i_7_n_0 : STD_LOGIC;
  signal W_21_19_i_8_n_0 : STD_LOGIC;
  signal W_21_19_i_9_n_0 : STD_LOGIC;
  signal W_21_23_i_10_n_0 : STD_LOGIC;
  signal W_21_23_i_11_n_0 : STD_LOGIC;
  signal W_21_23_i_12_n_0 : STD_LOGIC;
  signal W_21_23_i_13_n_0 : STD_LOGIC;
  signal W_21_23_i_14_n_0 : STD_LOGIC;
  signal W_21_23_i_15_n_0 : STD_LOGIC;
  signal W_21_23_i_16_n_0 : STD_LOGIC;
  signal W_21_23_i_17_n_0 : STD_LOGIC;
  signal W_21_23_i_2_n_0 : STD_LOGIC;
  signal W_21_23_i_3_n_0 : STD_LOGIC;
  signal W_21_23_i_4_n_0 : STD_LOGIC;
  signal W_21_23_i_5_n_0 : STD_LOGIC;
  signal W_21_23_i_6_n_0 : STD_LOGIC;
  signal W_21_23_i_7_n_0 : STD_LOGIC;
  signal W_21_23_i_8_n_0 : STD_LOGIC;
  signal W_21_23_i_9_n_0 : STD_LOGIC;
  signal W_21_27_i_10_n_0 : STD_LOGIC;
  signal W_21_27_i_11_n_0 : STD_LOGIC;
  signal W_21_27_i_12_n_0 : STD_LOGIC;
  signal W_21_27_i_13_n_0 : STD_LOGIC;
  signal W_21_27_i_14_n_0 : STD_LOGIC;
  signal W_21_27_i_15_n_0 : STD_LOGIC;
  signal W_21_27_i_16_n_0 : STD_LOGIC;
  signal W_21_27_i_17_n_0 : STD_LOGIC;
  signal W_21_27_i_2_n_0 : STD_LOGIC;
  signal W_21_27_i_3_n_0 : STD_LOGIC;
  signal W_21_27_i_4_n_0 : STD_LOGIC;
  signal W_21_27_i_5_n_0 : STD_LOGIC;
  signal W_21_27_i_6_n_0 : STD_LOGIC;
  signal W_21_27_i_7_n_0 : STD_LOGIC;
  signal W_21_27_i_8_n_0 : STD_LOGIC;
  signal W_21_27_i_9_n_0 : STD_LOGIC;
  signal W_21_31_i_10_n_0 : STD_LOGIC;
  signal W_21_31_i_11_n_0 : STD_LOGIC;
  signal W_21_31_i_12_n_0 : STD_LOGIC;
  signal W_21_31_i_13_n_0 : STD_LOGIC;
  signal W_21_31_i_14_n_0 : STD_LOGIC;
  signal W_21_31_i_15_n_0 : STD_LOGIC;
  signal W_21_31_i_17_n_0 : STD_LOGIC;
  signal W_21_31_i_19_n_0 : STD_LOGIC;
  signal W_21_31_i_2_n_0 : STD_LOGIC;
  signal W_21_31_i_3_n_0 : STD_LOGIC;
  signal W_21_31_i_4_n_0 : STD_LOGIC;
  signal W_21_31_i_5_n_0 : STD_LOGIC;
  signal W_21_31_i_6_n_0 : STD_LOGIC;
  signal W_21_31_i_7_n_0 : STD_LOGIC;
  signal W_21_31_i_8_n_0 : STD_LOGIC;
  signal W_21_31_i_9_n_0 : STD_LOGIC;
  signal W_21_3_i_10_n_0 : STD_LOGIC;
  signal W_21_3_i_11_n_0 : STD_LOGIC;
  signal W_21_3_i_13_n_0 : STD_LOGIC;
  signal W_21_3_i_2_n_0 : STD_LOGIC;
  signal W_21_3_i_3_n_0 : STD_LOGIC;
  signal W_21_3_i_4_n_0 : STD_LOGIC;
  signal W_21_3_i_5_n_0 : STD_LOGIC;
  signal W_21_3_i_6_n_0 : STD_LOGIC;
  signal W_21_3_i_7_n_0 : STD_LOGIC;
  signal W_21_3_i_8_n_0 : STD_LOGIC;
  signal W_21_3_i_9_n_0 : STD_LOGIC;
  signal W_21_7_i_10_n_0 : STD_LOGIC;
  signal W_21_7_i_11_n_0 : STD_LOGIC;
  signal W_21_7_i_12_n_0 : STD_LOGIC;
  signal W_21_7_i_13_n_0 : STD_LOGIC;
  signal W_21_7_i_14_n_0 : STD_LOGIC;
  signal W_21_7_i_15_n_0 : STD_LOGIC;
  signal W_21_7_i_16_n_0 : STD_LOGIC;
  signal W_21_7_i_17_n_0 : STD_LOGIC;
  signal W_21_7_i_2_n_0 : STD_LOGIC;
  signal W_21_7_i_3_n_0 : STD_LOGIC;
  signal W_21_7_i_4_n_0 : STD_LOGIC;
  signal W_21_7_i_5_n_0 : STD_LOGIC;
  signal W_21_7_i_6_n_0 : STD_LOGIC;
  signal W_21_7_i_7_n_0 : STD_LOGIC;
  signal W_21_7_i_8_n_0 : STD_LOGIC;
  signal W_21_7_i_9_n_0 : STD_LOGIC;
  signal W_22_11_i_10_n_0 : STD_LOGIC;
  signal W_22_11_i_11_n_0 : STD_LOGIC;
  signal W_22_11_i_12_n_0 : STD_LOGIC;
  signal W_22_11_i_13_n_0 : STD_LOGIC;
  signal W_22_11_i_14_n_0 : STD_LOGIC;
  signal W_22_11_i_15_n_0 : STD_LOGIC;
  signal W_22_11_i_16_n_0 : STD_LOGIC;
  signal W_22_11_i_17_n_0 : STD_LOGIC;
  signal W_22_11_i_2_n_0 : STD_LOGIC;
  signal W_22_11_i_3_n_0 : STD_LOGIC;
  signal W_22_11_i_4_n_0 : STD_LOGIC;
  signal W_22_11_i_5_n_0 : STD_LOGIC;
  signal W_22_11_i_6_n_0 : STD_LOGIC;
  signal W_22_11_i_7_n_0 : STD_LOGIC;
  signal W_22_11_i_8_n_0 : STD_LOGIC;
  signal W_22_11_i_9_n_0 : STD_LOGIC;
  signal W_22_15_i_10_n_0 : STD_LOGIC;
  signal W_22_15_i_11_n_0 : STD_LOGIC;
  signal W_22_15_i_12_n_0 : STD_LOGIC;
  signal W_22_15_i_13_n_0 : STD_LOGIC;
  signal W_22_15_i_14_n_0 : STD_LOGIC;
  signal W_22_15_i_15_n_0 : STD_LOGIC;
  signal W_22_15_i_16_n_0 : STD_LOGIC;
  signal W_22_15_i_17_n_0 : STD_LOGIC;
  signal W_22_15_i_2_n_0 : STD_LOGIC;
  signal W_22_15_i_3_n_0 : STD_LOGIC;
  signal W_22_15_i_4_n_0 : STD_LOGIC;
  signal W_22_15_i_5_n_0 : STD_LOGIC;
  signal W_22_15_i_6_n_0 : STD_LOGIC;
  signal W_22_15_i_7_n_0 : STD_LOGIC;
  signal W_22_15_i_8_n_0 : STD_LOGIC;
  signal W_22_15_i_9_n_0 : STD_LOGIC;
  signal W_22_19_i_10_n_0 : STD_LOGIC;
  signal W_22_19_i_11_n_0 : STD_LOGIC;
  signal W_22_19_i_12_n_0 : STD_LOGIC;
  signal W_22_19_i_13_n_0 : STD_LOGIC;
  signal W_22_19_i_14_n_0 : STD_LOGIC;
  signal W_22_19_i_15_n_0 : STD_LOGIC;
  signal W_22_19_i_16_n_0 : STD_LOGIC;
  signal W_22_19_i_17_n_0 : STD_LOGIC;
  signal W_22_19_i_2_n_0 : STD_LOGIC;
  signal W_22_19_i_3_n_0 : STD_LOGIC;
  signal W_22_19_i_4_n_0 : STD_LOGIC;
  signal W_22_19_i_5_n_0 : STD_LOGIC;
  signal W_22_19_i_6_n_0 : STD_LOGIC;
  signal W_22_19_i_7_n_0 : STD_LOGIC;
  signal W_22_19_i_8_n_0 : STD_LOGIC;
  signal W_22_19_i_9_n_0 : STD_LOGIC;
  signal W_22_23_i_10_n_0 : STD_LOGIC;
  signal W_22_23_i_11_n_0 : STD_LOGIC;
  signal W_22_23_i_12_n_0 : STD_LOGIC;
  signal W_22_23_i_13_n_0 : STD_LOGIC;
  signal W_22_23_i_14_n_0 : STD_LOGIC;
  signal W_22_23_i_15_n_0 : STD_LOGIC;
  signal W_22_23_i_16_n_0 : STD_LOGIC;
  signal W_22_23_i_17_n_0 : STD_LOGIC;
  signal W_22_23_i_2_n_0 : STD_LOGIC;
  signal W_22_23_i_3_n_0 : STD_LOGIC;
  signal W_22_23_i_4_n_0 : STD_LOGIC;
  signal W_22_23_i_5_n_0 : STD_LOGIC;
  signal W_22_23_i_6_n_0 : STD_LOGIC;
  signal W_22_23_i_7_n_0 : STD_LOGIC;
  signal W_22_23_i_8_n_0 : STD_LOGIC;
  signal W_22_23_i_9_n_0 : STD_LOGIC;
  signal W_22_27_i_10_n_0 : STD_LOGIC;
  signal W_22_27_i_11_n_0 : STD_LOGIC;
  signal W_22_27_i_12_n_0 : STD_LOGIC;
  signal W_22_27_i_13_n_0 : STD_LOGIC;
  signal W_22_27_i_14_n_0 : STD_LOGIC;
  signal W_22_27_i_15_n_0 : STD_LOGIC;
  signal W_22_27_i_16_n_0 : STD_LOGIC;
  signal W_22_27_i_17_n_0 : STD_LOGIC;
  signal W_22_27_i_2_n_0 : STD_LOGIC;
  signal W_22_27_i_3_n_0 : STD_LOGIC;
  signal W_22_27_i_4_n_0 : STD_LOGIC;
  signal W_22_27_i_5_n_0 : STD_LOGIC;
  signal W_22_27_i_6_n_0 : STD_LOGIC;
  signal W_22_27_i_7_n_0 : STD_LOGIC;
  signal W_22_27_i_8_n_0 : STD_LOGIC;
  signal W_22_27_i_9_n_0 : STD_LOGIC;
  signal W_22_31_i_10_n_0 : STD_LOGIC;
  signal W_22_31_i_11_n_0 : STD_LOGIC;
  signal W_22_31_i_12_n_0 : STD_LOGIC;
  signal W_22_31_i_13_n_0 : STD_LOGIC;
  signal W_22_31_i_14_n_0 : STD_LOGIC;
  signal W_22_31_i_15_n_0 : STD_LOGIC;
  signal W_22_31_i_17_n_0 : STD_LOGIC;
  signal W_22_31_i_19_n_0 : STD_LOGIC;
  signal W_22_31_i_2_n_0 : STD_LOGIC;
  signal W_22_31_i_3_n_0 : STD_LOGIC;
  signal W_22_31_i_4_n_0 : STD_LOGIC;
  signal W_22_31_i_5_n_0 : STD_LOGIC;
  signal W_22_31_i_6_n_0 : STD_LOGIC;
  signal W_22_31_i_7_n_0 : STD_LOGIC;
  signal W_22_31_i_8_n_0 : STD_LOGIC;
  signal W_22_31_i_9_n_0 : STD_LOGIC;
  signal W_22_3_i_10_n_0 : STD_LOGIC;
  signal W_22_3_i_11_n_0 : STD_LOGIC;
  signal W_22_3_i_13_n_0 : STD_LOGIC;
  signal W_22_3_i_2_n_0 : STD_LOGIC;
  signal W_22_3_i_3_n_0 : STD_LOGIC;
  signal W_22_3_i_4_n_0 : STD_LOGIC;
  signal W_22_3_i_5_n_0 : STD_LOGIC;
  signal W_22_3_i_6_n_0 : STD_LOGIC;
  signal W_22_3_i_7_n_0 : STD_LOGIC;
  signal W_22_3_i_8_n_0 : STD_LOGIC;
  signal W_22_3_i_9_n_0 : STD_LOGIC;
  signal W_22_7_i_10_n_0 : STD_LOGIC;
  signal W_22_7_i_11_n_0 : STD_LOGIC;
  signal W_22_7_i_12_n_0 : STD_LOGIC;
  signal W_22_7_i_13_n_0 : STD_LOGIC;
  signal W_22_7_i_14_n_0 : STD_LOGIC;
  signal W_22_7_i_15_n_0 : STD_LOGIC;
  signal W_22_7_i_16_n_0 : STD_LOGIC;
  signal W_22_7_i_17_n_0 : STD_LOGIC;
  signal W_22_7_i_2_n_0 : STD_LOGIC;
  signal W_22_7_i_3_n_0 : STD_LOGIC;
  signal W_22_7_i_4_n_0 : STD_LOGIC;
  signal W_22_7_i_5_n_0 : STD_LOGIC;
  signal W_22_7_i_6_n_0 : STD_LOGIC;
  signal W_22_7_i_7_n_0 : STD_LOGIC;
  signal W_22_7_i_8_n_0 : STD_LOGIC;
  signal W_22_7_i_9_n_0 : STD_LOGIC;
  signal W_23_11_i_10_n_0 : STD_LOGIC;
  signal W_23_11_i_11_n_0 : STD_LOGIC;
  signal W_23_11_i_12_n_0 : STD_LOGIC;
  signal W_23_11_i_13_n_0 : STD_LOGIC;
  signal W_23_11_i_14_n_0 : STD_LOGIC;
  signal W_23_11_i_15_n_0 : STD_LOGIC;
  signal W_23_11_i_16_n_0 : STD_LOGIC;
  signal W_23_11_i_17_n_0 : STD_LOGIC;
  signal W_23_11_i_2_n_0 : STD_LOGIC;
  signal W_23_11_i_3_n_0 : STD_LOGIC;
  signal W_23_11_i_4_n_0 : STD_LOGIC;
  signal W_23_11_i_5_n_0 : STD_LOGIC;
  signal W_23_11_i_6_n_0 : STD_LOGIC;
  signal W_23_11_i_7_n_0 : STD_LOGIC;
  signal W_23_11_i_8_n_0 : STD_LOGIC;
  signal W_23_11_i_9_n_0 : STD_LOGIC;
  signal W_23_15_i_10_n_0 : STD_LOGIC;
  signal W_23_15_i_11_n_0 : STD_LOGIC;
  signal W_23_15_i_12_n_0 : STD_LOGIC;
  signal W_23_15_i_13_n_0 : STD_LOGIC;
  signal W_23_15_i_14_n_0 : STD_LOGIC;
  signal W_23_15_i_15_n_0 : STD_LOGIC;
  signal W_23_15_i_16_n_0 : STD_LOGIC;
  signal W_23_15_i_17_n_0 : STD_LOGIC;
  signal W_23_15_i_2_n_0 : STD_LOGIC;
  signal W_23_15_i_3_n_0 : STD_LOGIC;
  signal W_23_15_i_4_n_0 : STD_LOGIC;
  signal W_23_15_i_5_n_0 : STD_LOGIC;
  signal W_23_15_i_6_n_0 : STD_LOGIC;
  signal W_23_15_i_7_n_0 : STD_LOGIC;
  signal W_23_15_i_8_n_0 : STD_LOGIC;
  signal W_23_15_i_9_n_0 : STD_LOGIC;
  signal W_23_19_i_10_n_0 : STD_LOGIC;
  signal W_23_19_i_11_n_0 : STD_LOGIC;
  signal W_23_19_i_12_n_0 : STD_LOGIC;
  signal W_23_19_i_13_n_0 : STD_LOGIC;
  signal W_23_19_i_14_n_0 : STD_LOGIC;
  signal W_23_19_i_15_n_0 : STD_LOGIC;
  signal W_23_19_i_16_n_0 : STD_LOGIC;
  signal W_23_19_i_17_n_0 : STD_LOGIC;
  signal W_23_19_i_2_n_0 : STD_LOGIC;
  signal W_23_19_i_3_n_0 : STD_LOGIC;
  signal W_23_19_i_4_n_0 : STD_LOGIC;
  signal W_23_19_i_5_n_0 : STD_LOGIC;
  signal W_23_19_i_6_n_0 : STD_LOGIC;
  signal W_23_19_i_7_n_0 : STD_LOGIC;
  signal W_23_19_i_8_n_0 : STD_LOGIC;
  signal W_23_19_i_9_n_0 : STD_LOGIC;
  signal W_23_23_i_10_n_0 : STD_LOGIC;
  signal W_23_23_i_11_n_0 : STD_LOGIC;
  signal W_23_23_i_12_n_0 : STD_LOGIC;
  signal W_23_23_i_13_n_0 : STD_LOGIC;
  signal W_23_23_i_14_n_0 : STD_LOGIC;
  signal W_23_23_i_15_n_0 : STD_LOGIC;
  signal W_23_23_i_16_n_0 : STD_LOGIC;
  signal W_23_23_i_17_n_0 : STD_LOGIC;
  signal W_23_23_i_2_n_0 : STD_LOGIC;
  signal W_23_23_i_3_n_0 : STD_LOGIC;
  signal W_23_23_i_4_n_0 : STD_LOGIC;
  signal W_23_23_i_5_n_0 : STD_LOGIC;
  signal W_23_23_i_6_n_0 : STD_LOGIC;
  signal W_23_23_i_7_n_0 : STD_LOGIC;
  signal W_23_23_i_8_n_0 : STD_LOGIC;
  signal W_23_23_i_9_n_0 : STD_LOGIC;
  signal W_23_27_i_10_n_0 : STD_LOGIC;
  signal W_23_27_i_11_n_0 : STD_LOGIC;
  signal W_23_27_i_12_n_0 : STD_LOGIC;
  signal W_23_27_i_13_n_0 : STD_LOGIC;
  signal W_23_27_i_14_n_0 : STD_LOGIC;
  signal W_23_27_i_15_n_0 : STD_LOGIC;
  signal W_23_27_i_16_n_0 : STD_LOGIC;
  signal W_23_27_i_17_n_0 : STD_LOGIC;
  signal W_23_27_i_2_n_0 : STD_LOGIC;
  signal W_23_27_i_3_n_0 : STD_LOGIC;
  signal W_23_27_i_4_n_0 : STD_LOGIC;
  signal W_23_27_i_5_n_0 : STD_LOGIC;
  signal W_23_27_i_6_n_0 : STD_LOGIC;
  signal W_23_27_i_7_n_0 : STD_LOGIC;
  signal W_23_27_i_8_n_0 : STD_LOGIC;
  signal W_23_27_i_9_n_0 : STD_LOGIC;
  signal W_23_31_i_10_n_0 : STD_LOGIC;
  signal W_23_31_i_11_n_0 : STD_LOGIC;
  signal W_23_31_i_12_n_0 : STD_LOGIC;
  signal W_23_31_i_13_n_0 : STD_LOGIC;
  signal W_23_31_i_14_n_0 : STD_LOGIC;
  signal W_23_31_i_15_n_0 : STD_LOGIC;
  signal W_23_31_i_17_n_0 : STD_LOGIC;
  signal W_23_31_i_19_n_0 : STD_LOGIC;
  signal W_23_31_i_2_n_0 : STD_LOGIC;
  signal W_23_31_i_3_n_0 : STD_LOGIC;
  signal W_23_31_i_4_n_0 : STD_LOGIC;
  signal W_23_31_i_5_n_0 : STD_LOGIC;
  signal W_23_31_i_6_n_0 : STD_LOGIC;
  signal W_23_31_i_7_n_0 : STD_LOGIC;
  signal W_23_31_i_8_n_0 : STD_LOGIC;
  signal W_23_31_i_9_n_0 : STD_LOGIC;
  signal W_23_3_i_10_n_0 : STD_LOGIC;
  signal W_23_3_i_11_n_0 : STD_LOGIC;
  signal W_23_3_i_2_n_0 : STD_LOGIC;
  signal W_23_3_i_3_n_0 : STD_LOGIC;
  signal W_23_3_i_4_n_0 : STD_LOGIC;
  signal W_23_3_i_5_n_0 : STD_LOGIC;
  signal W_23_3_i_6_n_0 : STD_LOGIC;
  signal W_23_3_i_7_n_0 : STD_LOGIC;
  signal W_23_3_i_8_n_0 : STD_LOGIC;
  signal W_23_3_i_9_n_0 : STD_LOGIC;
  signal W_23_7_i_10_n_0 : STD_LOGIC;
  signal W_23_7_i_11_n_0 : STD_LOGIC;
  signal W_23_7_i_12_n_0 : STD_LOGIC;
  signal W_23_7_i_13_n_0 : STD_LOGIC;
  signal W_23_7_i_14_n_0 : STD_LOGIC;
  signal W_23_7_i_15_n_0 : STD_LOGIC;
  signal W_23_7_i_16_n_0 : STD_LOGIC;
  signal W_23_7_i_17_n_0 : STD_LOGIC;
  signal W_23_7_i_2_n_0 : STD_LOGIC;
  signal W_23_7_i_3_n_0 : STD_LOGIC;
  signal W_23_7_i_4_n_0 : STD_LOGIC;
  signal W_23_7_i_5_n_0 : STD_LOGIC;
  signal W_23_7_i_6_n_0 : STD_LOGIC;
  signal W_23_7_i_7_n_0 : STD_LOGIC;
  signal W_23_7_i_8_n_0 : STD_LOGIC;
  signal W_23_7_i_9_n_0 : STD_LOGIC;
  signal W_24_11_i_10_n_0 : STD_LOGIC;
  signal W_24_11_i_11_n_0 : STD_LOGIC;
  signal W_24_11_i_12_n_0 : STD_LOGIC;
  signal W_24_11_i_13_n_0 : STD_LOGIC;
  signal W_24_11_i_14_n_0 : STD_LOGIC;
  signal W_24_11_i_15_n_0 : STD_LOGIC;
  signal W_24_11_i_16_n_0 : STD_LOGIC;
  signal W_24_11_i_17_n_0 : STD_LOGIC;
  signal W_24_11_i_2_n_0 : STD_LOGIC;
  signal W_24_11_i_3_n_0 : STD_LOGIC;
  signal W_24_11_i_4_n_0 : STD_LOGIC;
  signal W_24_11_i_5_n_0 : STD_LOGIC;
  signal W_24_11_i_6_n_0 : STD_LOGIC;
  signal W_24_11_i_7_n_0 : STD_LOGIC;
  signal W_24_11_i_8_n_0 : STD_LOGIC;
  signal W_24_11_i_9_n_0 : STD_LOGIC;
  signal W_24_15_i_10_n_0 : STD_LOGIC;
  signal W_24_15_i_11_n_0 : STD_LOGIC;
  signal W_24_15_i_12_n_0 : STD_LOGIC;
  signal W_24_15_i_13_n_0 : STD_LOGIC;
  signal W_24_15_i_14_n_0 : STD_LOGIC;
  signal W_24_15_i_15_n_0 : STD_LOGIC;
  signal W_24_15_i_16_n_0 : STD_LOGIC;
  signal W_24_15_i_17_n_0 : STD_LOGIC;
  signal W_24_15_i_2_n_0 : STD_LOGIC;
  signal W_24_15_i_3_n_0 : STD_LOGIC;
  signal W_24_15_i_4_n_0 : STD_LOGIC;
  signal W_24_15_i_5_n_0 : STD_LOGIC;
  signal W_24_15_i_6_n_0 : STD_LOGIC;
  signal W_24_15_i_7_n_0 : STD_LOGIC;
  signal W_24_15_i_8_n_0 : STD_LOGIC;
  signal W_24_15_i_9_n_0 : STD_LOGIC;
  signal W_24_19_i_10_n_0 : STD_LOGIC;
  signal W_24_19_i_11_n_0 : STD_LOGIC;
  signal W_24_19_i_12_n_0 : STD_LOGIC;
  signal W_24_19_i_13_n_0 : STD_LOGIC;
  signal W_24_19_i_14_n_0 : STD_LOGIC;
  signal W_24_19_i_15_n_0 : STD_LOGIC;
  signal W_24_19_i_16_n_0 : STD_LOGIC;
  signal W_24_19_i_17_n_0 : STD_LOGIC;
  signal W_24_19_i_2_n_0 : STD_LOGIC;
  signal W_24_19_i_3_n_0 : STD_LOGIC;
  signal W_24_19_i_4_n_0 : STD_LOGIC;
  signal W_24_19_i_5_n_0 : STD_LOGIC;
  signal W_24_19_i_6_n_0 : STD_LOGIC;
  signal W_24_19_i_7_n_0 : STD_LOGIC;
  signal W_24_19_i_8_n_0 : STD_LOGIC;
  signal W_24_19_i_9_n_0 : STD_LOGIC;
  signal W_24_23_i_10_n_0 : STD_LOGIC;
  signal W_24_23_i_11_n_0 : STD_LOGIC;
  signal W_24_23_i_12_n_0 : STD_LOGIC;
  signal W_24_23_i_13_n_0 : STD_LOGIC;
  signal W_24_23_i_14_n_0 : STD_LOGIC;
  signal W_24_23_i_15_n_0 : STD_LOGIC;
  signal W_24_23_i_16_n_0 : STD_LOGIC;
  signal W_24_23_i_17_n_0 : STD_LOGIC;
  signal W_24_23_i_2_n_0 : STD_LOGIC;
  signal W_24_23_i_3_n_0 : STD_LOGIC;
  signal W_24_23_i_4_n_0 : STD_LOGIC;
  signal W_24_23_i_5_n_0 : STD_LOGIC;
  signal W_24_23_i_6_n_0 : STD_LOGIC;
  signal W_24_23_i_7_n_0 : STD_LOGIC;
  signal W_24_23_i_8_n_0 : STD_LOGIC;
  signal W_24_23_i_9_n_0 : STD_LOGIC;
  signal W_24_27_i_10_n_0 : STD_LOGIC;
  signal W_24_27_i_11_n_0 : STD_LOGIC;
  signal W_24_27_i_12_n_0 : STD_LOGIC;
  signal W_24_27_i_13_n_0 : STD_LOGIC;
  signal W_24_27_i_14_n_0 : STD_LOGIC;
  signal W_24_27_i_15_n_0 : STD_LOGIC;
  signal W_24_27_i_16_n_0 : STD_LOGIC;
  signal W_24_27_i_17_n_0 : STD_LOGIC;
  signal W_24_27_i_2_n_0 : STD_LOGIC;
  signal W_24_27_i_3_n_0 : STD_LOGIC;
  signal W_24_27_i_4_n_0 : STD_LOGIC;
  signal W_24_27_i_5_n_0 : STD_LOGIC;
  signal W_24_27_i_6_n_0 : STD_LOGIC;
  signal W_24_27_i_7_n_0 : STD_LOGIC;
  signal W_24_27_i_8_n_0 : STD_LOGIC;
  signal W_24_27_i_9_n_0 : STD_LOGIC;
  signal W_24_31_i_10_n_0 : STD_LOGIC;
  signal W_24_31_i_11_n_0 : STD_LOGIC;
  signal W_24_31_i_12_n_0 : STD_LOGIC;
  signal W_24_31_i_13_n_0 : STD_LOGIC;
  signal W_24_31_i_14_n_0 : STD_LOGIC;
  signal W_24_31_i_15_n_0 : STD_LOGIC;
  signal W_24_31_i_17_n_0 : STD_LOGIC;
  signal W_24_31_i_19_n_0 : STD_LOGIC;
  signal W_24_31_i_2_n_0 : STD_LOGIC;
  signal W_24_31_i_3_n_0 : STD_LOGIC;
  signal W_24_31_i_4_n_0 : STD_LOGIC;
  signal W_24_31_i_5_n_0 : STD_LOGIC;
  signal W_24_31_i_6_n_0 : STD_LOGIC;
  signal W_24_31_i_7_n_0 : STD_LOGIC;
  signal W_24_31_i_8_n_0 : STD_LOGIC;
  signal W_24_31_i_9_n_0 : STD_LOGIC;
  signal W_24_3_i_10_n_0 : STD_LOGIC;
  signal W_24_3_i_11_n_0 : STD_LOGIC;
  signal W_24_3_i_2_n_0 : STD_LOGIC;
  signal W_24_3_i_3_n_0 : STD_LOGIC;
  signal W_24_3_i_4_n_0 : STD_LOGIC;
  signal W_24_3_i_5_n_0 : STD_LOGIC;
  signal W_24_3_i_6_n_0 : STD_LOGIC;
  signal W_24_3_i_7_n_0 : STD_LOGIC;
  signal W_24_3_i_8_n_0 : STD_LOGIC;
  signal W_24_3_i_9_n_0 : STD_LOGIC;
  signal W_24_7_i_10_n_0 : STD_LOGIC;
  signal W_24_7_i_11_n_0 : STD_LOGIC;
  signal W_24_7_i_12_n_0 : STD_LOGIC;
  signal W_24_7_i_13_n_0 : STD_LOGIC;
  signal W_24_7_i_14_n_0 : STD_LOGIC;
  signal W_24_7_i_15_n_0 : STD_LOGIC;
  signal W_24_7_i_16_n_0 : STD_LOGIC;
  signal W_24_7_i_17_n_0 : STD_LOGIC;
  signal W_24_7_i_2_n_0 : STD_LOGIC;
  signal W_24_7_i_3_n_0 : STD_LOGIC;
  signal W_24_7_i_4_n_0 : STD_LOGIC;
  signal W_24_7_i_5_n_0 : STD_LOGIC;
  signal W_24_7_i_6_n_0 : STD_LOGIC;
  signal W_24_7_i_7_n_0 : STD_LOGIC;
  signal W_24_7_i_8_n_0 : STD_LOGIC;
  signal W_24_7_i_9_n_0 : STD_LOGIC;
  signal W_25_11_i_10_n_0 : STD_LOGIC;
  signal W_25_11_i_11_n_0 : STD_LOGIC;
  signal W_25_11_i_12_n_0 : STD_LOGIC;
  signal W_25_11_i_13_n_0 : STD_LOGIC;
  signal W_25_11_i_14_n_0 : STD_LOGIC;
  signal W_25_11_i_15_n_0 : STD_LOGIC;
  signal W_25_11_i_16_n_0 : STD_LOGIC;
  signal W_25_11_i_17_n_0 : STD_LOGIC;
  signal W_25_11_i_2_n_0 : STD_LOGIC;
  signal W_25_11_i_3_n_0 : STD_LOGIC;
  signal W_25_11_i_4_n_0 : STD_LOGIC;
  signal W_25_11_i_5_n_0 : STD_LOGIC;
  signal W_25_11_i_6_n_0 : STD_LOGIC;
  signal W_25_11_i_7_n_0 : STD_LOGIC;
  signal W_25_11_i_8_n_0 : STD_LOGIC;
  signal W_25_11_i_9_n_0 : STD_LOGIC;
  signal W_25_15_i_10_n_0 : STD_LOGIC;
  signal W_25_15_i_11_n_0 : STD_LOGIC;
  signal W_25_15_i_12_n_0 : STD_LOGIC;
  signal W_25_15_i_13_n_0 : STD_LOGIC;
  signal W_25_15_i_14_n_0 : STD_LOGIC;
  signal W_25_15_i_15_n_0 : STD_LOGIC;
  signal W_25_15_i_16_n_0 : STD_LOGIC;
  signal W_25_15_i_17_n_0 : STD_LOGIC;
  signal W_25_15_i_2_n_0 : STD_LOGIC;
  signal W_25_15_i_3_n_0 : STD_LOGIC;
  signal W_25_15_i_4_n_0 : STD_LOGIC;
  signal W_25_15_i_5_n_0 : STD_LOGIC;
  signal W_25_15_i_6_n_0 : STD_LOGIC;
  signal W_25_15_i_7_n_0 : STD_LOGIC;
  signal W_25_15_i_8_n_0 : STD_LOGIC;
  signal W_25_15_i_9_n_0 : STD_LOGIC;
  signal W_25_19_i_10_n_0 : STD_LOGIC;
  signal W_25_19_i_11_n_0 : STD_LOGIC;
  signal W_25_19_i_12_n_0 : STD_LOGIC;
  signal W_25_19_i_13_n_0 : STD_LOGIC;
  signal W_25_19_i_14_n_0 : STD_LOGIC;
  signal W_25_19_i_15_n_0 : STD_LOGIC;
  signal W_25_19_i_16_n_0 : STD_LOGIC;
  signal W_25_19_i_17_n_0 : STD_LOGIC;
  signal W_25_19_i_2_n_0 : STD_LOGIC;
  signal W_25_19_i_3_n_0 : STD_LOGIC;
  signal W_25_19_i_4_n_0 : STD_LOGIC;
  signal W_25_19_i_5_n_0 : STD_LOGIC;
  signal W_25_19_i_6_n_0 : STD_LOGIC;
  signal W_25_19_i_7_n_0 : STD_LOGIC;
  signal W_25_19_i_8_n_0 : STD_LOGIC;
  signal W_25_19_i_9_n_0 : STD_LOGIC;
  signal W_25_23_i_10_n_0 : STD_LOGIC;
  signal W_25_23_i_11_n_0 : STD_LOGIC;
  signal W_25_23_i_12_n_0 : STD_LOGIC;
  signal W_25_23_i_13_n_0 : STD_LOGIC;
  signal W_25_23_i_14_n_0 : STD_LOGIC;
  signal W_25_23_i_15_n_0 : STD_LOGIC;
  signal W_25_23_i_16_n_0 : STD_LOGIC;
  signal W_25_23_i_17_n_0 : STD_LOGIC;
  signal W_25_23_i_2_n_0 : STD_LOGIC;
  signal W_25_23_i_3_n_0 : STD_LOGIC;
  signal W_25_23_i_4_n_0 : STD_LOGIC;
  signal W_25_23_i_5_n_0 : STD_LOGIC;
  signal W_25_23_i_6_n_0 : STD_LOGIC;
  signal W_25_23_i_7_n_0 : STD_LOGIC;
  signal W_25_23_i_8_n_0 : STD_LOGIC;
  signal W_25_23_i_9_n_0 : STD_LOGIC;
  signal W_25_27_i_10_n_0 : STD_LOGIC;
  signal W_25_27_i_11_n_0 : STD_LOGIC;
  signal W_25_27_i_12_n_0 : STD_LOGIC;
  signal W_25_27_i_13_n_0 : STD_LOGIC;
  signal W_25_27_i_14_n_0 : STD_LOGIC;
  signal W_25_27_i_15_n_0 : STD_LOGIC;
  signal W_25_27_i_16_n_0 : STD_LOGIC;
  signal W_25_27_i_17_n_0 : STD_LOGIC;
  signal W_25_27_i_2_n_0 : STD_LOGIC;
  signal W_25_27_i_3_n_0 : STD_LOGIC;
  signal W_25_27_i_4_n_0 : STD_LOGIC;
  signal W_25_27_i_5_n_0 : STD_LOGIC;
  signal W_25_27_i_6_n_0 : STD_LOGIC;
  signal W_25_27_i_7_n_0 : STD_LOGIC;
  signal W_25_27_i_8_n_0 : STD_LOGIC;
  signal W_25_27_i_9_n_0 : STD_LOGIC;
  signal W_25_31_i_10_n_0 : STD_LOGIC;
  signal W_25_31_i_11_n_0 : STD_LOGIC;
  signal W_25_31_i_12_n_0 : STD_LOGIC;
  signal W_25_31_i_13_n_0 : STD_LOGIC;
  signal W_25_31_i_14_n_0 : STD_LOGIC;
  signal W_25_31_i_15_n_0 : STD_LOGIC;
  signal W_25_31_i_17_n_0 : STD_LOGIC;
  signal W_25_31_i_19_n_0 : STD_LOGIC;
  signal W_25_31_i_2_n_0 : STD_LOGIC;
  signal W_25_31_i_3_n_0 : STD_LOGIC;
  signal W_25_31_i_4_n_0 : STD_LOGIC;
  signal W_25_31_i_5_n_0 : STD_LOGIC;
  signal W_25_31_i_6_n_0 : STD_LOGIC;
  signal W_25_31_i_7_n_0 : STD_LOGIC;
  signal W_25_31_i_8_n_0 : STD_LOGIC;
  signal W_25_31_i_9_n_0 : STD_LOGIC;
  signal W_25_3_i_10_n_0 : STD_LOGIC;
  signal W_25_3_i_11_n_0 : STD_LOGIC;
  signal W_25_3_i_2_n_0 : STD_LOGIC;
  signal W_25_3_i_3_n_0 : STD_LOGIC;
  signal W_25_3_i_4_n_0 : STD_LOGIC;
  signal W_25_3_i_5_n_0 : STD_LOGIC;
  signal W_25_3_i_6_n_0 : STD_LOGIC;
  signal W_25_3_i_7_n_0 : STD_LOGIC;
  signal W_25_3_i_8_n_0 : STD_LOGIC;
  signal W_25_3_i_9_n_0 : STD_LOGIC;
  signal W_25_7_i_10_n_0 : STD_LOGIC;
  signal W_25_7_i_11_n_0 : STD_LOGIC;
  signal W_25_7_i_12_n_0 : STD_LOGIC;
  signal W_25_7_i_13_n_0 : STD_LOGIC;
  signal W_25_7_i_14_n_0 : STD_LOGIC;
  signal W_25_7_i_15_n_0 : STD_LOGIC;
  signal W_25_7_i_16_n_0 : STD_LOGIC;
  signal W_25_7_i_17_n_0 : STD_LOGIC;
  signal W_25_7_i_2_n_0 : STD_LOGIC;
  signal W_25_7_i_3_n_0 : STD_LOGIC;
  signal W_25_7_i_4_n_0 : STD_LOGIC;
  signal W_25_7_i_5_n_0 : STD_LOGIC;
  signal W_25_7_i_6_n_0 : STD_LOGIC;
  signal W_25_7_i_7_n_0 : STD_LOGIC;
  signal W_25_7_i_8_n_0 : STD_LOGIC;
  signal W_25_7_i_9_n_0 : STD_LOGIC;
  signal W_26_11_i_10_n_0 : STD_LOGIC;
  signal W_26_11_i_11_n_0 : STD_LOGIC;
  signal W_26_11_i_12_n_0 : STD_LOGIC;
  signal W_26_11_i_13_n_0 : STD_LOGIC;
  signal W_26_11_i_14_n_0 : STD_LOGIC;
  signal W_26_11_i_15_n_0 : STD_LOGIC;
  signal W_26_11_i_16_n_0 : STD_LOGIC;
  signal W_26_11_i_17_n_0 : STD_LOGIC;
  signal W_26_11_i_2_n_0 : STD_LOGIC;
  signal W_26_11_i_3_n_0 : STD_LOGIC;
  signal W_26_11_i_4_n_0 : STD_LOGIC;
  signal W_26_11_i_5_n_0 : STD_LOGIC;
  signal W_26_11_i_6_n_0 : STD_LOGIC;
  signal W_26_11_i_7_n_0 : STD_LOGIC;
  signal W_26_11_i_8_n_0 : STD_LOGIC;
  signal W_26_11_i_9_n_0 : STD_LOGIC;
  signal W_26_15_i_10_n_0 : STD_LOGIC;
  signal W_26_15_i_11_n_0 : STD_LOGIC;
  signal W_26_15_i_12_n_0 : STD_LOGIC;
  signal W_26_15_i_13_n_0 : STD_LOGIC;
  signal W_26_15_i_14_n_0 : STD_LOGIC;
  signal W_26_15_i_15_n_0 : STD_LOGIC;
  signal W_26_15_i_16_n_0 : STD_LOGIC;
  signal W_26_15_i_17_n_0 : STD_LOGIC;
  signal W_26_15_i_2_n_0 : STD_LOGIC;
  signal W_26_15_i_3_n_0 : STD_LOGIC;
  signal W_26_15_i_4_n_0 : STD_LOGIC;
  signal W_26_15_i_5_n_0 : STD_LOGIC;
  signal W_26_15_i_6_n_0 : STD_LOGIC;
  signal W_26_15_i_7_n_0 : STD_LOGIC;
  signal W_26_15_i_8_n_0 : STD_LOGIC;
  signal W_26_15_i_9_n_0 : STD_LOGIC;
  signal W_26_19_i_10_n_0 : STD_LOGIC;
  signal W_26_19_i_11_n_0 : STD_LOGIC;
  signal W_26_19_i_12_n_0 : STD_LOGIC;
  signal W_26_19_i_13_n_0 : STD_LOGIC;
  signal W_26_19_i_14_n_0 : STD_LOGIC;
  signal W_26_19_i_15_n_0 : STD_LOGIC;
  signal W_26_19_i_16_n_0 : STD_LOGIC;
  signal W_26_19_i_17_n_0 : STD_LOGIC;
  signal W_26_19_i_2_n_0 : STD_LOGIC;
  signal W_26_19_i_3_n_0 : STD_LOGIC;
  signal W_26_19_i_4_n_0 : STD_LOGIC;
  signal W_26_19_i_5_n_0 : STD_LOGIC;
  signal W_26_19_i_6_n_0 : STD_LOGIC;
  signal W_26_19_i_7_n_0 : STD_LOGIC;
  signal W_26_19_i_8_n_0 : STD_LOGIC;
  signal W_26_19_i_9_n_0 : STD_LOGIC;
  signal W_26_23_i_10_n_0 : STD_LOGIC;
  signal W_26_23_i_11_n_0 : STD_LOGIC;
  signal W_26_23_i_12_n_0 : STD_LOGIC;
  signal W_26_23_i_13_n_0 : STD_LOGIC;
  signal W_26_23_i_14_n_0 : STD_LOGIC;
  signal W_26_23_i_15_n_0 : STD_LOGIC;
  signal W_26_23_i_16_n_0 : STD_LOGIC;
  signal W_26_23_i_17_n_0 : STD_LOGIC;
  signal W_26_23_i_2_n_0 : STD_LOGIC;
  signal W_26_23_i_3_n_0 : STD_LOGIC;
  signal W_26_23_i_4_n_0 : STD_LOGIC;
  signal W_26_23_i_5_n_0 : STD_LOGIC;
  signal W_26_23_i_6_n_0 : STD_LOGIC;
  signal W_26_23_i_7_n_0 : STD_LOGIC;
  signal W_26_23_i_8_n_0 : STD_LOGIC;
  signal W_26_23_i_9_n_0 : STD_LOGIC;
  signal W_26_27_i_10_n_0 : STD_LOGIC;
  signal W_26_27_i_11_n_0 : STD_LOGIC;
  signal W_26_27_i_12_n_0 : STD_LOGIC;
  signal W_26_27_i_13_n_0 : STD_LOGIC;
  signal W_26_27_i_14_n_0 : STD_LOGIC;
  signal W_26_27_i_15_n_0 : STD_LOGIC;
  signal W_26_27_i_16_n_0 : STD_LOGIC;
  signal W_26_27_i_17_n_0 : STD_LOGIC;
  signal W_26_27_i_2_n_0 : STD_LOGIC;
  signal W_26_27_i_3_n_0 : STD_LOGIC;
  signal W_26_27_i_4_n_0 : STD_LOGIC;
  signal W_26_27_i_5_n_0 : STD_LOGIC;
  signal W_26_27_i_6_n_0 : STD_LOGIC;
  signal W_26_27_i_7_n_0 : STD_LOGIC;
  signal W_26_27_i_8_n_0 : STD_LOGIC;
  signal W_26_27_i_9_n_0 : STD_LOGIC;
  signal W_26_31_i_10_n_0 : STD_LOGIC;
  signal W_26_31_i_11_n_0 : STD_LOGIC;
  signal W_26_31_i_12_n_0 : STD_LOGIC;
  signal W_26_31_i_13_n_0 : STD_LOGIC;
  signal W_26_31_i_14_n_0 : STD_LOGIC;
  signal W_26_31_i_15_n_0 : STD_LOGIC;
  signal W_26_31_i_17_n_0 : STD_LOGIC;
  signal W_26_31_i_19_n_0 : STD_LOGIC;
  signal W_26_31_i_2_n_0 : STD_LOGIC;
  signal W_26_31_i_3_n_0 : STD_LOGIC;
  signal W_26_31_i_4_n_0 : STD_LOGIC;
  signal W_26_31_i_5_n_0 : STD_LOGIC;
  signal W_26_31_i_6_n_0 : STD_LOGIC;
  signal W_26_31_i_7_n_0 : STD_LOGIC;
  signal W_26_31_i_8_n_0 : STD_LOGIC;
  signal W_26_31_i_9_n_0 : STD_LOGIC;
  signal W_26_3_i_10_n_0 : STD_LOGIC;
  signal W_26_3_i_11_n_0 : STD_LOGIC;
  signal W_26_3_i_2_n_0 : STD_LOGIC;
  signal W_26_3_i_3_n_0 : STD_LOGIC;
  signal W_26_3_i_4_n_0 : STD_LOGIC;
  signal W_26_3_i_5_n_0 : STD_LOGIC;
  signal W_26_3_i_6_n_0 : STD_LOGIC;
  signal W_26_3_i_7_n_0 : STD_LOGIC;
  signal W_26_3_i_8_n_0 : STD_LOGIC;
  signal W_26_3_i_9_n_0 : STD_LOGIC;
  signal W_26_7_i_10_n_0 : STD_LOGIC;
  signal W_26_7_i_11_n_0 : STD_LOGIC;
  signal W_26_7_i_12_n_0 : STD_LOGIC;
  signal W_26_7_i_13_n_0 : STD_LOGIC;
  signal W_26_7_i_14_n_0 : STD_LOGIC;
  signal W_26_7_i_15_n_0 : STD_LOGIC;
  signal W_26_7_i_16_n_0 : STD_LOGIC;
  signal W_26_7_i_17_n_0 : STD_LOGIC;
  signal W_26_7_i_2_n_0 : STD_LOGIC;
  signal W_26_7_i_3_n_0 : STD_LOGIC;
  signal W_26_7_i_4_n_0 : STD_LOGIC;
  signal W_26_7_i_5_n_0 : STD_LOGIC;
  signal W_26_7_i_6_n_0 : STD_LOGIC;
  signal W_26_7_i_7_n_0 : STD_LOGIC;
  signal W_26_7_i_8_n_0 : STD_LOGIC;
  signal W_26_7_i_9_n_0 : STD_LOGIC;
  signal W_27_11_i_10_n_0 : STD_LOGIC;
  signal W_27_11_i_11_n_0 : STD_LOGIC;
  signal W_27_11_i_12_n_0 : STD_LOGIC;
  signal W_27_11_i_13_n_0 : STD_LOGIC;
  signal W_27_11_i_14_n_0 : STD_LOGIC;
  signal W_27_11_i_15_n_0 : STD_LOGIC;
  signal W_27_11_i_16_n_0 : STD_LOGIC;
  signal W_27_11_i_17_n_0 : STD_LOGIC;
  signal W_27_11_i_2_n_0 : STD_LOGIC;
  signal W_27_11_i_3_n_0 : STD_LOGIC;
  signal W_27_11_i_4_n_0 : STD_LOGIC;
  signal W_27_11_i_5_n_0 : STD_LOGIC;
  signal W_27_11_i_6_n_0 : STD_LOGIC;
  signal W_27_11_i_7_n_0 : STD_LOGIC;
  signal W_27_11_i_8_n_0 : STD_LOGIC;
  signal W_27_11_i_9_n_0 : STD_LOGIC;
  signal W_27_15_i_10_n_0 : STD_LOGIC;
  signal W_27_15_i_11_n_0 : STD_LOGIC;
  signal W_27_15_i_12_n_0 : STD_LOGIC;
  signal W_27_15_i_13_n_0 : STD_LOGIC;
  signal W_27_15_i_14_n_0 : STD_LOGIC;
  signal W_27_15_i_15_n_0 : STD_LOGIC;
  signal W_27_15_i_16_n_0 : STD_LOGIC;
  signal W_27_15_i_17_n_0 : STD_LOGIC;
  signal W_27_15_i_2_n_0 : STD_LOGIC;
  signal W_27_15_i_3_n_0 : STD_LOGIC;
  signal W_27_15_i_4_n_0 : STD_LOGIC;
  signal W_27_15_i_5_n_0 : STD_LOGIC;
  signal W_27_15_i_6_n_0 : STD_LOGIC;
  signal W_27_15_i_7_n_0 : STD_LOGIC;
  signal W_27_15_i_8_n_0 : STD_LOGIC;
  signal W_27_15_i_9_n_0 : STD_LOGIC;
  signal W_27_19_i_10_n_0 : STD_LOGIC;
  signal W_27_19_i_11_n_0 : STD_LOGIC;
  signal W_27_19_i_12_n_0 : STD_LOGIC;
  signal W_27_19_i_13_n_0 : STD_LOGIC;
  signal W_27_19_i_14_n_0 : STD_LOGIC;
  signal W_27_19_i_15_n_0 : STD_LOGIC;
  signal W_27_19_i_16_n_0 : STD_LOGIC;
  signal W_27_19_i_17_n_0 : STD_LOGIC;
  signal W_27_19_i_2_n_0 : STD_LOGIC;
  signal W_27_19_i_3_n_0 : STD_LOGIC;
  signal W_27_19_i_4_n_0 : STD_LOGIC;
  signal W_27_19_i_5_n_0 : STD_LOGIC;
  signal W_27_19_i_6_n_0 : STD_LOGIC;
  signal W_27_19_i_7_n_0 : STD_LOGIC;
  signal W_27_19_i_8_n_0 : STD_LOGIC;
  signal W_27_19_i_9_n_0 : STD_LOGIC;
  signal W_27_23_i_10_n_0 : STD_LOGIC;
  signal W_27_23_i_11_n_0 : STD_LOGIC;
  signal W_27_23_i_12_n_0 : STD_LOGIC;
  signal W_27_23_i_13_n_0 : STD_LOGIC;
  signal W_27_23_i_14_n_0 : STD_LOGIC;
  signal W_27_23_i_15_n_0 : STD_LOGIC;
  signal W_27_23_i_16_n_0 : STD_LOGIC;
  signal W_27_23_i_17_n_0 : STD_LOGIC;
  signal W_27_23_i_2_n_0 : STD_LOGIC;
  signal W_27_23_i_3_n_0 : STD_LOGIC;
  signal W_27_23_i_4_n_0 : STD_LOGIC;
  signal W_27_23_i_5_n_0 : STD_LOGIC;
  signal W_27_23_i_6_n_0 : STD_LOGIC;
  signal W_27_23_i_7_n_0 : STD_LOGIC;
  signal W_27_23_i_8_n_0 : STD_LOGIC;
  signal W_27_23_i_9_n_0 : STD_LOGIC;
  signal W_27_27_i_10_n_0 : STD_LOGIC;
  signal W_27_27_i_11_n_0 : STD_LOGIC;
  signal W_27_27_i_12_n_0 : STD_LOGIC;
  signal W_27_27_i_13_n_0 : STD_LOGIC;
  signal W_27_27_i_14_n_0 : STD_LOGIC;
  signal W_27_27_i_15_n_0 : STD_LOGIC;
  signal W_27_27_i_16_n_0 : STD_LOGIC;
  signal W_27_27_i_17_n_0 : STD_LOGIC;
  signal W_27_27_i_2_n_0 : STD_LOGIC;
  signal W_27_27_i_3_n_0 : STD_LOGIC;
  signal W_27_27_i_4_n_0 : STD_LOGIC;
  signal W_27_27_i_5_n_0 : STD_LOGIC;
  signal W_27_27_i_6_n_0 : STD_LOGIC;
  signal W_27_27_i_7_n_0 : STD_LOGIC;
  signal W_27_27_i_8_n_0 : STD_LOGIC;
  signal W_27_27_i_9_n_0 : STD_LOGIC;
  signal W_27_31_i_10_n_0 : STD_LOGIC;
  signal W_27_31_i_11_n_0 : STD_LOGIC;
  signal W_27_31_i_12_n_0 : STD_LOGIC;
  signal W_27_31_i_13_n_0 : STD_LOGIC;
  signal W_27_31_i_14_n_0 : STD_LOGIC;
  signal W_27_31_i_15_n_0 : STD_LOGIC;
  signal W_27_31_i_17_n_0 : STD_LOGIC;
  signal W_27_31_i_19_n_0 : STD_LOGIC;
  signal W_27_31_i_2_n_0 : STD_LOGIC;
  signal W_27_31_i_3_n_0 : STD_LOGIC;
  signal W_27_31_i_4_n_0 : STD_LOGIC;
  signal W_27_31_i_5_n_0 : STD_LOGIC;
  signal W_27_31_i_6_n_0 : STD_LOGIC;
  signal W_27_31_i_7_n_0 : STD_LOGIC;
  signal W_27_31_i_8_n_0 : STD_LOGIC;
  signal W_27_31_i_9_n_0 : STD_LOGIC;
  signal W_27_3_i_10_n_0 : STD_LOGIC;
  signal W_27_3_i_11_n_0 : STD_LOGIC;
  signal W_27_3_i_2_n_0 : STD_LOGIC;
  signal W_27_3_i_3_n_0 : STD_LOGIC;
  signal W_27_3_i_4_n_0 : STD_LOGIC;
  signal W_27_3_i_5_n_0 : STD_LOGIC;
  signal W_27_3_i_6_n_0 : STD_LOGIC;
  signal W_27_3_i_7_n_0 : STD_LOGIC;
  signal W_27_3_i_8_n_0 : STD_LOGIC;
  signal W_27_3_i_9_n_0 : STD_LOGIC;
  signal W_27_7_i_10_n_0 : STD_LOGIC;
  signal W_27_7_i_11_n_0 : STD_LOGIC;
  signal W_27_7_i_12_n_0 : STD_LOGIC;
  signal W_27_7_i_13_n_0 : STD_LOGIC;
  signal W_27_7_i_14_n_0 : STD_LOGIC;
  signal W_27_7_i_15_n_0 : STD_LOGIC;
  signal W_27_7_i_16_n_0 : STD_LOGIC;
  signal W_27_7_i_17_n_0 : STD_LOGIC;
  signal W_27_7_i_2_n_0 : STD_LOGIC;
  signal W_27_7_i_3_n_0 : STD_LOGIC;
  signal W_27_7_i_4_n_0 : STD_LOGIC;
  signal W_27_7_i_5_n_0 : STD_LOGIC;
  signal W_27_7_i_6_n_0 : STD_LOGIC;
  signal W_27_7_i_7_n_0 : STD_LOGIC;
  signal W_27_7_i_8_n_0 : STD_LOGIC;
  signal W_27_7_i_9_n_0 : STD_LOGIC;
  signal W_28_11_i_10_n_0 : STD_LOGIC;
  signal W_28_11_i_11_n_0 : STD_LOGIC;
  signal W_28_11_i_12_n_0 : STD_LOGIC;
  signal W_28_11_i_13_n_0 : STD_LOGIC;
  signal W_28_11_i_14_n_0 : STD_LOGIC;
  signal W_28_11_i_15_n_0 : STD_LOGIC;
  signal W_28_11_i_16_n_0 : STD_LOGIC;
  signal W_28_11_i_17_n_0 : STD_LOGIC;
  signal W_28_11_i_2_n_0 : STD_LOGIC;
  signal W_28_11_i_3_n_0 : STD_LOGIC;
  signal W_28_11_i_4_n_0 : STD_LOGIC;
  signal W_28_11_i_5_n_0 : STD_LOGIC;
  signal W_28_11_i_6_n_0 : STD_LOGIC;
  signal W_28_11_i_7_n_0 : STD_LOGIC;
  signal W_28_11_i_8_n_0 : STD_LOGIC;
  signal W_28_11_i_9_n_0 : STD_LOGIC;
  signal W_28_15_i_10_n_0 : STD_LOGIC;
  signal W_28_15_i_11_n_0 : STD_LOGIC;
  signal W_28_15_i_12_n_0 : STD_LOGIC;
  signal W_28_15_i_13_n_0 : STD_LOGIC;
  signal W_28_15_i_14_n_0 : STD_LOGIC;
  signal W_28_15_i_15_n_0 : STD_LOGIC;
  signal W_28_15_i_16_n_0 : STD_LOGIC;
  signal W_28_15_i_17_n_0 : STD_LOGIC;
  signal W_28_15_i_2_n_0 : STD_LOGIC;
  signal W_28_15_i_3_n_0 : STD_LOGIC;
  signal W_28_15_i_4_n_0 : STD_LOGIC;
  signal W_28_15_i_5_n_0 : STD_LOGIC;
  signal W_28_15_i_6_n_0 : STD_LOGIC;
  signal W_28_15_i_7_n_0 : STD_LOGIC;
  signal W_28_15_i_8_n_0 : STD_LOGIC;
  signal W_28_15_i_9_n_0 : STD_LOGIC;
  signal W_28_19_i_10_n_0 : STD_LOGIC;
  signal W_28_19_i_11_n_0 : STD_LOGIC;
  signal W_28_19_i_12_n_0 : STD_LOGIC;
  signal W_28_19_i_13_n_0 : STD_LOGIC;
  signal W_28_19_i_14_n_0 : STD_LOGIC;
  signal W_28_19_i_15_n_0 : STD_LOGIC;
  signal W_28_19_i_16_n_0 : STD_LOGIC;
  signal W_28_19_i_17_n_0 : STD_LOGIC;
  signal W_28_19_i_2_n_0 : STD_LOGIC;
  signal W_28_19_i_3_n_0 : STD_LOGIC;
  signal W_28_19_i_4_n_0 : STD_LOGIC;
  signal W_28_19_i_5_n_0 : STD_LOGIC;
  signal W_28_19_i_6_n_0 : STD_LOGIC;
  signal W_28_19_i_7_n_0 : STD_LOGIC;
  signal W_28_19_i_8_n_0 : STD_LOGIC;
  signal W_28_19_i_9_n_0 : STD_LOGIC;
  signal W_28_23_i_10_n_0 : STD_LOGIC;
  signal W_28_23_i_11_n_0 : STD_LOGIC;
  signal W_28_23_i_12_n_0 : STD_LOGIC;
  signal W_28_23_i_13_n_0 : STD_LOGIC;
  signal W_28_23_i_14_n_0 : STD_LOGIC;
  signal W_28_23_i_15_n_0 : STD_LOGIC;
  signal W_28_23_i_16_n_0 : STD_LOGIC;
  signal W_28_23_i_17_n_0 : STD_LOGIC;
  signal W_28_23_i_2_n_0 : STD_LOGIC;
  signal W_28_23_i_3_n_0 : STD_LOGIC;
  signal W_28_23_i_4_n_0 : STD_LOGIC;
  signal W_28_23_i_5_n_0 : STD_LOGIC;
  signal W_28_23_i_6_n_0 : STD_LOGIC;
  signal W_28_23_i_7_n_0 : STD_LOGIC;
  signal W_28_23_i_8_n_0 : STD_LOGIC;
  signal W_28_23_i_9_n_0 : STD_LOGIC;
  signal W_28_27_i_10_n_0 : STD_LOGIC;
  signal W_28_27_i_11_n_0 : STD_LOGIC;
  signal W_28_27_i_12_n_0 : STD_LOGIC;
  signal W_28_27_i_13_n_0 : STD_LOGIC;
  signal W_28_27_i_14_n_0 : STD_LOGIC;
  signal W_28_27_i_15_n_0 : STD_LOGIC;
  signal W_28_27_i_16_n_0 : STD_LOGIC;
  signal W_28_27_i_17_n_0 : STD_LOGIC;
  signal W_28_27_i_2_n_0 : STD_LOGIC;
  signal W_28_27_i_3_n_0 : STD_LOGIC;
  signal W_28_27_i_4_n_0 : STD_LOGIC;
  signal W_28_27_i_5_n_0 : STD_LOGIC;
  signal W_28_27_i_6_n_0 : STD_LOGIC;
  signal W_28_27_i_7_n_0 : STD_LOGIC;
  signal W_28_27_i_8_n_0 : STD_LOGIC;
  signal W_28_27_i_9_n_0 : STD_LOGIC;
  signal W_28_31_i_10_n_0 : STD_LOGIC;
  signal W_28_31_i_11_n_0 : STD_LOGIC;
  signal W_28_31_i_12_n_0 : STD_LOGIC;
  signal W_28_31_i_13_n_0 : STD_LOGIC;
  signal W_28_31_i_14_n_0 : STD_LOGIC;
  signal W_28_31_i_15_n_0 : STD_LOGIC;
  signal W_28_31_i_17_n_0 : STD_LOGIC;
  signal W_28_31_i_19_n_0 : STD_LOGIC;
  signal W_28_31_i_2_n_0 : STD_LOGIC;
  signal W_28_31_i_3_n_0 : STD_LOGIC;
  signal W_28_31_i_4_n_0 : STD_LOGIC;
  signal W_28_31_i_5_n_0 : STD_LOGIC;
  signal W_28_31_i_6_n_0 : STD_LOGIC;
  signal W_28_31_i_7_n_0 : STD_LOGIC;
  signal W_28_31_i_8_n_0 : STD_LOGIC;
  signal W_28_31_i_9_n_0 : STD_LOGIC;
  signal W_28_3_i_10_n_0 : STD_LOGIC;
  signal W_28_3_i_11_n_0 : STD_LOGIC;
  signal W_28_3_i_2_n_0 : STD_LOGIC;
  signal W_28_3_i_3_n_0 : STD_LOGIC;
  signal W_28_3_i_4_n_0 : STD_LOGIC;
  signal W_28_3_i_5_n_0 : STD_LOGIC;
  signal W_28_3_i_6_n_0 : STD_LOGIC;
  signal W_28_3_i_7_n_0 : STD_LOGIC;
  signal W_28_3_i_8_n_0 : STD_LOGIC;
  signal W_28_3_i_9_n_0 : STD_LOGIC;
  signal W_28_7_i_10_n_0 : STD_LOGIC;
  signal W_28_7_i_11_n_0 : STD_LOGIC;
  signal W_28_7_i_12_n_0 : STD_LOGIC;
  signal W_28_7_i_13_n_0 : STD_LOGIC;
  signal W_28_7_i_14_n_0 : STD_LOGIC;
  signal W_28_7_i_15_n_0 : STD_LOGIC;
  signal W_28_7_i_16_n_0 : STD_LOGIC;
  signal W_28_7_i_17_n_0 : STD_LOGIC;
  signal W_28_7_i_2_n_0 : STD_LOGIC;
  signal W_28_7_i_3_n_0 : STD_LOGIC;
  signal W_28_7_i_4_n_0 : STD_LOGIC;
  signal W_28_7_i_5_n_0 : STD_LOGIC;
  signal W_28_7_i_6_n_0 : STD_LOGIC;
  signal W_28_7_i_7_n_0 : STD_LOGIC;
  signal W_28_7_i_8_n_0 : STD_LOGIC;
  signal W_28_7_i_9_n_0 : STD_LOGIC;
  signal W_29_11_i_10_n_0 : STD_LOGIC;
  signal W_29_11_i_11_n_0 : STD_LOGIC;
  signal W_29_11_i_12_n_0 : STD_LOGIC;
  signal W_29_11_i_13_n_0 : STD_LOGIC;
  signal W_29_11_i_14_n_0 : STD_LOGIC;
  signal W_29_11_i_15_n_0 : STD_LOGIC;
  signal W_29_11_i_16_n_0 : STD_LOGIC;
  signal W_29_11_i_17_n_0 : STD_LOGIC;
  signal W_29_11_i_2_n_0 : STD_LOGIC;
  signal W_29_11_i_3_n_0 : STD_LOGIC;
  signal W_29_11_i_4_n_0 : STD_LOGIC;
  signal W_29_11_i_5_n_0 : STD_LOGIC;
  signal W_29_11_i_6_n_0 : STD_LOGIC;
  signal W_29_11_i_7_n_0 : STD_LOGIC;
  signal W_29_11_i_8_n_0 : STD_LOGIC;
  signal W_29_11_i_9_n_0 : STD_LOGIC;
  signal W_29_15_i_10_n_0 : STD_LOGIC;
  signal W_29_15_i_11_n_0 : STD_LOGIC;
  signal W_29_15_i_12_n_0 : STD_LOGIC;
  signal W_29_15_i_13_n_0 : STD_LOGIC;
  signal W_29_15_i_14_n_0 : STD_LOGIC;
  signal W_29_15_i_15_n_0 : STD_LOGIC;
  signal W_29_15_i_16_n_0 : STD_LOGIC;
  signal W_29_15_i_17_n_0 : STD_LOGIC;
  signal W_29_15_i_2_n_0 : STD_LOGIC;
  signal W_29_15_i_3_n_0 : STD_LOGIC;
  signal W_29_15_i_4_n_0 : STD_LOGIC;
  signal W_29_15_i_5_n_0 : STD_LOGIC;
  signal W_29_15_i_6_n_0 : STD_LOGIC;
  signal W_29_15_i_7_n_0 : STD_LOGIC;
  signal W_29_15_i_8_n_0 : STD_LOGIC;
  signal W_29_15_i_9_n_0 : STD_LOGIC;
  signal W_29_19_i_10_n_0 : STD_LOGIC;
  signal W_29_19_i_11_n_0 : STD_LOGIC;
  signal W_29_19_i_12_n_0 : STD_LOGIC;
  signal W_29_19_i_13_n_0 : STD_LOGIC;
  signal W_29_19_i_14_n_0 : STD_LOGIC;
  signal W_29_19_i_15_n_0 : STD_LOGIC;
  signal W_29_19_i_16_n_0 : STD_LOGIC;
  signal W_29_19_i_17_n_0 : STD_LOGIC;
  signal W_29_19_i_2_n_0 : STD_LOGIC;
  signal W_29_19_i_3_n_0 : STD_LOGIC;
  signal W_29_19_i_4_n_0 : STD_LOGIC;
  signal W_29_19_i_5_n_0 : STD_LOGIC;
  signal W_29_19_i_6_n_0 : STD_LOGIC;
  signal W_29_19_i_7_n_0 : STD_LOGIC;
  signal W_29_19_i_8_n_0 : STD_LOGIC;
  signal W_29_19_i_9_n_0 : STD_LOGIC;
  signal W_29_23_i_10_n_0 : STD_LOGIC;
  signal W_29_23_i_11_n_0 : STD_LOGIC;
  signal W_29_23_i_12_n_0 : STD_LOGIC;
  signal W_29_23_i_13_n_0 : STD_LOGIC;
  signal W_29_23_i_14_n_0 : STD_LOGIC;
  signal W_29_23_i_15_n_0 : STD_LOGIC;
  signal W_29_23_i_16_n_0 : STD_LOGIC;
  signal W_29_23_i_17_n_0 : STD_LOGIC;
  signal W_29_23_i_2_n_0 : STD_LOGIC;
  signal W_29_23_i_3_n_0 : STD_LOGIC;
  signal W_29_23_i_4_n_0 : STD_LOGIC;
  signal W_29_23_i_5_n_0 : STD_LOGIC;
  signal W_29_23_i_6_n_0 : STD_LOGIC;
  signal W_29_23_i_7_n_0 : STD_LOGIC;
  signal W_29_23_i_8_n_0 : STD_LOGIC;
  signal W_29_23_i_9_n_0 : STD_LOGIC;
  signal W_29_27_i_10_n_0 : STD_LOGIC;
  signal W_29_27_i_11_n_0 : STD_LOGIC;
  signal W_29_27_i_12_n_0 : STD_LOGIC;
  signal W_29_27_i_13_n_0 : STD_LOGIC;
  signal W_29_27_i_14_n_0 : STD_LOGIC;
  signal W_29_27_i_15_n_0 : STD_LOGIC;
  signal W_29_27_i_16_n_0 : STD_LOGIC;
  signal W_29_27_i_17_n_0 : STD_LOGIC;
  signal W_29_27_i_2_n_0 : STD_LOGIC;
  signal W_29_27_i_3_n_0 : STD_LOGIC;
  signal W_29_27_i_4_n_0 : STD_LOGIC;
  signal W_29_27_i_5_n_0 : STD_LOGIC;
  signal W_29_27_i_6_n_0 : STD_LOGIC;
  signal W_29_27_i_7_n_0 : STD_LOGIC;
  signal W_29_27_i_8_n_0 : STD_LOGIC;
  signal W_29_27_i_9_n_0 : STD_LOGIC;
  signal W_29_31_i_10_n_0 : STD_LOGIC;
  signal W_29_31_i_11_n_0 : STD_LOGIC;
  signal W_29_31_i_12_n_0 : STD_LOGIC;
  signal W_29_31_i_13_n_0 : STD_LOGIC;
  signal W_29_31_i_14_n_0 : STD_LOGIC;
  signal W_29_31_i_15_n_0 : STD_LOGIC;
  signal W_29_31_i_17_n_0 : STD_LOGIC;
  signal W_29_31_i_19_n_0 : STD_LOGIC;
  signal W_29_31_i_2_n_0 : STD_LOGIC;
  signal W_29_31_i_3_n_0 : STD_LOGIC;
  signal W_29_31_i_4_n_0 : STD_LOGIC;
  signal W_29_31_i_5_n_0 : STD_LOGIC;
  signal W_29_31_i_6_n_0 : STD_LOGIC;
  signal W_29_31_i_7_n_0 : STD_LOGIC;
  signal W_29_31_i_8_n_0 : STD_LOGIC;
  signal W_29_31_i_9_n_0 : STD_LOGIC;
  signal W_29_3_i_10_n_0 : STD_LOGIC;
  signal W_29_3_i_11_n_0 : STD_LOGIC;
  signal W_29_3_i_2_n_0 : STD_LOGIC;
  signal W_29_3_i_3_n_0 : STD_LOGIC;
  signal W_29_3_i_4_n_0 : STD_LOGIC;
  signal W_29_3_i_5_n_0 : STD_LOGIC;
  signal W_29_3_i_6_n_0 : STD_LOGIC;
  signal W_29_3_i_7_n_0 : STD_LOGIC;
  signal W_29_3_i_8_n_0 : STD_LOGIC;
  signal W_29_3_i_9_n_0 : STD_LOGIC;
  signal W_29_7_i_10_n_0 : STD_LOGIC;
  signal W_29_7_i_11_n_0 : STD_LOGIC;
  signal W_29_7_i_12_n_0 : STD_LOGIC;
  signal W_29_7_i_13_n_0 : STD_LOGIC;
  signal W_29_7_i_14_n_0 : STD_LOGIC;
  signal W_29_7_i_15_n_0 : STD_LOGIC;
  signal W_29_7_i_16_n_0 : STD_LOGIC;
  signal W_29_7_i_17_n_0 : STD_LOGIC;
  signal W_29_7_i_2_n_0 : STD_LOGIC;
  signal W_29_7_i_3_n_0 : STD_LOGIC;
  signal W_29_7_i_4_n_0 : STD_LOGIC;
  signal W_29_7_i_5_n_0 : STD_LOGIC;
  signal W_29_7_i_6_n_0 : STD_LOGIC;
  signal W_29_7_i_7_n_0 : STD_LOGIC;
  signal W_29_7_i_8_n_0 : STD_LOGIC;
  signal W_29_7_i_9_n_0 : STD_LOGIC;
  signal W_30_11_i_10_n_0 : STD_LOGIC;
  signal W_30_11_i_11_n_0 : STD_LOGIC;
  signal W_30_11_i_12_n_0 : STD_LOGIC;
  signal W_30_11_i_13_n_0 : STD_LOGIC;
  signal W_30_11_i_14_n_0 : STD_LOGIC;
  signal W_30_11_i_15_n_0 : STD_LOGIC;
  signal W_30_11_i_16_n_0 : STD_LOGIC;
  signal W_30_11_i_17_n_0 : STD_LOGIC;
  signal W_30_11_i_2_n_0 : STD_LOGIC;
  signal W_30_11_i_3_n_0 : STD_LOGIC;
  signal W_30_11_i_4_n_0 : STD_LOGIC;
  signal W_30_11_i_5_n_0 : STD_LOGIC;
  signal W_30_11_i_6_n_0 : STD_LOGIC;
  signal W_30_11_i_7_n_0 : STD_LOGIC;
  signal W_30_11_i_8_n_0 : STD_LOGIC;
  signal W_30_11_i_9_n_0 : STD_LOGIC;
  signal W_30_15_i_10_n_0 : STD_LOGIC;
  signal W_30_15_i_11_n_0 : STD_LOGIC;
  signal W_30_15_i_12_n_0 : STD_LOGIC;
  signal W_30_15_i_13_n_0 : STD_LOGIC;
  signal W_30_15_i_14_n_0 : STD_LOGIC;
  signal W_30_15_i_15_n_0 : STD_LOGIC;
  signal W_30_15_i_16_n_0 : STD_LOGIC;
  signal W_30_15_i_17_n_0 : STD_LOGIC;
  signal W_30_15_i_2_n_0 : STD_LOGIC;
  signal W_30_15_i_3_n_0 : STD_LOGIC;
  signal W_30_15_i_4_n_0 : STD_LOGIC;
  signal W_30_15_i_5_n_0 : STD_LOGIC;
  signal W_30_15_i_6_n_0 : STD_LOGIC;
  signal W_30_15_i_7_n_0 : STD_LOGIC;
  signal W_30_15_i_8_n_0 : STD_LOGIC;
  signal W_30_15_i_9_n_0 : STD_LOGIC;
  signal W_30_19_i_10_n_0 : STD_LOGIC;
  signal W_30_19_i_11_n_0 : STD_LOGIC;
  signal W_30_19_i_12_n_0 : STD_LOGIC;
  signal W_30_19_i_13_n_0 : STD_LOGIC;
  signal W_30_19_i_14_n_0 : STD_LOGIC;
  signal W_30_19_i_15_n_0 : STD_LOGIC;
  signal W_30_19_i_16_n_0 : STD_LOGIC;
  signal W_30_19_i_17_n_0 : STD_LOGIC;
  signal W_30_19_i_2_n_0 : STD_LOGIC;
  signal W_30_19_i_3_n_0 : STD_LOGIC;
  signal W_30_19_i_4_n_0 : STD_LOGIC;
  signal W_30_19_i_5_n_0 : STD_LOGIC;
  signal W_30_19_i_6_n_0 : STD_LOGIC;
  signal W_30_19_i_7_n_0 : STD_LOGIC;
  signal W_30_19_i_8_n_0 : STD_LOGIC;
  signal W_30_19_i_9_n_0 : STD_LOGIC;
  signal W_30_23_i_10_n_0 : STD_LOGIC;
  signal W_30_23_i_11_n_0 : STD_LOGIC;
  signal W_30_23_i_12_n_0 : STD_LOGIC;
  signal W_30_23_i_13_n_0 : STD_LOGIC;
  signal W_30_23_i_14_n_0 : STD_LOGIC;
  signal W_30_23_i_15_n_0 : STD_LOGIC;
  signal W_30_23_i_16_n_0 : STD_LOGIC;
  signal W_30_23_i_17_n_0 : STD_LOGIC;
  signal W_30_23_i_2_n_0 : STD_LOGIC;
  signal W_30_23_i_3_n_0 : STD_LOGIC;
  signal W_30_23_i_4_n_0 : STD_LOGIC;
  signal W_30_23_i_5_n_0 : STD_LOGIC;
  signal W_30_23_i_6_n_0 : STD_LOGIC;
  signal W_30_23_i_7_n_0 : STD_LOGIC;
  signal W_30_23_i_8_n_0 : STD_LOGIC;
  signal W_30_23_i_9_n_0 : STD_LOGIC;
  signal W_30_27_i_10_n_0 : STD_LOGIC;
  signal W_30_27_i_11_n_0 : STD_LOGIC;
  signal W_30_27_i_12_n_0 : STD_LOGIC;
  signal W_30_27_i_13_n_0 : STD_LOGIC;
  signal W_30_27_i_14_n_0 : STD_LOGIC;
  signal W_30_27_i_15_n_0 : STD_LOGIC;
  signal W_30_27_i_16_n_0 : STD_LOGIC;
  signal W_30_27_i_17_n_0 : STD_LOGIC;
  signal W_30_27_i_2_n_0 : STD_LOGIC;
  signal W_30_27_i_3_n_0 : STD_LOGIC;
  signal W_30_27_i_4_n_0 : STD_LOGIC;
  signal W_30_27_i_5_n_0 : STD_LOGIC;
  signal W_30_27_i_6_n_0 : STD_LOGIC;
  signal W_30_27_i_7_n_0 : STD_LOGIC;
  signal W_30_27_i_8_n_0 : STD_LOGIC;
  signal W_30_27_i_9_n_0 : STD_LOGIC;
  signal W_30_31_i_10_n_0 : STD_LOGIC;
  signal W_30_31_i_11_n_0 : STD_LOGIC;
  signal W_30_31_i_12_n_0 : STD_LOGIC;
  signal W_30_31_i_13_n_0 : STD_LOGIC;
  signal W_30_31_i_14_n_0 : STD_LOGIC;
  signal W_30_31_i_15_n_0 : STD_LOGIC;
  signal W_30_31_i_17_n_0 : STD_LOGIC;
  signal W_30_31_i_19_n_0 : STD_LOGIC;
  signal W_30_31_i_2_n_0 : STD_LOGIC;
  signal W_30_31_i_3_n_0 : STD_LOGIC;
  signal W_30_31_i_4_n_0 : STD_LOGIC;
  signal W_30_31_i_5_n_0 : STD_LOGIC;
  signal W_30_31_i_6_n_0 : STD_LOGIC;
  signal W_30_31_i_7_n_0 : STD_LOGIC;
  signal W_30_31_i_8_n_0 : STD_LOGIC;
  signal W_30_31_i_9_n_0 : STD_LOGIC;
  signal W_30_3_i_10_n_0 : STD_LOGIC;
  signal W_30_3_i_11_n_0 : STD_LOGIC;
  signal W_30_3_i_2_n_0 : STD_LOGIC;
  signal W_30_3_i_3_n_0 : STD_LOGIC;
  signal W_30_3_i_4_n_0 : STD_LOGIC;
  signal W_30_3_i_5_n_0 : STD_LOGIC;
  signal W_30_3_i_6_n_0 : STD_LOGIC;
  signal W_30_3_i_7_n_0 : STD_LOGIC;
  signal W_30_3_i_8_n_0 : STD_LOGIC;
  signal W_30_3_i_9_n_0 : STD_LOGIC;
  signal W_30_7_i_10_n_0 : STD_LOGIC;
  signal W_30_7_i_11_n_0 : STD_LOGIC;
  signal W_30_7_i_12_n_0 : STD_LOGIC;
  signal W_30_7_i_13_n_0 : STD_LOGIC;
  signal W_30_7_i_14_n_0 : STD_LOGIC;
  signal W_30_7_i_15_n_0 : STD_LOGIC;
  signal W_30_7_i_16_n_0 : STD_LOGIC;
  signal W_30_7_i_17_n_0 : STD_LOGIC;
  signal W_30_7_i_2_n_0 : STD_LOGIC;
  signal W_30_7_i_3_n_0 : STD_LOGIC;
  signal W_30_7_i_4_n_0 : STD_LOGIC;
  signal W_30_7_i_5_n_0 : STD_LOGIC;
  signal W_30_7_i_6_n_0 : STD_LOGIC;
  signal W_30_7_i_7_n_0 : STD_LOGIC;
  signal W_30_7_i_8_n_0 : STD_LOGIC;
  signal W_30_7_i_9_n_0 : STD_LOGIC;
  signal W_31_11_i_10_n_0 : STD_LOGIC;
  signal W_31_11_i_11_n_0 : STD_LOGIC;
  signal W_31_11_i_12_n_0 : STD_LOGIC;
  signal W_31_11_i_13_n_0 : STD_LOGIC;
  signal W_31_11_i_14_n_0 : STD_LOGIC;
  signal W_31_11_i_15_n_0 : STD_LOGIC;
  signal W_31_11_i_16_n_0 : STD_LOGIC;
  signal W_31_11_i_17_n_0 : STD_LOGIC;
  signal W_31_11_i_2_n_0 : STD_LOGIC;
  signal W_31_11_i_3_n_0 : STD_LOGIC;
  signal W_31_11_i_4_n_0 : STD_LOGIC;
  signal W_31_11_i_5_n_0 : STD_LOGIC;
  signal W_31_11_i_6_n_0 : STD_LOGIC;
  signal W_31_11_i_7_n_0 : STD_LOGIC;
  signal W_31_11_i_8_n_0 : STD_LOGIC;
  signal W_31_11_i_9_n_0 : STD_LOGIC;
  signal W_31_15_i_10_n_0 : STD_LOGIC;
  signal W_31_15_i_11_n_0 : STD_LOGIC;
  signal W_31_15_i_12_n_0 : STD_LOGIC;
  signal W_31_15_i_13_n_0 : STD_LOGIC;
  signal W_31_15_i_14_n_0 : STD_LOGIC;
  signal W_31_15_i_15_n_0 : STD_LOGIC;
  signal W_31_15_i_16_n_0 : STD_LOGIC;
  signal W_31_15_i_17_n_0 : STD_LOGIC;
  signal W_31_15_i_2_n_0 : STD_LOGIC;
  signal W_31_15_i_3_n_0 : STD_LOGIC;
  signal W_31_15_i_4_n_0 : STD_LOGIC;
  signal W_31_15_i_5_n_0 : STD_LOGIC;
  signal W_31_15_i_6_n_0 : STD_LOGIC;
  signal W_31_15_i_7_n_0 : STD_LOGIC;
  signal W_31_15_i_8_n_0 : STD_LOGIC;
  signal W_31_15_i_9_n_0 : STD_LOGIC;
  signal W_31_19_i_10_n_0 : STD_LOGIC;
  signal W_31_19_i_11_n_0 : STD_LOGIC;
  signal W_31_19_i_12_n_0 : STD_LOGIC;
  signal W_31_19_i_13_n_0 : STD_LOGIC;
  signal W_31_19_i_14_n_0 : STD_LOGIC;
  signal W_31_19_i_15_n_0 : STD_LOGIC;
  signal W_31_19_i_16_n_0 : STD_LOGIC;
  signal W_31_19_i_17_n_0 : STD_LOGIC;
  signal W_31_19_i_2_n_0 : STD_LOGIC;
  signal W_31_19_i_3_n_0 : STD_LOGIC;
  signal W_31_19_i_4_n_0 : STD_LOGIC;
  signal W_31_19_i_5_n_0 : STD_LOGIC;
  signal W_31_19_i_6_n_0 : STD_LOGIC;
  signal W_31_19_i_7_n_0 : STD_LOGIC;
  signal W_31_19_i_8_n_0 : STD_LOGIC;
  signal W_31_19_i_9_n_0 : STD_LOGIC;
  signal W_31_23_i_10_n_0 : STD_LOGIC;
  signal W_31_23_i_11_n_0 : STD_LOGIC;
  signal W_31_23_i_12_n_0 : STD_LOGIC;
  signal W_31_23_i_13_n_0 : STD_LOGIC;
  signal W_31_23_i_14_n_0 : STD_LOGIC;
  signal W_31_23_i_15_n_0 : STD_LOGIC;
  signal W_31_23_i_16_n_0 : STD_LOGIC;
  signal W_31_23_i_17_n_0 : STD_LOGIC;
  signal W_31_23_i_2_n_0 : STD_LOGIC;
  signal W_31_23_i_3_n_0 : STD_LOGIC;
  signal W_31_23_i_4_n_0 : STD_LOGIC;
  signal W_31_23_i_5_n_0 : STD_LOGIC;
  signal W_31_23_i_6_n_0 : STD_LOGIC;
  signal W_31_23_i_7_n_0 : STD_LOGIC;
  signal W_31_23_i_8_n_0 : STD_LOGIC;
  signal W_31_23_i_9_n_0 : STD_LOGIC;
  signal W_31_27_i_10_n_0 : STD_LOGIC;
  signal W_31_27_i_11_n_0 : STD_LOGIC;
  signal W_31_27_i_12_n_0 : STD_LOGIC;
  signal W_31_27_i_13_n_0 : STD_LOGIC;
  signal W_31_27_i_14_n_0 : STD_LOGIC;
  signal W_31_27_i_15_n_0 : STD_LOGIC;
  signal W_31_27_i_16_n_0 : STD_LOGIC;
  signal W_31_27_i_17_n_0 : STD_LOGIC;
  signal W_31_27_i_2_n_0 : STD_LOGIC;
  signal W_31_27_i_3_n_0 : STD_LOGIC;
  signal W_31_27_i_4_n_0 : STD_LOGIC;
  signal W_31_27_i_5_n_0 : STD_LOGIC;
  signal W_31_27_i_6_n_0 : STD_LOGIC;
  signal W_31_27_i_7_n_0 : STD_LOGIC;
  signal W_31_27_i_8_n_0 : STD_LOGIC;
  signal W_31_27_i_9_n_0 : STD_LOGIC;
  signal W_31_31_i_10_n_0 : STD_LOGIC;
  signal W_31_31_i_11_n_0 : STD_LOGIC;
  signal W_31_31_i_12_n_0 : STD_LOGIC;
  signal W_31_31_i_13_n_0 : STD_LOGIC;
  signal W_31_31_i_14_n_0 : STD_LOGIC;
  signal W_31_31_i_15_n_0 : STD_LOGIC;
  signal W_31_31_i_17_n_0 : STD_LOGIC;
  signal W_31_31_i_19_n_0 : STD_LOGIC;
  signal W_31_31_i_2_n_0 : STD_LOGIC;
  signal W_31_31_i_3_n_0 : STD_LOGIC;
  signal W_31_31_i_4_n_0 : STD_LOGIC;
  signal W_31_31_i_5_n_0 : STD_LOGIC;
  signal W_31_31_i_6_n_0 : STD_LOGIC;
  signal W_31_31_i_7_n_0 : STD_LOGIC;
  signal W_31_31_i_8_n_0 : STD_LOGIC;
  signal W_31_31_i_9_n_0 : STD_LOGIC;
  signal W_31_3_i_10_n_0 : STD_LOGIC;
  signal W_31_3_i_11_n_0 : STD_LOGIC;
  signal W_31_3_i_15_n_0 : STD_LOGIC;
  signal W_31_3_i_2_n_0 : STD_LOGIC;
  signal W_31_3_i_3_n_0 : STD_LOGIC;
  signal W_31_3_i_4_n_0 : STD_LOGIC;
  signal W_31_3_i_5_n_0 : STD_LOGIC;
  signal W_31_3_i_6_n_0 : STD_LOGIC;
  signal W_31_3_i_7_n_0 : STD_LOGIC;
  signal W_31_3_i_8_n_0 : STD_LOGIC;
  signal W_31_3_i_9_n_0 : STD_LOGIC;
  signal W_31_7_i_10_n_0 : STD_LOGIC;
  signal W_31_7_i_11_n_0 : STD_LOGIC;
  signal W_31_7_i_12_n_0 : STD_LOGIC;
  signal W_31_7_i_13_n_0 : STD_LOGIC;
  signal W_31_7_i_14_n_0 : STD_LOGIC;
  signal W_31_7_i_15_n_0 : STD_LOGIC;
  signal W_31_7_i_16_n_0 : STD_LOGIC;
  signal W_31_7_i_17_n_0 : STD_LOGIC;
  signal W_31_7_i_2_n_0 : STD_LOGIC;
  signal W_31_7_i_3_n_0 : STD_LOGIC;
  signal W_31_7_i_4_n_0 : STD_LOGIC;
  signal W_31_7_i_5_n_0 : STD_LOGIC;
  signal W_31_7_i_6_n_0 : STD_LOGIC;
  signal W_31_7_i_7_n_0 : STD_LOGIC;
  signal W_31_7_i_8_n_0 : STD_LOGIC;
  signal W_31_7_i_9_n_0 : STD_LOGIC;
  signal W_32 : STD_LOGIC;
  signal W_32_11_i_10_n_0 : STD_LOGIC;
  signal W_32_11_i_11_n_0 : STD_LOGIC;
  signal W_32_11_i_12_n_0 : STD_LOGIC;
  signal W_32_11_i_13_n_0 : STD_LOGIC;
  signal W_32_11_i_14_n_0 : STD_LOGIC;
  signal W_32_11_i_15_n_0 : STD_LOGIC;
  signal W_32_11_i_16_n_0 : STD_LOGIC;
  signal W_32_11_i_17_n_0 : STD_LOGIC;
  signal W_32_11_i_2_n_0 : STD_LOGIC;
  signal W_32_11_i_3_n_0 : STD_LOGIC;
  signal W_32_11_i_4_n_0 : STD_LOGIC;
  signal W_32_11_i_5_n_0 : STD_LOGIC;
  signal W_32_11_i_6_n_0 : STD_LOGIC;
  signal W_32_11_i_7_n_0 : STD_LOGIC;
  signal W_32_11_i_8_n_0 : STD_LOGIC;
  signal W_32_11_i_9_n_0 : STD_LOGIC;
  signal W_32_15_i_10_n_0 : STD_LOGIC;
  signal W_32_15_i_11_n_0 : STD_LOGIC;
  signal W_32_15_i_12_n_0 : STD_LOGIC;
  signal W_32_15_i_13_n_0 : STD_LOGIC;
  signal W_32_15_i_14_n_0 : STD_LOGIC;
  signal W_32_15_i_15_n_0 : STD_LOGIC;
  signal W_32_15_i_16_n_0 : STD_LOGIC;
  signal W_32_15_i_17_n_0 : STD_LOGIC;
  signal W_32_15_i_2_n_0 : STD_LOGIC;
  signal W_32_15_i_3_n_0 : STD_LOGIC;
  signal W_32_15_i_4_n_0 : STD_LOGIC;
  signal W_32_15_i_5_n_0 : STD_LOGIC;
  signal W_32_15_i_6_n_0 : STD_LOGIC;
  signal W_32_15_i_7_n_0 : STD_LOGIC;
  signal W_32_15_i_8_n_0 : STD_LOGIC;
  signal W_32_15_i_9_n_0 : STD_LOGIC;
  signal W_32_19_i_10_n_0 : STD_LOGIC;
  signal W_32_19_i_11_n_0 : STD_LOGIC;
  signal W_32_19_i_12_n_0 : STD_LOGIC;
  signal W_32_19_i_13_n_0 : STD_LOGIC;
  signal W_32_19_i_14_n_0 : STD_LOGIC;
  signal W_32_19_i_15_n_0 : STD_LOGIC;
  signal W_32_19_i_16_n_0 : STD_LOGIC;
  signal W_32_19_i_17_n_0 : STD_LOGIC;
  signal W_32_19_i_2_n_0 : STD_LOGIC;
  signal W_32_19_i_3_n_0 : STD_LOGIC;
  signal W_32_19_i_4_n_0 : STD_LOGIC;
  signal W_32_19_i_5_n_0 : STD_LOGIC;
  signal W_32_19_i_6_n_0 : STD_LOGIC;
  signal W_32_19_i_7_n_0 : STD_LOGIC;
  signal W_32_19_i_8_n_0 : STD_LOGIC;
  signal W_32_19_i_9_n_0 : STD_LOGIC;
  signal W_32_23_i_10_n_0 : STD_LOGIC;
  signal W_32_23_i_11_n_0 : STD_LOGIC;
  signal W_32_23_i_12_n_0 : STD_LOGIC;
  signal W_32_23_i_13_n_0 : STD_LOGIC;
  signal W_32_23_i_14_n_0 : STD_LOGIC;
  signal W_32_23_i_15_n_0 : STD_LOGIC;
  signal W_32_23_i_16_n_0 : STD_LOGIC;
  signal W_32_23_i_17_n_0 : STD_LOGIC;
  signal W_32_23_i_2_n_0 : STD_LOGIC;
  signal W_32_23_i_3_n_0 : STD_LOGIC;
  signal W_32_23_i_4_n_0 : STD_LOGIC;
  signal W_32_23_i_5_n_0 : STD_LOGIC;
  signal W_32_23_i_6_n_0 : STD_LOGIC;
  signal W_32_23_i_7_n_0 : STD_LOGIC;
  signal W_32_23_i_8_n_0 : STD_LOGIC;
  signal W_32_23_i_9_n_0 : STD_LOGIC;
  signal W_32_27_i_10_n_0 : STD_LOGIC;
  signal W_32_27_i_11_n_0 : STD_LOGIC;
  signal W_32_27_i_12_n_0 : STD_LOGIC;
  signal W_32_27_i_13_n_0 : STD_LOGIC;
  signal W_32_27_i_14_n_0 : STD_LOGIC;
  signal W_32_27_i_15_n_0 : STD_LOGIC;
  signal W_32_27_i_16_n_0 : STD_LOGIC;
  signal W_32_27_i_17_n_0 : STD_LOGIC;
  signal W_32_27_i_2_n_0 : STD_LOGIC;
  signal W_32_27_i_3_n_0 : STD_LOGIC;
  signal W_32_27_i_4_n_0 : STD_LOGIC;
  signal W_32_27_i_5_n_0 : STD_LOGIC;
  signal W_32_27_i_6_n_0 : STD_LOGIC;
  signal W_32_27_i_7_n_0 : STD_LOGIC;
  signal W_32_27_i_8_n_0 : STD_LOGIC;
  signal W_32_27_i_9_n_0 : STD_LOGIC;
  signal W_32_31_i_10_n_0 : STD_LOGIC;
  signal W_32_31_i_11_n_0 : STD_LOGIC;
  signal W_32_31_i_12_n_0 : STD_LOGIC;
  signal W_32_31_i_13_n_0 : STD_LOGIC;
  signal W_32_31_i_14_n_0 : STD_LOGIC;
  signal W_32_31_i_15_n_0 : STD_LOGIC;
  signal W_32_31_i_16_n_0 : STD_LOGIC;
  signal W_32_31_i_18_n_0 : STD_LOGIC;
  signal W_32_31_i_20_n_0 : STD_LOGIC;
  signal W_32_31_i_3_n_0 : STD_LOGIC;
  signal W_32_31_i_4_n_0 : STD_LOGIC;
  signal W_32_31_i_5_n_0 : STD_LOGIC;
  signal W_32_31_i_6_n_0 : STD_LOGIC;
  signal W_32_31_i_7_n_0 : STD_LOGIC;
  signal W_32_31_i_8_n_0 : STD_LOGIC;
  signal W_32_31_i_9_n_0 : STD_LOGIC;
  signal W_32_3_i_10_n_0 : STD_LOGIC;
  signal W_32_3_i_11_n_0 : STD_LOGIC;
  signal W_32_3_i_15_n_0 : STD_LOGIC;
  signal W_32_3_i_2_n_0 : STD_LOGIC;
  signal W_32_3_i_3_n_0 : STD_LOGIC;
  signal W_32_3_i_4_n_0 : STD_LOGIC;
  signal W_32_3_i_5_n_0 : STD_LOGIC;
  signal W_32_3_i_6_n_0 : STD_LOGIC;
  signal W_32_3_i_7_n_0 : STD_LOGIC;
  signal W_32_3_i_8_n_0 : STD_LOGIC;
  signal W_32_3_i_9_n_0 : STD_LOGIC;
  signal W_32_7_i_10_n_0 : STD_LOGIC;
  signal W_32_7_i_11_n_0 : STD_LOGIC;
  signal W_32_7_i_12_n_0 : STD_LOGIC;
  signal W_32_7_i_13_n_0 : STD_LOGIC;
  signal W_32_7_i_14_n_0 : STD_LOGIC;
  signal W_32_7_i_15_n_0 : STD_LOGIC;
  signal W_32_7_i_16_n_0 : STD_LOGIC;
  signal W_32_7_i_17_n_0 : STD_LOGIC;
  signal W_32_7_i_2_n_0 : STD_LOGIC;
  signal W_32_7_i_3_n_0 : STD_LOGIC;
  signal W_32_7_i_4_n_0 : STD_LOGIC;
  signal W_32_7_i_5_n_0 : STD_LOGIC;
  signal W_32_7_i_6_n_0 : STD_LOGIC;
  signal W_32_7_i_7_n_0 : STD_LOGIC;
  signal W_32_7_i_8_n_0 : STD_LOGIC;
  signal W_32_7_i_9_n_0 : STD_LOGIC;
  signal W_33_11_i_10_n_0 : STD_LOGIC;
  signal W_33_11_i_11_n_0 : STD_LOGIC;
  signal W_33_11_i_12_n_0 : STD_LOGIC;
  signal W_33_11_i_13_n_0 : STD_LOGIC;
  signal W_33_11_i_14_n_0 : STD_LOGIC;
  signal W_33_11_i_15_n_0 : STD_LOGIC;
  signal W_33_11_i_16_n_0 : STD_LOGIC;
  signal W_33_11_i_17_n_0 : STD_LOGIC;
  signal W_33_11_i_2_n_0 : STD_LOGIC;
  signal W_33_11_i_3_n_0 : STD_LOGIC;
  signal W_33_11_i_4_n_0 : STD_LOGIC;
  signal W_33_11_i_5_n_0 : STD_LOGIC;
  signal W_33_11_i_6_n_0 : STD_LOGIC;
  signal W_33_11_i_7_n_0 : STD_LOGIC;
  signal W_33_11_i_8_n_0 : STD_LOGIC;
  signal W_33_11_i_9_n_0 : STD_LOGIC;
  signal W_33_15_i_10_n_0 : STD_LOGIC;
  signal W_33_15_i_11_n_0 : STD_LOGIC;
  signal W_33_15_i_12_n_0 : STD_LOGIC;
  signal W_33_15_i_13_n_0 : STD_LOGIC;
  signal W_33_15_i_14_n_0 : STD_LOGIC;
  signal W_33_15_i_15_n_0 : STD_LOGIC;
  signal W_33_15_i_16_n_0 : STD_LOGIC;
  signal W_33_15_i_17_n_0 : STD_LOGIC;
  signal W_33_15_i_2_n_0 : STD_LOGIC;
  signal W_33_15_i_3_n_0 : STD_LOGIC;
  signal W_33_15_i_4_n_0 : STD_LOGIC;
  signal W_33_15_i_5_n_0 : STD_LOGIC;
  signal W_33_15_i_6_n_0 : STD_LOGIC;
  signal W_33_15_i_7_n_0 : STD_LOGIC;
  signal W_33_15_i_8_n_0 : STD_LOGIC;
  signal W_33_15_i_9_n_0 : STD_LOGIC;
  signal W_33_19_i_10_n_0 : STD_LOGIC;
  signal W_33_19_i_11_n_0 : STD_LOGIC;
  signal W_33_19_i_12_n_0 : STD_LOGIC;
  signal W_33_19_i_13_n_0 : STD_LOGIC;
  signal W_33_19_i_14_n_0 : STD_LOGIC;
  signal W_33_19_i_15_n_0 : STD_LOGIC;
  signal W_33_19_i_16_n_0 : STD_LOGIC;
  signal W_33_19_i_17_n_0 : STD_LOGIC;
  signal W_33_19_i_2_n_0 : STD_LOGIC;
  signal W_33_19_i_3_n_0 : STD_LOGIC;
  signal W_33_19_i_4_n_0 : STD_LOGIC;
  signal W_33_19_i_5_n_0 : STD_LOGIC;
  signal W_33_19_i_6_n_0 : STD_LOGIC;
  signal W_33_19_i_7_n_0 : STD_LOGIC;
  signal W_33_19_i_8_n_0 : STD_LOGIC;
  signal W_33_19_i_9_n_0 : STD_LOGIC;
  signal W_33_23_i_10_n_0 : STD_LOGIC;
  signal W_33_23_i_11_n_0 : STD_LOGIC;
  signal W_33_23_i_12_n_0 : STD_LOGIC;
  signal W_33_23_i_13_n_0 : STD_LOGIC;
  signal W_33_23_i_14_n_0 : STD_LOGIC;
  signal W_33_23_i_15_n_0 : STD_LOGIC;
  signal W_33_23_i_16_n_0 : STD_LOGIC;
  signal W_33_23_i_17_n_0 : STD_LOGIC;
  signal W_33_23_i_2_n_0 : STD_LOGIC;
  signal W_33_23_i_3_n_0 : STD_LOGIC;
  signal W_33_23_i_4_n_0 : STD_LOGIC;
  signal W_33_23_i_5_n_0 : STD_LOGIC;
  signal W_33_23_i_6_n_0 : STD_LOGIC;
  signal W_33_23_i_7_n_0 : STD_LOGIC;
  signal W_33_23_i_8_n_0 : STD_LOGIC;
  signal W_33_23_i_9_n_0 : STD_LOGIC;
  signal W_33_27_i_10_n_0 : STD_LOGIC;
  signal W_33_27_i_11_n_0 : STD_LOGIC;
  signal W_33_27_i_12_n_0 : STD_LOGIC;
  signal W_33_27_i_13_n_0 : STD_LOGIC;
  signal W_33_27_i_14_n_0 : STD_LOGIC;
  signal W_33_27_i_15_n_0 : STD_LOGIC;
  signal W_33_27_i_16_n_0 : STD_LOGIC;
  signal W_33_27_i_17_n_0 : STD_LOGIC;
  signal W_33_27_i_2_n_0 : STD_LOGIC;
  signal W_33_27_i_3_n_0 : STD_LOGIC;
  signal W_33_27_i_4_n_0 : STD_LOGIC;
  signal W_33_27_i_5_n_0 : STD_LOGIC;
  signal W_33_27_i_6_n_0 : STD_LOGIC;
  signal W_33_27_i_7_n_0 : STD_LOGIC;
  signal W_33_27_i_8_n_0 : STD_LOGIC;
  signal W_33_27_i_9_n_0 : STD_LOGIC;
  signal W_33_31_i_10_n_0 : STD_LOGIC;
  signal W_33_31_i_11_n_0 : STD_LOGIC;
  signal W_33_31_i_12_n_0 : STD_LOGIC;
  signal W_33_31_i_13_n_0 : STD_LOGIC;
  signal W_33_31_i_14_n_0 : STD_LOGIC;
  signal W_33_31_i_15_n_0 : STD_LOGIC;
  signal W_33_31_i_17_n_0 : STD_LOGIC;
  signal W_33_31_i_19_n_0 : STD_LOGIC;
  signal W_33_31_i_2_n_0 : STD_LOGIC;
  signal W_33_31_i_3_n_0 : STD_LOGIC;
  signal W_33_31_i_4_n_0 : STD_LOGIC;
  signal W_33_31_i_5_n_0 : STD_LOGIC;
  signal W_33_31_i_6_n_0 : STD_LOGIC;
  signal W_33_31_i_7_n_0 : STD_LOGIC;
  signal W_33_31_i_8_n_0 : STD_LOGIC;
  signal W_33_31_i_9_n_0 : STD_LOGIC;
  signal W_33_3_i_10_n_0 : STD_LOGIC;
  signal W_33_3_i_11_n_0 : STD_LOGIC;
  signal W_33_3_i_15_n_0 : STD_LOGIC;
  signal W_33_3_i_2_n_0 : STD_LOGIC;
  signal W_33_3_i_3_n_0 : STD_LOGIC;
  signal W_33_3_i_4_n_0 : STD_LOGIC;
  signal W_33_3_i_5_n_0 : STD_LOGIC;
  signal W_33_3_i_6_n_0 : STD_LOGIC;
  signal W_33_3_i_7_n_0 : STD_LOGIC;
  signal W_33_3_i_8_n_0 : STD_LOGIC;
  signal W_33_3_i_9_n_0 : STD_LOGIC;
  signal W_33_7_i_10_n_0 : STD_LOGIC;
  signal W_33_7_i_11_n_0 : STD_LOGIC;
  signal W_33_7_i_12_n_0 : STD_LOGIC;
  signal W_33_7_i_13_n_0 : STD_LOGIC;
  signal W_33_7_i_14_n_0 : STD_LOGIC;
  signal W_33_7_i_15_n_0 : STD_LOGIC;
  signal W_33_7_i_16_n_0 : STD_LOGIC;
  signal W_33_7_i_17_n_0 : STD_LOGIC;
  signal W_33_7_i_2_n_0 : STD_LOGIC;
  signal W_33_7_i_3_n_0 : STD_LOGIC;
  signal W_33_7_i_4_n_0 : STD_LOGIC;
  signal W_33_7_i_5_n_0 : STD_LOGIC;
  signal W_33_7_i_6_n_0 : STD_LOGIC;
  signal W_33_7_i_7_n_0 : STD_LOGIC;
  signal W_33_7_i_8_n_0 : STD_LOGIC;
  signal W_33_7_i_9_n_0 : STD_LOGIC;
  signal W_34_11_i_10_n_0 : STD_LOGIC;
  signal W_34_11_i_11_n_0 : STD_LOGIC;
  signal W_34_11_i_12_n_0 : STD_LOGIC;
  signal W_34_11_i_13_n_0 : STD_LOGIC;
  signal W_34_11_i_14_n_0 : STD_LOGIC;
  signal W_34_11_i_15_n_0 : STD_LOGIC;
  signal W_34_11_i_16_n_0 : STD_LOGIC;
  signal W_34_11_i_17_n_0 : STD_LOGIC;
  signal W_34_11_i_2_n_0 : STD_LOGIC;
  signal W_34_11_i_3_n_0 : STD_LOGIC;
  signal W_34_11_i_4_n_0 : STD_LOGIC;
  signal W_34_11_i_5_n_0 : STD_LOGIC;
  signal W_34_11_i_6_n_0 : STD_LOGIC;
  signal W_34_11_i_7_n_0 : STD_LOGIC;
  signal W_34_11_i_8_n_0 : STD_LOGIC;
  signal W_34_11_i_9_n_0 : STD_LOGIC;
  signal W_34_15_i_10_n_0 : STD_LOGIC;
  signal W_34_15_i_11_n_0 : STD_LOGIC;
  signal W_34_15_i_12_n_0 : STD_LOGIC;
  signal W_34_15_i_13_n_0 : STD_LOGIC;
  signal W_34_15_i_14_n_0 : STD_LOGIC;
  signal W_34_15_i_15_n_0 : STD_LOGIC;
  signal W_34_15_i_16_n_0 : STD_LOGIC;
  signal W_34_15_i_17_n_0 : STD_LOGIC;
  signal W_34_15_i_2_n_0 : STD_LOGIC;
  signal W_34_15_i_3_n_0 : STD_LOGIC;
  signal W_34_15_i_4_n_0 : STD_LOGIC;
  signal W_34_15_i_5_n_0 : STD_LOGIC;
  signal W_34_15_i_6_n_0 : STD_LOGIC;
  signal W_34_15_i_7_n_0 : STD_LOGIC;
  signal W_34_15_i_8_n_0 : STD_LOGIC;
  signal W_34_15_i_9_n_0 : STD_LOGIC;
  signal W_34_19_i_10_n_0 : STD_LOGIC;
  signal W_34_19_i_11_n_0 : STD_LOGIC;
  signal W_34_19_i_12_n_0 : STD_LOGIC;
  signal W_34_19_i_13_n_0 : STD_LOGIC;
  signal W_34_19_i_14_n_0 : STD_LOGIC;
  signal W_34_19_i_15_n_0 : STD_LOGIC;
  signal W_34_19_i_16_n_0 : STD_LOGIC;
  signal W_34_19_i_17_n_0 : STD_LOGIC;
  signal W_34_19_i_2_n_0 : STD_LOGIC;
  signal W_34_19_i_3_n_0 : STD_LOGIC;
  signal W_34_19_i_4_n_0 : STD_LOGIC;
  signal W_34_19_i_5_n_0 : STD_LOGIC;
  signal W_34_19_i_6_n_0 : STD_LOGIC;
  signal W_34_19_i_7_n_0 : STD_LOGIC;
  signal W_34_19_i_8_n_0 : STD_LOGIC;
  signal W_34_19_i_9_n_0 : STD_LOGIC;
  signal W_34_23_i_10_n_0 : STD_LOGIC;
  signal W_34_23_i_11_n_0 : STD_LOGIC;
  signal W_34_23_i_12_n_0 : STD_LOGIC;
  signal W_34_23_i_13_n_0 : STD_LOGIC;
  signal W_34_23_i_14_n_0 : STD_LOGIC;
  signal W_34_23_i_15_n_0 : STD_LOGIC;
  signal W_34_23_i_16_n_0 : STD_LOGIC;
  signal W_34_23_i_17_n_0 : STD_LOGIC;
  signal W_34_23_i_2_n_0 : STD_LOGIC;
  signal W_34_23_i_3_n_0 : STD_LOGIC;
  signal W_34_23_i_4_n_0 : STD_LOGIC;
  signal W_34_23_i_5_n_0 : STD_LOGIC;
  signal W_34_23_i_6_n_0 : STD_LOGIC;
  signal W_34_23_i_7_n_0 : STD_LOGIC;
  signal W_34_23_i_8_n_0 : STD_LOGIC;
  signal W_34_23_i_9_n_0 : STD_LOGIC;
  signal W_34_27_i_10_n_0 : STD_LOGIC;
  signal W_34_27_i_11_n_0 : STD_LOGIC;
  signal W_34_27_i_12_n_0 : STD_LOGIC;
  signal W_34_27_i_13_n_0 : STD_LOGIC;
  signal W_34_27_i_14_n_0 : STD_LOGIC;
  signal W_34_27_i_15_n_0 : STD_LOGIC;
  signal W_34_27_i_16_n_0 : STD_LOGIC;
  signal W_34_27_i_17_n_0 : STD_LOGIC;
  signal W_34_27_i_2_n_0 : STD_LOGIC;
  signal W_34_27_i_3_n_0 : STD_LOGIC;
  signal W_34_27_i_4_n_0 : STD_LOGIC;
  signal W_34_27_i_5_n_0 : STD_LOGIC;
  signal W_34_27_i_6_n_0 : STD_LOGIC;
  signal W_34_27_i_7_n_0 : STD_LOGIC;
  signal W_34_27_i_8_n_0 : STD_LOGIC;
  signal W_34_27_i_9_n_0 : STD_LOGIC;
  signal W_34_31_i_10_n_0 : STD_LOGIC;
  signal W_34_31_i_11_n_0 : STD_LOGIC;
  signal W_34_31_i_12_n_0 : STD_LOGIC;
  signal W_34_31_i_13_n_0 : STD_LOGIC;
  signal W_34_31_i_14_n_0 : STD_LOGIC;
  signal W_34_31_i_15_n_0 : STD_LOGIC;
  signal W_34_31_i_17_n_0 : STD_LOGIC;
  signal W_34_31_i_19_n_0 : STD_LOGIC;
  signal W_34_31_i_2_n_0 : STD_LOGIC;
  signal W_34_31_i_3_n_0 : STD_LOGIC;
  signal W_34_31_i_4_n_0 : STD_LOGIC;
  signal W_34_31_i_5_n_0 : STD_LOGIC;
  signal W_34_31_i_6_n_0 : STD_LOGIC;
  signal W_34_31_i_7_n_0 : STD_LOGIC;
  signal W_34_31_i_8_n_0 : STD_LOGIC;
  signal W_34_31_i_9_n_0 : STD_LOGIC;
  signal W_34_3_i_10_n_0 : STD_LOGIC;
  signal W_34_3_i_11_n_0 : STD_LOGIC;
  signal W_34_3_i_15_n_0 : STD_LOGIC;
  signal W_34_3_i_2_n_0 : STD_LOGIC;
  signal W_34_3_i_3_n_0 : STD_LOGIC;
  signal W_34_3_i_4_n_0 : STD_LOGIC;
  signal W_34_3_i_5_n_0 : STD_LOGIC;
  signal W_34_3_i_6_n_0 : STD_LOGIC;
  signal W_34_3_i_7_n_0 : STD_LOGIC;
  signal W_34_3_i_8_n_0 : STD_LOGIC;
  signal W_34_3_i_9_n_0 : STD_LOGIC;
  signal W_34_7_i_10_n_0 : STD_LOGIC;
  signal W_34_7_i_11_n_0 : STD_LOGIC;
  signal W_34_7_i_12_n_0 : STD_LOGIC;
  signal W_34_7_i_13_n_0 : STD_LOGIC;
  signal W_34_7_i_14_n_0 : STD_LOGIC;
  signal W_34_7_i_15_n_0 : STD_LOGIC;
  signal W_34_7_i_16_n_0 : STD_LOGIC;
  signal W_34_7_i_17_n_0 : STD_LOGIC;
  signal W_34_7_i_2_n_0 : STD_LOGIC;
  signal W_34_7_i_3_n_0 : STD_LOGIC;
  signal W_34_7_i_4_n_0 : STD_LOGIC;
  signal W_34_7_i_5_n_0 : STD_LOGIC;
  signal W_34_7_i_6_n_0 : STD_LOGIC;
  signal W_34_7_i_7_n_0 : STD_LOGIC;
  signal W_34_7_i_8_n_0 : STD_LOGIC;
  signal W_34_7_i_9_n_0 : STD_LOGIC;
  signal W_35_11_i_10_n_0 : STD_LOGIC;
  signal W_35_11_i_11_n_0 : STD_LOGIC;
  signal W_35_11_i_12_n_0 : STD_LOGIC;
  signal W_35_11_i_13_n_0 : STD_LOGIC;
  signal W_35_11_i_14_n_0 : STD_LOGIC;
  signal W_35_11_i_15_n_0 : STD_LOGIC;
  signal W_35_11_i_16_n_0 : STD_LOGIC;
  signal W_35_11_i_17_n_0 : STD_LOGIC;
  signal W_35_11_i_2_n_0 : STD_LOGIC;
  signal W_35_11_i_3_n_0 : STD_LOGIC;
  signal W_35_11_i_4_n_0 : STD_LOGIC;
  signal W_35_11_i_5_n_0 : STD_LOGIC;
  signal W_35_11_i_6_n_0 : STD_LOGIC;
  signal W_35_11_i_7_n_0 : STD_LOGIC;
  signal W_35_11_i_8_n_0 : STD_LOGIC;
  signal W_35_11_i_9_n_0 : STD_LOGIC;
  signal W_35_15_i_10_n_0 : STD_LOGIC;
  signal W_35_15_i_11_n_0 : STD_LOGIC;
  signal W_35_15_i_12_n_0 : STD_LOGIC;
  signal W_35_15_i_13_n_0 : STD_LOGIC;
  signal W_35_15_i_14_n_0 : STD_LOGIC;
  signal W_35_15_i_15_n_0 : STD_LOGIC;
  signal W_35_15_i_16_n_0 : STD_LOGIC;
  signal W_35_15_i_17_n_0 : STD_LOGIC;
  signal W_35_15_i_2_n_0 : STD_LOGIC;
  signal W_35_15_i_3_n_0 : STD_LOGIC;
  signal W_35_15_i_4_n_0 : STD_LOGIC;
  signal W_35_15_i_5_n_0 : STD_LOGIC;
  signal W_35_15_i_6_n_0 : STD_LOGIC;
  signal W_35_15_i_7_n_0 : STD_LOGIC;
  signal W_35_15_i_8_n_0 : STD_LOGIC;
  signal W_35_15_i_9_n_0 : STD_LOGIC;
  signal W_35_19_i_10_n_0 : STD_LOGIC;
  signal W_35_19_i_11_n_0 : STD_LOGIC;
  signal W_35_19_i_12_n_0 : STD_LOGIC;
  signal W_35_19_i_13_n_0 : STD_LOGIC;
  signal W_35_19_i_14_n_0 : STD_LOGIC;
  signal W_35_19_i_15_n_0 : STD_LOGIC;
  signal W_35_19_i_16_n_0 : STD_LOGIC;
  signal W_35_19_i_17_n_0 : STD_LOGIC;
  signal W_35_19_i_2_n_0 : STD_LOGIC;
  signal W_35_19_i_3_n_0 : STD_LOGIC;
  signal W_35_19_i_4_n_0 : STD_LOGIC;
  signal W_35_19_i_5_n_0 : STD_LOGIC;
  signal W_35_19_i_6_n_0 : STD_LOGIC;
  signal W_35_19_i_7_n_0 : STD_LOGIC;
  signal W_35_19_i_8_n_0 : STD_LOGIC;
  signal W_35_19_i_9_n_0 : STD_LOGIC;
  signal W_35_23_i_10_n_0 : STD_LOGIC;
  signal W_35_23_i_11_n_0 : STD_LOGIC;
  signal W_35_23_i_12_n_0 : STD_LOGIC;
  signal W_35_23_i_13_n_0 : STD_LOGIC;
  signal W_35_23_i_14_n_0 : STD_LOGIC;
  signal W_35_23_i_15_n_0 : STD_LOGIC;
  signal W_35_23_i_16_n_0 : STD_LOGIC;
  signal W_35_23_i_17_n_0 : STD_LOGIC;
  signal W_35_23_i_2_n_0 : STD_LOGIC;
  signal W_35_23_i_3_n_0 : STD_LOGIC;
  signal W_35_23_i_4_n_0 : STD_LOGIC;
  signal W_35_23_i_5_n_0 : STD_LOGIC;
  signal W_35_23_i_6_n_0 : STD_LOGIC;
  signal W_35_23_i_7_n_0 : STD_LOGIC;
  signal W_35_23_i_8_n_0 : STD_LOGIC;
  signal W_35_23_i_9_n_0 : STD_LOGIC;
  signal W_35_27_i_10_n_0 : STD_LOGIC;
  signal W_35_27_i_11_n_0 : STD_LOGIC;
  signal W_35_27_i_12_n_0 : STD_LOGIC;
  signal W_35_27_i_13_n_0 : STD_LOGIC;
  signal W_35_27_i_14_n_0 : STD_LOGIC;
  signal W_35_27_i_15_n_0 : STD_LOGIC;
  signal W_35_27_i_16_n_0 : STD_LOGIC;
  signal W_35_27_i_17_n_0 : STD_LOGIC;
  signal W_35_27_i_2_n_0 : STD_LOGIC;
  signal W_35_27_i_3_n_0 : STD_LOGIC;
  signal W_35_27_i_4_n_0 : STD_LOGIC;
  signal W_35_27_i_5_n_0 : STD_LOGIC;
  signal W_35_27_i_6_n_0 : STD_LOGIC;
  signal W_35_27_i_7_n_0 : STD_LOGIC;
  signal W_35_27_i_8_n_0 : STD_LOGIC;
  signal W_35_27_i_9_n_0 : STD_LOGIC;
  signal W_35_31_i_10_n_0 : STD_LOGIC;
  signal W_35_31_i_11_n_0 : STD_LOGIC;
  signal W_35_31_i_12_n_0 : STD_LOGIC;
  signal W_35_31_i_13_n_0 : STD_LOGIC;
  signal W_35_31_i_14_n_0 : STD_LOGIC;
  signal W_35_31_i_15_n_0 : STD_LOGIC;
  signal W_35_31_i_17_n_0 : STD_LOGIC;
  signal W_35_31_i_19_n_0 : STD_LOGIC;
  signal W_35_31_i_2_n_0 : STD_LOGIC;
  signal W_35_31_i_3_n_0 : STD_LOGIC;
  signal W_35_31_i_4_n_0 : STD_LOGIC;
  signal W_35_31_i_5_n_0 : STD_LOGIC;
  signal W_35_31_i_6_n_0 : STD_LOGIC;
  signal W_35_31_i_7_n_0 : STD_LOGIC;
  signal W_35_31_i_8_n_0 : STD_LOGIC;
  signal W_35_31_i_9_n_0 : STD_LOGIC;
  signal W_35_3_i_10_n_0 : STD_LOGIC;
  signal W_35_3_i_11_n_0 : STD_LOGIC;
  signal W_35_3_i_15_n_0 : STD_LOGIC;
  signal W_35_3_i_2_n_0 : STD_LOGIC;
  signal W_35_3_i_3_n_0 : STD_LOGIC;
  signal W_35_3_i_4_n_0 : STD_LOGIC;
  signal W_35_3_i_5_n_0 : STD_LOGIC;
  signal W_35_3_i_6_n_0 : STD_LOGIC;
  signal W_35_3_i_7_n_0 : STD_LOGIC;
  signal W_35_3_i_8_n_0 : STD_LOGIC;
  signal W_35_3_i_9_n_0 : STD_LOGIC;
  signal W_35_7_i_10_n_0 : STD_LOGIC;
  signal W_35_7_i_11_n_0 : STD_LOGIC;
  signal W_35_7_i_12_n_0 : STD_LOGIC;
  signal W_35_7_i_13_n_0 : STD_LOGIC;
  signal W_35_7_i_14_n_0 : STD_LOGIC;
  signal W_35_7_i_15_n_0 : STD_LOGIC;
  signal W_35_7_i_16_n_0 : STD_LOGIC;
  signal W_35_7_i_17_n_0 : STD_LOGIC;
  signal W_35_7_i_2_n_0 : STD_LOGIC;
  signal W_35_7_i_3_n_0 : STD_LOGIC;
  signal W_35_7_i_4_n_0 : STD_LOGIC;
  signal W_35_7_i_5_n_0 : STD_LOGIC;
  signal W_35_7_i_6_n_0 : STD_LOGIC;
  signal W_35_7_i_7_n_0 : STD_LOGIC;
  signal W_35_7_i_8_n_0 : STD_LOGIC;
  signal W_35_7_i_9_n_0 : STD_LOGIC;
  signal W_36_11_i_10_n_0 : STD_LOGIC;
  signal W_36_11_i_11_n_0 : STD_LOGIC;
  signal W_36_11_i_12_n_0 : STD_LOGIC;
  signal W_36_11_i_13_n_0 : STD_LOGIC;
  signal W_36_11_i_14_n_0 : STD_LOGIC;
  signal W_36_11_i_15_n_0 : STD_LOGIC;
  signal W_36_11_i_16_n_0 : STD_LOGIC;
  signal W_36_11_i_17_n_0 : STD_LOGIC;
  signal W_36_11_i_2_n_0 : STD_LOGIC;
  signal W_36_11_i_3_n_0 : STD_LOGIC;
  signal W_36_11_i_4_n_0 : STD_LOGIC;
  signal W_36_11_i_5_n_0 : STD_LOGIC;
  signal W_36_11_i_6_n_0 : STD_LOGIC;
  signal W_36_11_i_7_n_0 : STD_LOGIC;
  signal W_36_11_i_8_n_0 : STD_LOGIC;
  signal W_36_11_i_9_n_0 : STD_LOGIC;
  signal W_36_15_i_10_n_0 : STD_LOGIC;
  signal W_36_15_i_11_n_0 : STD_LOGIC;
  signal W_36_15_i_12_n_0 : STD_LOGIC;
  signal W_36_15_i_13_n_0 : STD_LOGIC;
  signal W_36_15_i_14_n_0 : STD_LOGIC;
  signal W_36_15_i_15_n_0 : STD_LOGIC;
  signal W_36_15_i_16_n_0 : STD_LOGIC;
  signal W_36_15_i_17_n_0 : STD_LOGIC;
  signal W_36_15_i_2_n_0 : STD_LOGIC;
  signal W_36_15_i_3_n_0 : STD_LOGIC;
  signal W_36_15_i_4_n_0 : STD_LOGIC;
  signal W_36_15_i_5_n_0 : STD_LOGIC;
  signal W_36_15_i_6_n_0 : STD_LOGIC;
  signal W_36_15_i_7_n_0 : STD_LOGIC;
  signal W_36_15_i_8_n_0 : STD_LOGIC;
  signal W_36_15_i_9_n_0 : STD_LOGIC;
  signal W_36_19_i_10_n_0 : STD_LOGIC;
  signal W_36_19_i_11_n_0 : STD_LOGIC;
  signal W_36_19_i_12_n_0 : STD_LOGIC;
  signal W_36_19_i_13_n_0 : STD_LOGIC;
  signal W_36_19_i_14_n_0 : STD_LOGIC;
  signal W_36_19_i_15_n_0 : STD_LOGIC;
  signal W_36_19_i_16_n_0 : STD_LOGIC;
  signal W_36_19_i_17_n_0 : STD_LOGIC;
  signal W_36_19_i_2_n_0 : STD_LOGIC;
  signal W_36_19_i_3_n_0 : STD_LOGIC;
  signal W_36_19_i_4_n_0 : STD_LOGIC;
  signal W_36_19_i_5_n_0 : STD_LOGIC;
  signal W_36_19_i_6_n_0 : STD_LOGIC;
  signal W_36_19_i_7_n_0 : STD_LOGIC;
  signal W_36_19_i_8_n_0 : STD_LOGIC;
  signal W_36_19_i_9_n_0 : STD_LOGIC;
  signal W_36_23_i_10_n_0 : STD_LOGIC;
  signal W_36_23_i_11_n_0 : STD_LOGIC;
  signal W_36_23_i_12_n_0 : STD_LOGIC;
  signal W_36_23_i_13_n_0 : STD_LOGIC;
  signal W_36_23_i_14_n_0 : STD_LOGIC;
  signal W_36_23_i_15_n_0 : STD_LOGIC;
  signal W_36_23_i_16_n_0 : STD_LOGIC;
  signal W_36_23_i_17_n_0 : STD_LOGIC;
  signal W_36_23_i_2_n_0 : STD_LOGIC;
  signal W_36_23_i_3_n_0 : STD_LOGIC;
  signal W_36_23_i_4_n_0 : STD_LOGIC;
  signal W_36_23_i_5_n_0 : STD_LOGIC;
  signal W_36_23_i_6_n_0 : STD_LOGIC;
  signal W_36_23_i_7_n_0 : STD_LOGIC;
  signal W_36_23_i_8_n_0 : STD_LOGIC;
  signal W_36_23_i_9_n_0 : STD_LOGIC;
  signal W_36_27_i_10_n_0 : STD_LOGIC;
  signal W_36_27_i_11_n_0 : STD_LOGIC;
  signal W_36_27_i_12_n_0 : STD_LOGIC;
  signal W_36_27_i_13_n_0 : STD_LOGIC;
  signal W_36_27_i_14_n_0 : STD_LOGIC;
  signal W_36_27_i_15_n_0 : STD_LOGIC;
  signal W_36_27_i_16_n_0 : STD_LOGIC;
  signal W_36_27_i_17_n_0 : STD_LOGIC;
  signal W_36_27_i_2_n_0 : STD_LOGIC;
  signal W_36_27_i_3_n_0 : STD_LOGIC;
  signal W_36_27_i_4_n_0 : STD_LOGIC;
  signal W_36_27_i_5_n_0 : STD_LOGIC;
  signal W_36_27_i_6_n_0 : STD_LOGIC;
  signal W_36_27_i_7_n_0 : STD_LOGIC;
  signal W_36_27_i_8_n_0 : STD_LOGIC;
  signal W_36_27_i_9_n_0 : STD_LOGIC;
  signal W_36_31_i_10_n_0 : STD_LOGIC;
  signal W_36_31_i_11_n_0 : STD_LOGIC;
  signal W_36_31_i_12_n_0 : STD_LOGIC;
  signal W_36_31_i_13_n_0 : STD_LOGIC;
  signal W_36_31_i_14_n_0 : STD_LOGIC;
  signal W_36_31_i_15_n_0 : STD_LOGIC;
  signal W_36_31_i_17_n_0 : STD_LOGIC;
  signal W_36_31_i_19_n_0 : STD_LOGIC;
  signal W_36_31_i_2_n_0 : STD_LOGIC;
  signal W_36_31_i_3_n_0 : STD_LOGIC;
  signal W_36_31_i_4_n_0 : STD_LOGIC;
  signal W_36_31_i_5_n_0 : STD_LOGIC;
  signal W_36_31_i_6_n_0 : STD_LOGIC;
  signal W_36_31_i_7_n_0 : STD_LOGIC;
  signal W_36_31_i_8_n_0 : STD_LOGIC;
  signal W_36_31_i_9_n_0 : STD_LOGIC;
  signal W_36_3_i_10_n_0 : STD_LOGIC;
  signal W_36_3_i_11_n_0 : STD_LOGIC;
  signal W_36_3_i_15_n_0 : STD_LOGIC;
  signal W_36_3_i_2_n_0 : STD_LOGIC;
  signal W_36_3_i_3_n_0 : STD_LOGIC;
  signal W_36_3_i_4_n_0 : STD_LOGIC;
  signal W_36_3_i_5_n_0 : STD_LOGIC;
  signal W_36_3_i_6_n_0 : STD_LOGIC;
  signal W_36_3_i_7_n_0 : STD_LOGIC;
  signal W_36_3_i_8_n_0 : STD_LOGIC;
  signal W_36_3_i_9_n_0 : STD_LOGIC;
  signal W_36_7_i_10_n_0 : STD_LOGIC;
  signal W_36_7_i_11_n_0 : STD_LOGIC;
  signal W_36_7_i_12_n_0 : STD_LOGIC;
  signal W_36_7_i_13_n_0 : STD_LOGIC;
  signal W_36_7_i_14_n_0 : STD_LOGIC;
  signal W_36_7_i_15_n_0 : STD_LOGIC;
  signal W_36_7_i_16_n_0 : STD_LOGIC;
  signal W_36_7_i_17_n_0 : STD_LOGIC;
  signal W_36_7_i_2_n_0 : STD_LOGIC;
  signal W_36_7_i_3_n_0 : STD_LOGIC;
  signal W_36_7_i_4_n_0 : STD_LOGIC;
  signal W_36_7_i_5_n_0 : STD_LOGIC;
  signal W_36_7_i_6_n_0 : STD_LOGIC;
  signal W_36_7_i_7_n_0 : STD_LOGIC;
  signal W_36_7_i_8_n_0 : STD_LOGIC;
  signal W_36_7_i_9_n_0 : STD_LOGIC;
  signal W_37_11_i_10_n_0 : STD_LOGIC;
  signal W_37_11_i_11_n_0 : STD_LOGIC;
  signal W_37_11_i_12_n_0 : STD_LOGIC;
  signal W_37_11_i_13_n_0 : STD_LOGIC;
  signal W_37_11_i_14_n_0 : STD_LOGIC;
  signal W_37_11_i_15_n_0 : STD_LOGIC;
  signal W_37_11_i_16_n_0 : STD_LOGIC;
  signal W_37_11_i_17_n_0 : STD_LOGIC;
  signal W_37_11_i_2_n_0 : STD_LOGIC;
  signal W_37_11_i_3_n_0 : STD_LOGIC;
  signal W_37_11_i_4_n_0 : STD_LOGIC;
  signal W_37_11_i_5_n_0 : STD_LOGIC;
  signal W_37_11_i_6_n_0 : STD_LOGIC;
  signal W_37_11_i_7_n_0 : STD_LOGIC;
  signal W_37_11_i_8_n_0 : STD_LOGIC;
  signal W_37_11_i_9_n_0 : STD_LOGIC;
  signal W_37_15_i_10_n_0 : STD_LOGIC;
  signal W_37_15_i_11_n_0 : STD_LOGIC;
  signal W_37_15_i_12_n_0 : STD_LOGIC;
  signal W_37_15_i_13_n_0 : STD_LOGIC;
  signal W_37_15_i_14_n_0 : STD_LOGIC;
  signal W_37_15_i_15_n_0 : STD_LOGIC;
  signal W_37_15_i_16_n_0 : STD_LOGIC;
  signal W_37_15_i_17_n_0 : STD_LOGIC;
  signal W_37_15_i_2_n_0 : STD_LOGIC;
  signal W_37_15_i_3_n_0 : STD_LOGIC;
  signal W_37_15_i_4_n_0 : STD_LOGIC;
  signal W_37_15_i_5_n_0 : STD_LOGIC;
  signal W_37_15_i_6_n_0 : STD_LOGIC;
  signal W_37_15_i_7_n_0 : STD_LOGIC;
  signal W_37_15_i_8_n_0 : STD_LOGIC;
  signal W_37_15_i_9_n_0 : STD_LOGIC;
  signal W_37_19_i_10_n_0 : STD_LOGIC;
  signal W_37_19_i_11_n_0 : STD_LOGIC;
  signal W_37_19_i_12_n_0 : STD_LOGIC;
  signal W_37_19_i_13_n_0 : STD_LOGIC;
  signal W_37_19_i_14_n_0 : STD_LOGIC;
  signal W_37_19_i_15_n_0 : STD_LOGIC;
  signal W_37_19_i_16_n_0 : STD_LOGIC;
  signal W_37_19_i_17_n_0 : STD_LOGIC;
  signal W_37_19_i_2_n_0 : STD_LOGIC;
  signal W_37_19_i_3_n_0 : STD_LOGIC;
  signal W_37_19_i_4_n_0 : STD_LOGIC;
  signal W_37_19_i_5_n_0 : STD_LOGIC;
  signal W_37_19_i_6_n_0 : STD_LOGIC;
  signal W_37_19_i_7_n_0 : STD_LOGIC;
  signal W_37_19_i_8_n_0 : STD_LOGIC;
  signal W_37_19_i_9_n_0 : STD_LOGIC;
  signal W_37_23_i_10_n_0 : STD_LOGIC;
  signal W_37_23_i_11_n_0 : STD_LOGIC;
  signal W_37_23_i_12_n_0 : STD_LOGIC;
  signal W_37_23_i_13_n_0 : STD_LOGIC;
  signal W_37_23_i_14_n_0 : STD_LOGIC;
  signal W_37_23_i_15_n_0 : STD_LOGIC;
  signal W_37_23_i_16_n_0 : STD_LOGIC;
  signal W_37_23_i_17_n_0 : STD_LOGIC;
  signal W_37_23_i_2_n_0 : STD_LOGIC;
  signal W_37_23_i_3_n_0 : STD_LOGIC;
  signal W_37_23_i_4_n_0 : STD_LOGIC;
  signal W_37_23_i_5_n_0 : STD_LOGIC;
  signal W_37_23_i_6_n_0 : STD_LOGIC;
  signal W_37_23_i_7_n_0 : STD_LOGIC;
  signal W_37_23_i_8_n_0 : STD_LOGIC;
  signal W_37_23_i_9_n_0 : STD_LOGIC;
  signal W_37_27_i_10_n_0 : STD_LOGIC;
  signal W_37_27_i_11_n_0 : STD_LOGIC;
  signal W_37_27_i_12_n_0 : STD_LOGIC;
  signal W_37_27_i_13_n_0 : STD_LOGIC;
  signal W_37_27_i_14_n_0 : STD_LOGIC;
  signal W_37_27_i_15_n_0 : STD_LOGIC;
  signal W_37_27_i_16_n_0 : STD_LOGIC;
  signal W_37_27_i_17_n_0 : STD_LOGIC;
  signal W_37_27_i_2_n_0 : STD_LOGIC;
  signal W_37_27_i_3_n_0 : STD_LOGIC;
  signal W_37_27_i_4_n_0 : STD_LOGIC;
  signal W_37_27_i_5_n_0 : STD_LOGIC;
  signal W_37_27_i_6_n_0 : STD_LOGIC;
  signal W_37_27_i_7_n_0 : STD_LOGIC;
  signal W_37_27_i_8_n_0 : STD_LOGIC;
  signal W_37_27_i_9_n_0 : STD_LOGIC;
  signal W_37_31_i_10_n_0 : STD_LOGIC;
  signal W_37_31_i_11_n_0 : STD_LOGIC;
  signal W_37_31_i_12_n_0 : STD_LOGIC;
  signal W_37_31_i_13_n_0 : STD_LOGIC;
  signal W_37_31_i_14_n_0 : STD_LOGIC;
  signal W_37_31_i_15_n_0 : STD_LOGIC;
  signal W_37_31_i_17_n_0 : STD_LOGIC;
  signal W_37_31_i_19_n_0 : STD_LOGIC;
  signal W_37_31_i_2_n_0 : STD_LOGIC;
  signal W_37_31_i_3_n_0 : STD_LOGIC;
  signal W_37_31_i_4_n_0 : STD_LOGIC;
  signal W_37_31_i_5_n_0 : STD_LOGIC;
  signal W_37_31_i_6_n_0 : STD_LOGIC;
  signal W_37_31_i_7_n_0 : STD_LOGIC;
  signal W_37_31_i_8_n_0 : STD_LOGIC;
  signal W_37_31_i_9_n_0 : STD_LOGIC;
  signal W_37_3_i_10_n_0 : STD_LOGIC;
  signal W_37_3_i_11_n_0 : STD_LOGIC;
  signal W_37_3_i_15_n_0 : STD_LOGIC;
  signal W_37_3_i_2_n_0 : STD_LOGIC;
  signal W_37_3_i_3_n_0 : STD_LOGIC;
  signal W_37_3_i_4_n_0 : STD_LOGIC;
  signal W_37_3_i_5_n_0 : STD_LOGIC;
  signal W_37_3_i_6_n_0 : STD_LOGIC;
  signal W_37_3_i_7_n_0 : STD_LOGIC;
  signal W_37_3_i_8_n_0 : STD_LOGIC;
  signal W_37_3_i_9_n_0 : STD_LOGIC;
  signal W_37_7_i_10_n_0 : STD_LOGIC;
  signal W_37_7_i_11_n_0 : STD_LOGIC;
  signal W_37_7_i_12_n_0 : STD_LOGIC;
  signal W_37_7_i_13_n_0 : STD_LOGIC;
  signal W_37_7_i_14_n_0 : STD_LOGIC;
  signal W_37_7_i_15_n_0 : STD_LOGIC;
  signal W_37_7_i_16_n_0 : STD_LOGIC;
  signal W_37_7_i_17_n_0 : STD_LOGIC;
  signal W_37_7_i_2_n_0 : STD_LOGIC;
  signal W_37_7_i_3_n_0 : STD_LOGIC;
  signal W_37_7_i_4_n_0 : STD_LOGIC;
  signal W_37_7_i_5_n_0 : STD_LOGIC;
  signal W_37_7_i_6_n_0 : STD_LOGIC;
  signal W_37_7_i_7_n_0 : STD_LOGIC;
  signal W_37_7_i_8_n_0 : STD_LOGIC;
  signal W_37_7_i_9_n_0 : STD_LOGIC;
  signal W_38_11_i_10_n_0 : STD_LOGIC;
  signal W_38_11_i_11_n_0 : STD_LOGIC;
  signal W_38_11_i_12_n_0 : STD_LOGIC;
  signal W_38_11_i_13_n_0 : STD_LOGIC;
  signal W_38_11_i_14_n_0 : STD_LOGIC;
  signal W_38_11_i_15_n_0 : STD_LOGIC;
  signal W_38_11_i_16_n_0 : STD_LOGIC;
  signal W_38_11_i_17_n_0 : STD_LOGIC;
  signal W_38_11_i_2_n_0 : STD_LOGIC;
  signal W_38_11_i_3_n_0 : STD_LOGIC;
  signal W_38_11_i_4_n_0 : STD_LOGIC;
  signal W_38_11_i_5_n_0 : STD_LOGIC;
  signal W_38_11_i_6_n_0 : STD_LOGIC;
  signal W_38_11_i_7_n_0 : STD_LOGIC;
  signal W_38_11_i_8_n_0 : STD_LOGIC;
  signal W_38_11_i_9_n_0 : STD_LOGIC;
  signal W_38_15_i_10_n_0 : STD_LOGIC;
  signal W_38_15_i_11_n_0 : STD_LOGIC;
  signal W_38_15_i_12_n_0 : STD_LOGIC;
  signal W_38_15_i_13_n_0 : STD_LOGIC;
  signal W_38_15_i_14_n_0 : STD_LOGIC;
  signal W_38_15_i_15_n_0 : STD_LOGIC;
  signal W_38_15_i_16_n_0 : STD_LOGIC;
  signal W_38_15_i_17_n_0 : STD_LOGIC;
  signal W_38_15_i_2_n_0 : STD_LOGIC;
  signal W_38_15_i_3_n_0 : STD_LOGIC;
  signal W_38_15_i_4_n_0 : STD_LOGIC;
  signal W_38_15_i_5_n_0 : STD_LOGIC;
  signal W_38_15_i_6_n_0 : STD_LOGIC;
  signal W_38_15_i_7_n_0 : STD_LOGIC;
  signal W_38_15_i_8_n_0 : STD_LOGIC;
  signal W_38_15_i_9_n_0 : STD_LOGIC;
  signal W_38_19_i_10_n_0 : STD_LOGIC;
  signal W_38_19_i_11_n_0 : STD_LOGIC;
  signal W_38_19_i_12_n_0 : STD_LOGIC;
  signal W_38_19_i_13_n_0 : STD_LOGIC;
  signal W_38_19_i_14_n_0 : STD_LOGIC;
  signal W_38_19_i_15_n_0 : STD_LOGIC;
  signal W_38_19_i_16_n_0 : STD_LOGIC;
  signal W_38_19_i_17_n_0 : STD_LOGIC;
  signal W_38_19_i_2_n_0 : STD_LOGIC;
  signal W_38_19_i_3_n_0 : STD_LOGIC;
  signal W_38_19_i_4_n_0 : STD_LOGIC;
  signal W_38_19_i_5_n_0 : STD_LOGIC;
  signal W_38_19_i_6_n_0 : STD_LOGIC;
  signal W_38_19_i_7_n_0 : STD_LOGIC;
  signal W_38_19_i_8_n_0 : STD_LOGIC;
  signal W_38_19_i_9_n_0 : STD_LOGIC;
  signal W_38_23_i_10_n_0 : STD_LOGIC;
  signal W_38_23_i_11_n_0 : STD_LOGIC;
  signal W_38_23_i_12_n_0 : STD_LOGIC;
  signal W_38_23_i_13_n_0 : STD_LOGIC;
  signal W_38_23_i_14_n_0 : STD_LOGIC;
  signal W_38_23_i_15_n_0 : STD_LOGIC;
  signal W_38_23_i_16_n_0 : STD_LOGIC;
  signal W_38_23_i_17_n_0 : STD_LOGIC;
  signal W_38_23_i_2_n_0 : STD_LOGIC;
  signal W_38_23_i_3_n_0 : STD_LOGIC;
  signal W_38_23_i_4_n_0 : STD_LOGIC;
  signal W_38_23_i_5_n_0 : STD_LOGIC;
  signal W_38_23_i_6_n_0 : STD_LOGIC;
  signal W_38_23_i_7_n_0 : STD_LOGIC;
  signal W_38_23_i_8_n_0 : STD_LOGIC;
  signal W_38_23_i_9_n_0 : STD_LOGIC;
  signal W_38_27_i_10_n_0 : STD_LOGIC;
  signal W_38_27_i_11_n_0 : STD_LOGIC;
  signal W_38_27_i_12_n_0 : STD_LOGIC;
  signal W_38_27_i_13_n_0 : STD_LOGIC;
  signal W_38_27_i_14_n_0 : STD_LOGIC;
  signal W_38_27_i_15_n_0 : STD_LOGIC;
  signal W_38_27_i_16_n_0 : STD_LOGIC;
  signal W_38_27_i_17_n_0 : STD_LOGIC;
  signal W_38_27_i_2_n_0 : STD_LOGIC;
  signal W_38_27_i_3_n_0 : STD_LOGIC;
  signal W_38_27_i_4_n_0 : STD_LOGIC;
  signal W_38_27_i_5_n_0 : STD_LOGIC;
  signal W_38_27_i_6_n_0 : STD_LOGIC;
  signal W_38_27_i_7_n_0 : STD_LOGIC;
  signal W_38_27_i_8_n_0 : STD_LOGIC;
  signal W_38_27_i_9_n_0 : STD_LOGIC;
  signal W_38_31_i_10_n_0 : STD_LOGIC;
  signal W_38_31_i_11_n_0 : STD_LOGIC;
  signal W_38_31_i_12_n_0 : STD_LOGIC;
  signal W_38_31_i_13_n_0 : STD_LOGIC;
  signal W_38_31_i_14_n_0 : STD_LOGIC;
  signal W_38_31_i_15_n_0 : STD_LOGIC;
  signal W_38_31_i_17_n_0 : STD_LOGIC;
  signal W_38_31_i_19_n_0 : STD_LOGIC;
  signal W_38_31_i_2_n_0 : STD_LOGIC;
  signal W_38_31_i_3_n_0 : STD_LOGIC;
  signal W_38_31_i_4_n_0 : STD_LOGIC;
  signal W_38_31_i_5_n_0 : STD_LOGIC;
  signal W_38_31_i_6_n_0 : STD_LOGIC;
  signal W_38_31_i_7_n_0 : STD_LOGIC;
  signal W_38_31_i_8_n_0 : STD_LOGIC;
  signal W_38_31_i_9_n_0 : STD_LOGIC;
  signal W_38_3_i_10_n_0 : STD_LOGIC;
  signal W_38_3_i_11_n_0 : STD_LOGIC;
  signal W_38_3_i_15_n_0 : STD_LOGIC;
  signal W_38_3_i_2_n_0 : STD_LOGIC;
  signal W_38_3_i_3_n_0 : STD_LOGIC;
  signal W_38_3_i_4_n_0 : STD_LOGIC;
  signal W_38_3_i_5_n_0 : STD_LOGIC;
  signal W_38_3_i_6_n_0 : STD_LOGIC;
  signal W_38_3_i_7_n_0 : STD_LOGIC;
  signal W_38_3_i_8_n_0 : STD_LOGIC;
  signal W_38_3_i_9_n_0 : STD_LOGIC;
  signal W_38_7_i_10_n_0 : STD_LOGIC;
  signal W_38_7_i_11_n_0 : STD_LOGIC;
  signal W_38_7_i_12_n_0 : STD_LOGIC;
  signal W_38_7_i_13_n_0 : STD_LOGIC;
  signal W_38_7_i_14_n_0 : STD_LOGIC;
  signal W_38_7_i_15_n_0 : STD_LOGIC;
  signal W_38_7_i_16_n_0 : STD_LOGIC;
  signal W_38_7_i_17_n_0 : STD_LOGIC;
  signal W_38_7_i_2_n_0 : STD_LOGIC;
  signal W_38_7_i_3_n_0 : STD_LOGIC;
  signal W_38_7_i_4_n_0 : STD_LOGIC;
  signal W_38_7_i_5_n_0 : STD_LOGIC;
  signal W_38_7_i_6_n_0 : STD_LOGIC;
  signal W_38_7_i_7_n_0 : STD_LOGIC;
  signal W_38_7_i_8_n_0 : STD_LOGIC;
  signal W_38_7_i_9_n_0 : STD_LOGIC;
  signal W_39_11_i_10_n_0 : STD_LOGIC;
  signal W_39_11_i_11_n_0 : STD_LOGIC;
  signal W_39_11_i_12_n_0 : STD_LOGIC;
  signal W_39_11_i_13_n_0 : STD_LOGIC;
  signal W_39_11_i_14_n_0 : STD_LOGIC;
  signal W_39_11_i_15_n_0 : STD_LOGIC;
  signal W_39_11_i_16_n_0 : STD_LOGIC;
  signal W_39_11_i_17_n_0 : STD_LOGIC;
  signal W_39_11_i_2_n_0 : STD_LOGIC;
  signal W_39_11_i_3_n_0 : STD_LOGIC;
  signal W_39_11_i_4_n_0 : STD_LOGIC;
  signal W_39_11_i_5_n_0 : STD_LOGIC;
  signal W_39_11_i_6_n_0 : STD_LOGIC;
  signal W_39_11_i_7_n_0 : STD_LOGIC;
  signal W_39_11_i_8_n_0 : STD_LOGIC;
  signal W_39_11_i_9_n_0 : STD_LOGIC;
  signal W_39_15_i_10_n_0 : STD_LOGIC;
  signal W_39_15_i_11_n_0 : STD_LOGIC;
  signal W_39_15_i_12_n_0 : STD_LOGIC;
  signal W_39_15_i_13_n_0 : STD_LOGIC;
  signal W_39_15_i_14_n_0 : STD_LOGIC;
  signal W_39_15_i_15_n_0 : STD_LOGIC;
  signal W_39_15_i_16_n_0 : STD_LOGIC;
  signal W_39_15_i_17_n_0 : STD_LOGIC;
  signal W_39_15_i_2_n_0 : STD_LOGIC;
  signal W_39_15_i_3_n_0 : STD_LOGIC;
  signal W_39_15_i_4_n_0 : STD_LOGIC;
  signal W_39_15_i_5_n_0 : STD_LOGIC;
  signal W_39_15_i_6_n_0 : STD_LOGIC;
  signal W_39_15_i_7_n_0 : STD_LOGIC;
  signal W_39_15_i_8_n_0 : STD_LOGIC;
  signal W_39_15_i_9_n_0 : STD_LOGIC;
  signal W_39_19_i_10_n_0 : STD_LOGIC;
  signal W_39_19_i_11_n_0 : STD_LOGIC;
  signal W_39_19_i_12_n_0 : STD_LOGIC;
  signal W_39_19_i_13_n_0 : STD_LOGIC;
  signal W_39_19_i_14_n_0 : STD_LOGIC;
  signal W_39_19_i_15_n_0 : STD_LOGIC;
  signal W_39_19_i_16_n_0 : STD_LOGIC;
  signal W_39_19_i_17_n_0 : STD_LOGIC;
  signal W_39_19_i_2_n_0 : STD_LOGIC;
  signal W_39_19_i_3_n_0 : STD_LOGIC;
  signal W_39_19_i_4_n_0 : STD_LOGIC;
  signal W_39_19_i_5_n_0 : STD_LOGIC;
  signal W_39_19_i_6_n_0 : STD_LOGIC;
  signal W_39_19_i_7_n_0 : STD_LOGIC;
  signal W_39_19_i_8_n_0 : STD_LOGIC;
  signal W_39_19_i_9_n_0 : STD_LOGIC;
  signal W_39_23_i_10_n_0 : STD_LOGIC;
  signal W_39_23_i_11_n_0 : STD_LOGIC;
  signal W_39_23_i_12_n_0 : STD_LOGIC;
  signal W_39_23_i_13_n_0 : STD_LOGIC;
  signal W_39_23_i_14_n_0 : STD_LOGIC;
  signal W_39_23_i_15_n_0 : STD_LOGIC;
  signal W_39_23_i_16_n_0 : STD_LOGIC;
  signal W_39_23_i_17_n_0 : STD_LOGIC;
  signal W_39_23_i_2_n_0 : STD_LOGIC;
  signal W_39_23_i_3_n_0 : STD_LOGIC;
  signal W_39_23_i_4_n_0 : STD_LOGIC;
  signal W_39_23_i_5_n_0 : STD_LOGIC;
  signal W_39_23_i_6_n_0 : STD_LOGIC;
  signal W_39_23_i_7_n_0 : STD_LOGIC;
  signal W_39_23_i_8_n_0 : STD_LOGIC;
  signal W_39_23_i_9_n_0 : STD_LOGIC;
  signal W_39_27_i_10_n_0 : STD_LOGIC;
  signal W_39_27_i_11_n_0 : STD_LOGIC;
  signal W_39_27_i_12_n_0 : STD_LOGIC;
  signal W_39_27_i_13_n_0 : STD_LOGIC;
  signal W_39_27_i_14_n_0 : STD_LOGIC;
  signal W_39_27_i_15_n_0 : STD_LOGIC;
  signal W_39_27_i_16_n_0 : STD_LOGIC;
  signal W_39_27_i_17_n_0 : STD_LOGIC;
  signal W_39_27_i_2_n_0 : STD_LOGIC;
  signal W_39_27_i_3_n_0 : STD_LOGIC;
  signal W_39_27_i_4_n_0 : STD_LOGIC;
  signal W_39_27_i_5_n_0 : STD_LOGIC;
  signal W_39_27_i_6_n_0 : STD_LOGIC;
  signal W_39_27_i_7_n_0 : STD_LOGIC;
  signal W_39_27_i_8_n_0 : STD_LOGIC;
  signal W_39_27_i_9_n_0 : STD_LOGIC;
  signal W_39_31_i_10_n_0 : STD_LOGIC;
  signal W_39_31_i_11_n_0 : STD_LOGIC;
  signal W_39_31_i_12_n_0 : STD_LOGIC;
  signal W_39_31_i_13_n_0 : STD_LOGIC;
  signal W_39_31_i_14_n_0 : STD_LOGIC;
  signal W_39_31_i_15_n_0 : STD_LOGIC;
  signal W_39_31_i_17_n_0 : STD_LOGIC;
  signal W_39_31_i_19_n_0 : STD_LOGIC;
  signal W_39_31_i_2_n_0 : STD_LOGIC;
  signal W_39_31_i_3_n_0 : STD_LOGIC;
  signal W_39_31_i_4_n_0 : STD_LOGIC;
  signal W_39_31_i_5_n_0 : STD_LOGIC;
  signal W_39_31_i_6_n_0 : STD_LOGIC;
  signal W_39_31_i_7_n_0 : STD_LOGIC;
  signal W_39_31_i_8_n_0 : STD_LOGIC;
  signal W_39_31_i_9_n_0 : STD_LOGIC;
  signal W_39_3_i_10_n_0 : STD_LOGIC;
  signal W_39_3_i_11_n_0 : STD_LOGIC;
  signal W_39_3_i_15_n_0 : STD_LOGIC;
  signal W_39_3_i_2_n_0 : STD_LOGIC;
  signal W_39_3_i_3_n_0 : STD_LOGIC;
  signal W_39_3_i_4_n_0 : STD_LOGIC;
  signal W_39_3_i_5_n_0 : STD_LOGIC;
  signal W_39_3_i_6_n_0 : STD_LOGIC;
  signal W_39_3_i_7_n_0 : STD_LOGIC;
  signal W_39_3_i_8_n_0 : STD_LOGIC;
  signal W_39_3_i_9_n_0 : STD_LOGIC;
  signal W_39_7_i_10_n_0 : STD_LOGIC;
  signal W_39_7_i_11_n_0 : STD_LOGIC;
  signal W_39_7_i_12_n_0 : STD_LOGIC;
  signal W_39_7_i_13_n_0 : STD_LOGIC;
  signal W_39_7_i_14_n_0 : STD_LOGIC;
  signal W_39_7_i_15_n_0 : STD_LOGIC;
  signal W_39_7_i_16_n_0 : STD_LOGIC;
  signal W_39_7_i_17_n_0 : STD_LOGIC;
  signal W_39_7_i_2_n_0 : STD_LOGIC;
  signal W_39_7_i_3_n_0 : STD_LOGIC;
  signal W_39_7_i_4_n_0 : STD_LOGIC;
  signal W_39_7_i_5_n_0 : STD_LOGIC;
  signal W_39_7_i_6_n_0 : STD_LOGIC;
  signal W_39_7_i_7_n_0 : STD_LOGIC;
  signal W_39_7_i_8_n_0 : STD_LOGIC;
  signal W_39_7_i_9_n_0 : STD_LOGIC;
  signal W_40_11_i_10_n_0 : STD_LOGIC;
  signal W_40_11_i_11_n_0 : STD_LOGIC;
  signal W_40_11_i_12_n_0 : STD_LOGIC;
  signal W_40_11_i_13_n_0 : STD_LOGIC;
  signal W_40_11_i_14_n_0 : STD_LOGIC;
  signal W_40_11_i_15_n_0 : STD_LOGIC;
  signal W_40_11_i_16_n_0 : STD_LOGIC;
  signal W_40_11_i_17_n_0 : STD_LOGIC;
  signal W_40_11_i_2_n_0 : STD_LOGIC;
  signal W_40_11_i_3_n_0 : STD_LOGIC;
  signal W_40_11_i_4_n_0 : STD_LOGIC;
  signal W_40_11_i_5_n_0 : STD_LOGIC;
  signal W_40_11_i_6_n_0 : STD_LOGIC;
  signal W_40_11_i_7_n_0 : STD_LOGIC;
  signal W_40_11_i_8_n_0 : STD_LOGIC;
  signal W_40_11_i_9_n_0 : STD_LOGIC;
  signal W_40_15_i_10_n_0 : STD_LOGIC;
  signal W_40_15_i_11_n_0 : STD_LOGIC;
  signal W_40_15_i_12_n_0 : STD_LOGIC;
  signal W_40_15_i_13_n_0 : STD_LOGIC;
  signal W_40_15_i_14_n_0 : STD_LOGIC;
  signal W_40_15_i_15_n_0 : STD_LOGIC;
  signal W_40_15_i_16_n_0 : STD_LOGIC;
  signal W_40_15_i_17_n_0 : STD_LOGIC;
  signal W_40_15_i_2_n_0 : STD_LOGIC;
  signal W_40_15_i_3_n_0 : STD_LOGIC;
  signal W_40_15_i_4_n_0 : STD_LOGIC;
  signal W_40_15_i_5_n_0 : STD_LOGIC;
  signal W_40_15_i_6_n_0 : STD_LOGIC;
  signal W_40_15_i_7_n_0 : STD_LOGIC;
  signal W_40_15_i_8_n_0 : STD_LOGIC;
  signal W_40_15_i_9_n_0 : STD_LOGIC;
  signal W_40_19_i_10_n_0 : STD_LOGIC;
  signal W_40_19_i_11_n_0 : STD_LOGIC;
  signal W_40_19_i_12_n_0 : STD_LOGIC;
  signal W_40_19_i_13_n_0 : STD_LOGIC;
  signal W_40_19_i_14_n_0 : STD_LOGIC;
  signal W_40_19_i_15_n_0 : STD_LOGIC;
  signal W_40_19_i_16_n_0 : STD_LOGIC;
  signal W_40_19_i_17_n_0 : STD_LOGIC;
  signal W_40_19_i_2_n_0 : STD_LOGIC;
  signal W_40_19_i_3_n_0 : STD_LOGIC;
  signal W_40_19_i_4_n_0 : STD_LOGIC;
  signal W_40_19_i_5_n_0 : STD_LOGIC;
  signal W_40_19_i_6_n_0 : STD_LOGIC;
  signal W_40_19_i_7_n_0 : STD_LOGIC;
  signal W_40_19_i_8_n_0 : STD_LOGIC;
  signal W_40_19_i_9_n_0 : STD_LOGIC;
  signal W_40_23_i_10_n_0 : STD_LOGIC;
  signal W_40_23_i_11_n_0 : STD_LOGIC;
  signal W_40_23_i_12_n_0 : STD_LOGIC;
  signal W_40_23_i_13_n_0 : STD_LOGIC;
  signal W_40_23_i_14_n_0 : STD_LOGIC;
  signal W_40_23_i_15_n_0 : STD_LOGIC;
  signal W_40_23_i_16_n_0 : STD_LOGIC;
  signal W_40_23_i_17_n_0 : STD_LOGIC;
  signal W_40_23_i_2_n_0 : STD_LOGIC;
  signal W_40_23_i_3_n_0 : STD_LOGIC;
  signal W_40_23_i_4_n_0 : STD_LOGIC;
  signal W_40_23_i_5_n_0 : STD_LOGIC;
  signal W_40_23_i_6_n_0 : STD_LOGIC;
  signal W_40_23_i_7_n_0 : STD_LOGIC;
  signal W_40_23_i_8_n_0 : STD_LOGIC;
  signal W_40_23_i_9_n_0 : STD_LOGIC;
  signal W_40_27_i_10_n_0 : STD_LOGIC;
  signal W_40_27_i_11_n_0 : STD_LOGIC;
  signal W_40_27_i_12_n_0 : STD_LOGIC;
  signal W_40_27_i_13_n_0 : STD_LOGIC;
  signal W_40_27_i_14_n_0 : STD_LOGIC;
  signal W_40_27_i_15_n_0 : STD_LOGIC;
  signal W_40_27_i_16_n_0 : STD_LOGIC;
  signal W_40_27_i_17_n_0 : STD_LOGIC;
  signal W_40_27_i_2_n_0 : STD_LOGIC;
  signal W_40_27_i_3_n_0 : STD_LOGIC;
  signal W_40_27_i_4_n_0 : STD_LOGIC;
  signal W_40_27_i_5_n_0 : STD_LOGIC;
  signal W_40_27_i_6_n_0 : STD_LOGIC;
  signal W_40_27_i_7_n_0 : STD_LOGIC;
  signal W_40_27_i_8_n_0 : STD_LOGIC;
  signal W_40_27_i_9_n_0 : STD_LOGIC;
  signal W_40_31_i_10_n_0 : STD_LOGIC;
  signal W_40_31_i_11_n_0 : STD_LOGIC;
  signal W_40_31_i_12_n_0 : STD_LOGIC;
  signal W_40_31_i_13_n_0 : STD_LOGIC;
  signal W_40_31_i_14_n_0 : STD_LOGIC;
  signal W_40_31_i_15_n_0 : STD_LOGIC;
  signal W_40_31_i_17_n_0 : STD_LOGIC;
  signal W_40_31_i_19_n_0 : STD_LOGIC;
  signal W_40_31_i_2_n_0 : STD_LOGIC;
  signal W_40_31_i_3_n_0 : STD_LOGIC;
  signal W_40_31_i_4_n_0 : STD_LOGIC;
  signal W_40_31_i_5_n_0 : STD_LOGIC;
  signal W_40_31_i_6_n_0 : STD_LOGIC;
  signal W_40_31_i_7_n_0 : STD_LOGIC;
  signal W_40_31_i_8_n_0 : STD_LOGIC;
  signal W_40_31_i_9_n_0 : STD_LOGIC;
  signal W_40_3_i_10_n_0 : STD_LOGIC;
  signal W_40_3_i_11_n_0 : STD_LOGIC;
  signal W_40_3_i_15_n_0 : STD_LOGIC;
  signal W_40_3_i_2_n_0 : STD_LOGIC;
  signal W_40_3_i_3_n_0 : STD_LOGIC;
  signal W_40_3_i_4_n_0 : STD_LOGIC;
  signal W_40_3_i_5_n_0 : STD_LOGIC;
  signal W_40_3_i_6_n_0 : STD_LOGIC;
  signal W_40_3_i_7_n_0 : STD_LOGIC;
  signal W_40_3_i_8_n_0 : STD_LOGIC;
  signal W_40_3_i_9_n_0 : STD_LOGIC;
  signal W_40_7_i_10_n_0 : STD_LOGIC;
  signal W_40_7_i_11_n_0 : STD_LOGIC;
  signal W_40_7_i_12_n_0 : STD_LOGIC;
  signal W_40_7_i_13_n_0 : STD_LOGIC;
  signal W_40_7_i_14_n_0 : STD_LOGIC;
  signal W_40_7_i_15_n_0 : STD_LOGIC;
  signal W_40_7_i_16_n_0 : STD_LOGIC;
  signal W_40_7_i_17_n_0 : STD_LOGIC;
  signal W_40_7_i_2_n_0 : STD_LOGIC;
  signal W_40_7_i_3_n_0 : STD_LOGIC;
  signal W_40_7_i_4_n_0 : STD_LOGIC;
  signal W_40_7_i_5_n_0 : STD_LOGIC;
  signal W_40_7_i_6_n_0 : STD_LOGIC;
  signal W_40_7_i_7_n_0 : STD_LOGIC;
  signal W_40_7_i_8_n_0 : STD_LOGIC;
  signal W_40_7_i_9_n_0 : STD_LOGIC;
  signal W_41_11_i_10_n_0 : STD_LOGIC;
  signal W_41_11_i_11_n_0 : STD_LOGIC;
  signal W_41_11_i_12_n_0 : STD_LOGIC;
  signal W_41_11_i_13_n_0 : STD_LOGIC;
  signal W_41_11_i_14_n_0 : STD_LOGIC;
  signal W_41_11_i_15_n_0 : STD_LOGIC;
  signal W_41_11_i_16_n_0 : STD_LOGIC;
  signal W_41_11_i_17_n_0 : STD_LOGIC;
  signal W_41_11_i_2_n_0 : STD_LOGIC;
  signal W_41_11_i_3_n_0 : STD_LOGIC;
  signal W_41_11_i_4_n_0 : STD_LOGIC;
  signal W_41_11_i_5_n_0 : STD_LOGIC;
  signal W_41_11_i_6_n_0 : STD_LOGIC;
  signal W_41_11_i_7_n_0 : STD_LOGIC;
  signal W_41_11_i_8_n_0 : STD_LOGIC;
  signal W_41_11_i_9_n_0 : STD_LOGIC;
  signal W_41_15_i_10_n_0 : STD_LOGIC;
  signal W_41_15_i_11_n_0 : STD_LOGIC;
  signal W_41_15_i_12_n_0 : STD_LOGIC;
  signal W_41_15_i_13_n_0 : STD_LOGIC;
  signal W_41_15_i_14_n_0 : STD_LOGIC;
  signal W_41_15_i_15_n_0 : STD_LOGIC;
  signal W_41_15_i_16_n_0 : STD_LOGIC;
  signal W_41_15_i_17_n_0 : STD_LOGIC;
  signal W_41_15_i_2_n_0 : STD_LOGIC;
  signal W_41_15_i_3_n_0 : STD_LOGIC;
  signal W_41_15_i_4_n_0 : STD_LOGIC;
  signal W_41_15_i_5_n_0 : STD_LOGIC;
  signal W_41_15_i_6_n_0 : STD_LOGIC;
  signal W_41_15_i_7_n_0 : STD_LOGIC;
  signal W_41_15_i_8_n_0 : STD_LOGIC;
  signal W_41_15_i_9_n_0 : STD_LOGIC;
  signal W_41_19_i_10_n_0 : STD_LOGIC;
  signal W_41_19_i_11_n_0 : STD_LOGIC;
  signal W_41_19_i_12_n_0 : STD_LOGIC;
  signal W_41_19_i_13_n_0 : STD_LOGIC;
  signal W_41_19_i_14_n_0 : STD_LOGIC;
  signal W_41_19_i_15_n_0 : STD_LOGIC;
  signal W_41_19_i_16_n_0 : STD_LOGIC;
  signal W_41_19_i_17_n_0 : STD_LOGIC;
  signal W_41_19_i_2_n_0 : STD_LOGIC;
  signal W_41_19_i_3_n_0 : STD_LOGIC;
  signal W_41_19_i_4_n_0 : STD_LOGIC;
  signal W_41_19_i_5_n_0 : STD_LOGIC;
  signal W_41_19_i_6_n_0 : STD_LOGIC;
  signal W_41_19_i_7_n_0 : STD_LOGIC;
  signal W_41_19_i_8_n_0 : STD_LOGIC;
  signal W_41_19_i_9_n_0 : STD_LOGIC;
  signal W_41_23_i_10_n_0 : STD_LOGIC;
  signal W_41_23_i_11_n_0 : STD_LOGIC;
  signal W_41_23_i_12_n_0 : STD_LOGIC;
  signal W_41_23_i_13_n_0 : STD_LOGIC;
  signal W_41_23_i_14_n_0 : STD_LOGIC;
  signal W_41_23_i_15_n_0 : STD_LOGIC;
  signal W_41_23_i_16_n_0 : STD_LOGIC;
  signal W_41_23_i_17_n_0 : STD_LOGIC;
  signal W_41_23_i_2_n_0 : STD_LOGIC;
  signal W_41_23_i_3_n_0 : STD_LOGIC;
  signal W_41_23_i_4_n_0 : STD_LOGIC;
  signal W_41_23_i_5_n_0 : STD_LOGIC;
  signal W_41_23_i_6_n_0 : STD_LOGIC;
  signal W_41_23_i_7_n_0 : STD_LOGIC;
  signal W_41_23_i_8_n_0 : STD_LOGIC;
  signal W_41_23_i_9_n_0 : STD_LOGIC;
  signal W_41_27_i_10_n_0 : STD_LOGIC;
  signal W_41_27_i_11_n_0 : STD_LOGIC;
  signal W_41_27_i_12_n_0 : STD_LOGIC;
  signal W_41_27_i_13_n_0 : STD_LOGIC;
  signal W_41_27_i_14_n_0 : STD_LOGIC;
  signal W_41_27_i_15_n_0 : STD_LOGIC;
  signal W_41_27_i_16_n_0 : STD_LOGIC;
  signal W_41_27_i_17_n_0 : STD_LOGIC;
  signal W_41_27_i_2_n_0 : STD_LOGIC;
  signal W_41_27_i_3_n_0 : STD_LOGIC;
  signal W_41_27_i_4_n_0 : STD_LOGIC;
  signal W_41_27_i_5_n_0 : STD_LOGIC;
  signal W_41_27_i_6_n_0 : STD_LOGIC;
  signal W_41_27_i_7_n_0 : STD_LOGIC;
  signal W_41_27_i_8_n_0 : STD_LOGIC;
  signal W_41_27_i_9_n_0 : STD_LOGIC;
  signal W_41_31_i_10_n_0 : STD_LOGIC;
  signal W_41_31_i_11_n_0 : STD_LOGIC;
  signal W_41_31_i_12_n_0 : STD_LOGIC;
  signal W_41_31_i_13_n_0 : STD_LOGIC;
  signal W_41_31_i_14_n_0 : STD_LOGIC;
  signal W_41_31_i_15_n_0 : STD_LOGIC;
  signal W_41_31_i_17_n_0 : STD_LOGIC;
  signal W_41_31_i_19_n_0 : STD_LOGIC;
  signal W_41_31_i_2_n_0 : STD_LOGIC;
  signal W_41_31_i_3_n_0 : STD_LOGIC;
  signal W_41_31_i_4_n_0 : STD_LOGIC;
  signal W_41_31_i_5_n_0 : STD_LOGIC;
  signal W_41_31_i_6_n_0 : STD_LOGIC;
  signal W_41_31_i_7_n_0 : STD_LOGIC;
  signal W_41_31_i_8_n_0 : STD_LOGIC;
  signal W_41_31_i_9_n_0 : STD_LOGIC;
  signal W_41_3_i_10_n_0 : STD_LOGIC;
  signal W_41_3_i_11_n_0 : STD_LOGIC;
  signal W_41_3_i_15_n_0 : STD_LOGIC;
  signal W_41_3_i_2_n_0 : STD_LOGIC;
  signal W_41_3_i_3_n_0 : STD_LOGIC;
  signal W_41_3_i_4_n_0 : STD_LOGIC;
  signal W_41_3_i_5_n_0 : STD_LOGIC;
  signal W_41_3_i_6_n_0 : STD_LOGIC;
  signal W_41_3_i_7_n_0 : STD_LOGIC;
  signal W_41_3_i_8_n_0 : STD_LOGIC;
  signal W_41_3_i_9_n_0 : STD_LOGIC;
  signal W_41_7_i_10_n_0 : STD_LOGIC;
  signal W_41_7_i_11_n_0 : STD_LOGIC;
  signal W_41_7_i_12_n_0 : STD_LOGIC;
  signal W_41_7_i_13_n_0 : STD_LOGIC;
  signal W_41_7_i_14_n_0 : STD_LOGIC;
  signal W_41_7_i_15_n_0 : STD_LOGIC;
  signal W_41_7_i_16_n_0 : STD_LOGIC;
  signal W_41_7_i_17_n_0 : STD_LOGIC;
  signal W_41_7_i_2_n_0 : STD_LOGIC;
  signal W_41_7_i_3_n_0 : STD_LOGIC;
  signal W_41_7_i_4_n_0 : STD_LOGIC;
  signal W_41_7_i_5_n_0 : STD_LOGIC;
  signal W_41_7_i_6_n_0 : STD_LOGIC;
  signal W_41_7_i_7_n_0 : STD_LOGIC;
  signal W_41_7_i_8_n_0 : STD_LOGIC;
  signal W_41_7_i_9_n_0 : STD_LOGIC;
  signal W_42_11_i_10_n_0 : STD_LOGIC;
  signal W_42_11_i_11_n_0 : STD_LOGIC;
  signal W_42_11_i_12_n_0 : STD_LOGIC;
  signal W_42_11_i_13_n_0 : STD_LOGIC;
  signal W_42_11_i_14_n_0 : STD_LOGIC;
  signal W_42_11_i_15_n_0 : STD_LOGIC;
  signal W_42_11_i_16_n_0 : STD_LOGIC;
  signal W_42_11_i_17_n_0 : STD_LOGIC;
  signal W_42_11_i_2_n_0 : STD_LOGIC;
  signal W_42_11_i_3_n_0 : STD_LOGIC;
  signal W_42_11_i_4_n_0 : STD_LOGIC;
  signal W_42_11_i_5_n_0 : STD_LOGIC;
  signal W_42_11_i_6_n_0 : STD_LOGIC;
  signal W_42_11_i_7_n_0 : STD_LOGIC;
  signal W_42_11_i_8_n_0 : STD_LOGIC;
  signal W_42_11_i_9_n_0 : STD_LOGIC;
  signal W_42_15_i_10_n_0 : STD_LOGIC;
  signal W_42_15_i_11_n_0 : STD_LOGIC;
  signal W_42_15_i_12_n_0 : STD_LOGIC;
  signal W_42_15_i_13_n_0 : STD_LOGIC;
  signal W_42_15_i_14_n_0 : STD_LOGIC;
  signal W_42_15_i_15_n_0 : STD_LOGIC;
  signal W_42_15_i_16_n_0 : STD_LOGIC;
  signal W_42_15_i_17_n_0 : STD_LOGIC;
  signal W_42_15_i_2_n_0 : STD_LOGIC;
  signal W_42_15_i_3_n_0 : STD_LOGIC;
  signal W_42_15_i_4_n_0 : STD_LOGIC;
  signal W_42_15_i_5_n_0 : STD_LOGIC;
  signal W_42_15_i_6_n_0 : STD_LOGIC;
  signal W_42_15_i_7_n_0 : STD_LOGIC;
  signal W_42_15_i_8_n_0 : STD_LOGIC;
  signal W_42_15_i_9_n_0 : STD_LOGIC;
  signal W_42_19_i_10_n_0 : STD_LOGIC;
  signal W_42_19_i_11_n_0 : STD_LOGIC;
  signal W_42_19_i_12_n_0 : STD_LOGIC;
  signal W_42_19_i_13_n_0 : STD_LOGIC;
  signal W_42_19_i_14_n_0 : STD_LOGIC;
  signal W_42_19_i_15_n_0 : STD_LOGIC;
  signal W_42_19_i_16_n_0 : STD_LOGIC;
  signal W_42_19_i_17_n_0 : STD_LOGIC;
  signal W_42_19_i_2_n_0 : STD_LOGIC;
  signal W_42_19_i_3_n_0 : STD_LOGIC;
  signal W_42_19_i_4_n_0 : STD_LOGIC;
  signal W_42_19_i_5_n_0 : STD_LOGIC;
  signal W_42_19_i_6_n_0 : STD_LOGIC;
  signal W_42_19_i_7_n_0 : STD_LOGIC;
  signal W_42_19_i_8_n_0 : STD_LOGIC;
  signal W_42_19_i_9_n_0 : STD_LOGIC;
  signal W_42_23_i_10_n_0 : STD_LOGIC;
  signal W_42_23_i_11_n_0 : STD_LOGIC;
  signal W_42_23_i_12_n_0 : STD_LOGIC;
  signal W_42_23_i_13_n_0 : STD_LOGIC;
  signal W_42_23_i_14_n_0 : STD_LOGIC;
  signal W_42_23_i_15_n_0 : STD_LOGIC;
  signal W_42_23_i_16_n_0 : STD_LOGIC;
  signal W_42_23_i_17_n_0 : STD_LOGIC;
  signal W_42_23_i_2_n_0 : STD_LOGIC;
  signal W_42_23_i_3_n_0 : STD_LOGIC;
  signal W_42_23_i_4_n_0 : STD_LOGIC;
  signal W_42_23_i_5_n_0 : STD_LOGIC;
  signal W_42_23_i_6_n_0 : STD_LOGIC;
  signal W_42_23_i_7_n_0 : STD_LOGIC;
  signal W_42_23_i_8_n_0 : STD_LOGIC;
  signal W_42_23_i_9_n_0 : STD_LOGIC;
  signal W_42_27_i_10_n_0 : STD_LOGIC;
  signal W_42_27_i_11_n_0 : STD_LOGIC;
  signal W_42_27_i_12_n_0 : STD_LOGIC;
  signal W_42_27_i_13_n_0 : STD_LOGIC;
  signal W_42_27_i_14_n_0 : STD_LOGIC;
  signal W_42_27_i_15_n_0 : STD_LOGIC;
  signal W_42_27_i_16_n_0 : STD_LOGIC;
  signal W_42_27_i_17_n_0 : STD_LOGIC;
  signal W_42_27_i_2_n_0 : STD_LOGIC;
  signal W_42_27_i_3_n_0 : STD_LOGIC;
  signal W_42_27_i_4_n_0 : STD_LOGIC;
  signal W_42_27_i_5_n_0 : STD_LOGIC;
  signal W_42_27_i_6_n_0 : STD_LOGIC;
  signal W_42_27_i_7_n_0 : STD_LOGIC;
  signal W_42_27_i_8_n_0 : STD_LOGIC;
  signal W_42_27_i_9_n_0 : STD_LOGIC;
  signal W_42_31_i_10_n_0 : STD_LOGIC;
  signal W_42_31_i_11_n_0 : STD_LOGIC;
  signal W_42_31_i_12_n_0 : STD_LOGIC;
  signal W_42_31_i_13_n_0 : STD_LOGIC;
  signal W_42_31_i_14_n_0 : STD_LOGIC;
  signal W_42_31_i_15_n_0 : STD_LOGIC;
  signal W_42_31_i_17_n_0 : STD_LOGIC;
  signal W_42_31_i_19_n_0 : STD_LOGIC;
  signal W_42_31_i_2_n_0 : STD_LOGIC;
  signal W_42_31_i_3_n_0 : STD_LOGIC;
  signal W_42_31_i_4_n_0 : STD_LOGIC;
  signal W_42_31_i_5_n_0 : STD_LOGIC;
  signal W_42_31_i_6_n_0 : STD_LOGIC;
  signal W_42_31_i_7_n_0 : STD_LOGIC;
  signal W_42_31_i_8_n_0 : STD_LOGIC;
  signal W_42_31_i_9_n_0 : STD_LOGIC;
  signal W_42_3_i_10_n_0 : STD_LOGIC;
  signal W_42_3_i_11_n_0 : STD_LOGIC;
  signal W_42_3_i_15_n_0 : STD_LOGIC;
  signal W_42_3_i_2_n_0 : STD_LOGIC;
  signal W_42_3_i_3_n_0 : STD_LOGIC;
  signal W_42_3_i_4_n_0 : STD_LOGIC;
  signal W_42_3_i_5_n_0 : STD_LOGIC;
  signal W_42_3_i_6_n_0 : STD_LOGIC;
  signal W_42_3_i_7_n_0 : STD_LOGIC;
  signal W_42_3_i_8_n_0 : STD_LOGIC;
  signal W_42_3_i_9_n_0 : STD_LOGIC;
  signal W_42_7_i_10_n_0 : STD_LOGIC;
  signal W_42_7_i_11_n_0 : STD_LOGIC;
  signal W_42_7_i_12_n_0 : STD_LOGIC;
  signal W_42_7_i_13_n_0 : STD_LOGIC;
  signal W_42_7_i_14_n_0 : STD_LOGIC;
  signal W_42_7_i_15_n_0 : STD_LOGIC;
  signal W_42_7_i_16_n_0 : STD_LOGIC;
  signal W_42_7_i_17_n_0 : STD_LOGIC;
  signal W_42_7_i_2_n_0 : STD_LOGIC;
  signal W_42_7_i_3_n_0 : STD_LOGIC;
  signal W_42_7_i_4_n_0 : STD_LOGIC;
  signal W_42_7_i_5_n_0 : STD_LOGIC;
  signal W_42_7_i_6_n_0 : STD_LOGIC;
  signal W_42_7_i_7_n_0 : STD_LOGIC;
  signal W_42_7_i_8_n_0 : STD_LOGIC;
  signal W_42_7_i_9_n_0 : STD_LOGIC;
  signal W_43_11_i_10_n_0 : STD_LOGIC;
  signal W_43_11_i_11_n_0 : STD_LOGIC;
  signal W_43_11_i_12_n_0 : STD_LOGIC;
  signal W_43_11_i_13_n_0 : STD_LOGIC;
  signal W_43_11_i_14_n_0 : STD_LOGIC;
  signal W_43_11_i_15_n_0 : STD_LOGIC;
  signal W_43_11_i_16_n_0 : STD_LOGIC;
  signal W_43_11_i_17_n_0 : STD_LOGIC;
  signal W_43_11_i_2_n_0 : STD_LOGIC;
  signal W_43_11_i_3_n_0 : STD_LOGIC;
  signal W_43_11_i_4_n_0 : STD_LOGIC;
  signal W_43_11_i_5_n_0 : STD_LOGIC;
  signal W_43_11_i_6_n_0 : STD_LOGIC;
  signal W_43_11_i_7_n_0 : STD_LOGIC;
  signal W_43_11_i_8_n_0 : STD_LOGIC;
  signal W_43_11_i_9_n_0 : STD_LOGIC;
  signal W_43_15_i_10_n_0 : STD_LOGIC;
  signal W_43_15_i_11_n_0 : STD_LOGIC;
  signal W_43_15_i_12_n_0 : STD_LOGIC;
  signal W_43_15_i_13_n_0 : STD_LOGIC;
  signal W_43_15_i_14_n_0 : STD_LOGIC;
  signal W_43_15_i_15_n_0 : STD_LOGIC;
  signal W_43_15_i_16_n_0 : STD_LOGIC;
  signal W_43_15_i_17_n_0 : STD_LOGIC;
  signal W_43_15_i_2_n_0 : STD_LOGIC;
  signal W_43_15_i_3_n_0 : STD_LOGIC;
  signal W_43_15_i_4_n_0 : STD_LOGIC;
  signal W_43_15_i_5_n_0 : STD_LOGIC;
  signal W_43_15_i_6_n_0 : STD_LOGIC;
  signal W_43_15_i_7_n_0 : STD_LOGIC;
  signal W_43_15_i_8_n_0 : STD_LOGIC;
  signal W_43_15_i_9_n_0 : STD_LOGIC;
  signal W_43_19_i_10_n_0 : STD_LOGIC;
  signal W_43_19_i_11_n_0 : STD_LOGIC;
  signal W_43_19_i_12_n_0 : STD_LOGIC;
  signal W_43_19_i_13_n_0 : STD_LOGIC;
  signal W_43_19_i_14_n_0 : STD_LOGIC;
  signal W_43_19_i_15_n_0 : STD_LOGIC;
  signal W_43_19_i_16_n_0 : STD_LOGIC;
  signal W_43_19_i_17_n_0 : STD_LOGIC;
  signal W_43_19_i_2_n_0 : STD_LOGIC;
  signal W_43_19_i_3_n_0 : STD_LOGIC;
  signal W_43_19_i_4_n_0 : STD_LOGIC;
  signal W_43_19_i_5_n_0 : STD_LOGIC;
  signal W_43_19_i_6_n_0 : STD_LOGIC;
  signal W_43_19_i_7_n_0 : STD_LOGIC;
  signal W_43_19_i_8_n_0 : STD_LOGIC;
  signal W_43_19_i_9_n_0 : STD_LOGIC;
  signal W_43_23_i_10_n_0 : STD_LOGIC;
  signal W_43_23_i_11_n_0 : STD_LOGIC;
  signal W_43_23_i_12_n_0 : STD_LOGIC;
  signal W_43_23_i_13_n_0 : STD_LOGIC;
  signal W_43_23_i_14_n_0 : STD_LOGIC;
  signal W_43_23_i_15_n_0 : STD_LOGIC;
  signal W_43_23_i_16_n_0 : STD_LOGIC;
  signal W_43_23_i_17_n_0 : STD_LOGIC;
  signal W_43_23_i_2_n_0 : STD_LOGIC;
  signal W_43_23_i_3_n_0 : STD_LOGIC;
  signal W_43_23_i_4_n_0 : STD_LOGIC;
  signal W_43_23_i_5_n_0 : STD_LOGIC;
  signal W_43_23_i_6_n_0 : STD_LOGIC;
  signal W_43_23_i_7_n_0 : STD_LOGIC;
  signal W_43_23_i_8_n_0 : STD_LOGIC;
  signal W_43_23_i_9_n_0 : STD_LOGIC;
  signal W_43_27_i_10_n_0 : STD_LOGIC;
  signal W_43_27_i_11_n_0 : STD_LOGIC;
  signal W_43_27_i_12_n_0 : STD_LOGIC;
  signal W_43_27_i_13_n_0 : STD_LOGIC;
  signal W_43_27_i_14_n_0 : STD_LOGIC;
  signal W_43_27_i_15_n_0 : STD_LOGIC;
  signal W_43_27_i_16_n_0 : STD_LOGIC;
  signal W_43_27_i_17_n_0 : STD_LOGIC;
  signal W_43_27_i_2_n_0 : STD_LOGIC;
  signal W_43_27_i_3_n_0 : STD_LOGIC;
  signal W_43_27_i_4_n_0 : STD_LOGIC;
  signal W_43_27_i_5_n_0 : STD_LOGIC;
  signal W_43_27_i_6_n_0 : STD_LOGIC;
  signal W_43_27_i_7_n_0 : STD_LOGIC;
  signal W_43_27_i_8_n_0 : STD_LOGIC;
  signal W_43_27_i_9_n_0 : STD_LOGIC;
  signal W_43_31_i_10_n_0 : STD_LOGIC;
  signal W_43_31_i_11_n_0 : STD_LOGIC;
  signal W_43_31_i_12_n_0 : STD_LOGIC;
  signal W_43_31_i_13_n_0 : STD_LOGIC;
  signal W_43_31_i_14_n_0 : STD_LOGIC;
  signal W_43_31_i_15_n_0 : STD_LOGIC;
  signal W_43_31_i_17_n_0 : STD_LOGIC;
  signal W_43_31_i_19_n_0 : STD_LOGIC;
  signal W_43_31_i_2_n_0 : STD_LOGIC;
  signal W_43_31_i_3_n_0 : STD_LOGIC;
  signal W_43_31_i_4_n_0 : STD_LOGIC;
  signal W_43_31_i_5_n_0 : STD_LOGIC;
  signal W_43_31_i_6_n_0 : STD_LOGIC;
  signal W_43_31_i_7_n_0 : STD_LOGIC;
  signal W_43_31_i_8_n_0 : STD_LOGIC;
  signal W_43_31_i_9_n_0 : STD_LOGIC;
  signal W_43_3_i_10_n_0 : STD_LOGIC;
  signal W_43_3_i_11_n_0 : STD_LOGIC;
  signal W_43_3_i_15_n_0 : STD_LOGIC;
  signal W_43_3_i_2_n_0 : STD_LOGIC;
  signal W_43_3_i_3_n_0 : STD_LOGIC;
  signal W_43_3_i_4_n_0 : STD_LOGIC;
  signal W_43_3_i_5_n_0 : STD_LOGIC;
  signal W_43_3_i_6_n_0 : STD_LOGIC;
  signal W_43_3_i_7_n_0 : STD_LOGIC;
  signal W_43_3_i_8_n_0 : STD_LOGIC;
  signal W_43_3_i_9_n_0 : STD_LOGIC;
  signal W_43_7_i_10_n_0 : STD_LOGIC;
  signal W_43_7_i_11_n_0 : STD_LOGIC;
  signal W_43_7_i_12_n_0 : STD_LOGIC;
  signal W_43_7_i_13_n_0 : STD_LOGIC;
  signal W_43_7_i_14_n_0 : STD_LOGIC;
  signal W_43_7_i_15_n_0 : STD_LOGIC;
  signal W_43_7_i_16_n_0 : STD_LOGIC;
  signal W_43_7_i_17_n_0 : STD_LOGIC;
  signal W_43_7_i_2_n_0 : STD_LOGIC;
  signal W_43_7_i_3_n_0 : STD_LOGIC;
  signal W_43_7_i_4_n_0 : STD_LOGIC;
  signal W_43_7_i_5_n_0 : STD_LOGIC;
  signal W_43_7_i_6_n_0 : STD_LOGIC;
  signal W_43_7_i_7_n_0 : STD_LOGIC;
  signal W_43_7_i_8_n_0 : STD_LOGIC;
  signal W_43_7_i_9_n_0 : STD_LOGIC;
  signal W_44_11_i_10_n_0 : STD_LOGIC;
  signal W_44_11_i_11_n_0 : STD_LOGIC;
  signal W_44_11_i_12_n_0 : STD_LOGIC;
  signal W_44_11_i_13_n_0 : STD_LOGIC;
  signal W_44_11_i_14_n_0 : STD_LOGIC;
  signal W_44_11_i_15_n_0 : STD_LOGIC;
  signal W_44_11_i_16_n_0 : STD_LOGIC;
  signal W_44_11_i_17_n_0 : STD_LOGIC;
  signal W_44_11_i_2_n_0 : STD_LOGIC;
  signal W_44_11_i_3_n_0 : STD_LOGIC;
  signal W_44_11_i_4_n_0 : STD_LOGIC;
  signal W_44_11_i_5_n_0 : STD_LOGIC;
  signal W_44_11_i_6_n_0 : STD_LOGIC;
  signal W_44_11_i_7_n_0 : STD_LOGIC;
  signal W_44_11_i_8_n_0 : STD_LOGIC;
  signal W_44_11_i_9_n_0 : STD_LOGIC;
  signal W_44_15_i_10_n_0 : STD_LOGIC;
  signal W_44_15_i_11_n_0 : STD_LOGIC;
  signal W_44_15_i_12_n_0 : STD_LOGIC;
  signal W_44_15_i_13_n_0 : STD_LOGIC;
  signal W_44_15_i_14_n_0 : STD_LOGIC;
  signal W_44_15_i_15_n_0 : STD_LOGIC;
  signal W_44_15_i_16_n_0 : STD_LOGIC;
  signal W_44_15_i_17_n_0 : STD_LOGIC;
  signal W_44_15_i_2_n_0 : STD_LOGIC;
  signal W_44_15_i_3_n_0 : STD_LOGIC;
  signal W_44_15_i_4_n_0 : STD_LOGIC;
  signal W_44_15_i_5_n_0 : STD_LOGIC;
  signal W_44_15_i_6_n_0 : STD_LOGIC;
  signal W_44_15_i_7_n_0 : STD_LOGIC;
  signal W_44_15_i_8_n_0 : STD_LOGIC;
  signal W_44_15_i_9_n_0 : STD_LOGIC;
  signal W_44_19_i_10_n_0 : STD_LOGIC;
  signal W_44_19_i_11_n_0 : STD_LOGIC;
  signal W_44_19_i_12_n_0 : STD_LOGIC;
  signal W_44_19_i_13_n_0 : STD_LOGIC;
  signal W_44_19_i_14_n_0 : STD_LOGIC;
  signal W_44_19_i_15_n_0 : STD_LOGIC;
  signal W_44_19_i_16_n_0 : STD_LOGIC;
  signal W_44_19_i_17_n_0 : STD_LOGIC;
  signal W_44_19_i_2_n_0 : STD_LOGIC;
  signal W_44_19_i_3_n_0 : STD_LOGIC;
  signal W_44_19_i_4_n_0 : STD_LOGIC;
  signal W_44_19_i_5_n_0 : STD_LOGIC;
  signal W_44_19_i_6_n_0 : STD_LOGIC;
  signal W_44_19_i_7_n_0 : STD_LOGIC;
  signal W_44_19_i_8_n_0 : STD_LOGIC;
  signal W_44_19_i_9_n_0 : STD_LOGIC;
  signal W_44_23_i_10_n_0 : STD_LOGIC;
  signal W_44_23_i_11_n_0 : STD_LOGIC;
  signal W_44_23_i_12_n_0 : STD_LOGIC;
  signal W_44_23_i_13_n_0 : STD_LOGIC;
  signal W_44_23_i_14_n_0 : STD_LOGIC;
  signal W_44_23_i_15_n_0 : STD_LOGIC;
  signal W_44_23_i_16_n_0 : STD_LOGIC;
  signal W_44_23_i_17_n_0 : STD_LOGIC;
  signal W_44_23_i_2_n_0 : STD_LOGIC;
  signal W_44_23_i_3_n_0 : STD_LOGIC;
  signal W_44_23_i_4_n_0 : STD_LOGIC;
  signal W_44_23_i_5_n_0 : STD_LOGIC;
  signal W_44_23_i_6_n_0 : STD_LOGIC;
  signal W_44_23_i_7_n_0 : STD_LOGIC;
  signal W_44_23_i_8_n_0 : STD_LOGIC;
  signal W_44_23_i_9_n_0 : STD_LOGIC;
  signal W_44_27_i_10_n_0 : STD_LOGIC;
  signal W_44_27_i_11_n_0 : STD_LOGIC;
  signal W_44_27_i_12_n_0 : STD_LOGIC;
  signal W_44_27_i_13_n_0 : STD_LOGIC;
  signal W_44_27_i_14_n_0 : STD_LOGIC;
  signal W_44_27_i_15_n_0 : STD_LOGIC;
  signal W_44_27_i_16_n_0 : STD_LOGIC;
  signal W_44_27_i_17_n_0 : STD_LOGIC;
  signal W_44_27_i_2_n_0 : STD_LOGIC;
  signal W_44_27_i_3_n_0 : STD_LOGIC;
  signal W_44_27_i_4_n_0 : STD_LOGIC;
  signal W_44_27_i_5_n_0 : STD_LOGIC;
  signal W_44_27_i_6_n_0 : STD_LOGIC;
  signal W_44_27_i_7_n_0 : STD_LOGIC;
  signal W_44_27_i_8_n_0 : STD_LOGIC;
  signal W_44_27_i_9_n_0 : STD_LOGIC;
  signal W_44_31_i_10_n_0 : STD_LOGIC;
  signal W_44_31_i_11_n_0 : STD_LOGIC;
  signal W_44_31_i_12_n_0 : STD_LOGIC;
  signal W_44_31_i_13_n_0 : STD_LOGIC;
  signal W_44_31_i_14_n_0 : STD_LOGIC;
  signal W_44_31_i_15_n_0 : STD_LOGIC;
  signal W_44_31_i_17_n_0 : STD_LOGIC;
  signal W_44_31_i_19_n_0 : STD_LOGIC;
  signal W_44_31_i_2_n_0 : STD_LOGIC;
  signal W_44_31_i_3_n_0 : STD_LOGIC;
  signal W_44_31_i_4_n_0 : STD_LOGIC;
  signal W_44_31_i_5_n_0 : STD_LOGIC;
  signal W_44_31_i_6_n_0 : STD_LOGIC;
  signal W_44_31_i_7_n_0 : STD_LOGIC;
  signal W_44_31_i_8_n_0 : STD_LOGIC;
  signal W_44_31_i_9_n_0 : STD_LOGIC;
  signal W_44_3_i_10_n_0 : STD_LOGIC;
  signal W_44_3_i_11_n_0 : STD_LOGIC;
  signal W_44_3_i_15_n_0 : STD_LOGIC;
  signal W_44_3_i_2_n_0 : STD_LOGIC;
  signal W_44_3_i_3_n_0 : STD_LOGIC;
  signal W_44_3_i_4_n_0 : STD_LOGIC;
  signal W_44_3_i_5_n_0 : STD_LOGIC;
  signal W_44_3_i_6_n_0 : STD_LOGIC;
  signal W_44_3_i_7_n_0 : STD_LOGIC;
  signal W_44_3_i_8_n_0 : STD_LOGIC;
  signal W_44_3_i_9_n_0 : STD_LOGIC;
  signal W_44_7_i_10_n_0 : STD_LOGIC;
  signal W_44_7_i_11_n_0 : STD_LOGIC;
  signal W_44_7_i_12_n_0 : STD_LOGIC;
  signal W_44_7_i_13_n_0 : STD_LOGIC;
  signal W_44_7_i_14_n_0 : STD_LOGIC;
  signal W_44_7_i_15_n_0 : STD_LOGIC;
  signal W_44_7_i_16_n_0 : STD_LOGIC;
  signal W_44_7_i_17_n_0 : STD_LOGIC;
  signal W_44_7_i_2_n_0 : STD_LOGIC;
  signal W_44_7_i_3_n_0 : STD_LOGIC;
  signal W_44_7_i_4_n_0 : STD_LOGIC;
  signal W_44_7_i_5_n_0 : STD_LOGIC;
  signal W_44_7_i_6_n_0 : STD_LOGIC;
  signal W_44_7_i_7_n_0 : STD_LOGIC;
  signal W_44_7_i_8_n_0 : STD_LOGIC;
  signal W_44_7_i_9_n_0 : STD_LOGIC;
  signal W_45_11_i_10_n_0 : STD_LOGIC;
  signal W_45_11_i_11_n_0 : STD_LOGIC;
  signal W_45_11_i_12_n_0 : STD_LOGIC;
  signal W_45_11_i_13_n_0 : STD_LOGIC;
  signal W_45_11_i_14_n_0 : STD_LOGIC;
  signal W_45_11_i_15_n_0 : STD_LOGIC;
  signal W_45_11_i_16_n_0 : STD_LOGIC;
  signal W_45_11_i_17_n_0 : STD_LOGIC;
  signal W_45_11_i_2_n_0 : STD_LOGIC;
  signal W_45_11_i_3_n_0 : STD_LOGIC;
  signal W_45_11_i_4_n_0 : STD_LOGIC;
  signal W_45_11_i_5_n_0 : STD_LOGIC;
  signal W_45_11_i_6_n_0 : STD_LOGIC;
  signal W_45_11_i_7_n_0 : STD_LOGIC;
  signal W_45_11_i_8_n_0 : STD_LOGIC;
  signal W_45_11_i_9_n_0 : STD_LOGIC;
  signal W_45_15_i_10_n_0 : STD_LOGIC;
  signal W_45_15_i_11_n_0 : STD_LOGIC;
  signal W_45_15_i_12_n_0 : STD_LOGIC;
  signal W_45_15_i_13_n_0 : STD_LOGIC;
  signal W_45_15_i_14_n_0 : STD_LOGIC;
  signal W_45_15_i_15_n_0 : STD_LOGIC;
  signal W_45_15_i_16_n_0 : STD_LOGIC;
  signal W_45_15_i_17_n_0 : STD_LOGIC;
  signal W_45_15_i_2_n_0 : STD_LOGIC;
  signal W_45_15_i_3_n_0 : STD_LOGIC;
  signal W_45_15_i_4_n_0 : STD_LOGIC;
  signal W_45_15_i_5_n_0 : STD_LOGIC;
  signal W_45_15_i_6_n_0 : STD_LOGIC;
  signal W_45_15_i_7_n_0 : STD_LOGIC;
  signal W_45_15_i_8_n_0 : STD_LOGIC;
  signal W_45_15_i_9_n_0 : STD_LOGIC;
  signal W_45_19_i_10_n_0 : STD_LOGIC;
  signal W_45_19_i_11_n_0 : STD_LOGIC;
  signal W_45_19_i_12_n_0 : STD_LOGIC;
  signal W_45_19_i_13_n_0 : STD_LOGIC;
  signal W_45_19_i_14_n_0 : STD_LOGIC;
  signal W_45_19_i_15_n_0 : STD_LOGIC;
  signal W_45_19_i_16_n_0 : STD_LOGIC;
  signal W_45_19_i_17_n_0 : STD_LOGIC;
  signal W_45_19_i_2_n_0 : STD_LOGIC;
  signal W_45_19_i_3_n_0 : STD_LOGIC;
  signal W_45_19_i_4_n_0 : STD_LOGIC;
  signal W_45_19_i_5_n_0 : STD_LOGIC;
  signal W_45_19_i_6_n_0 : STD_LOGIC;
  signal W_45_19_i_7_n_0 : STD_LOGIC;
  signal W_45_19_i_8_n_0 : STD_LOGIC;
  signal W_45_19_i_9_n_0 : STD_LOGIC;
  signal W_45_23_i_10_n_0 : STD_LOGIC;
  signal W_45_23_i_11_n_0 : STD_LOGIC;
  signal W_45_23_i_12_n_0 : STD_LOGIC;
  signal W_45_23_i_13_n_0 : STD_LOGIC;
  signal W_45_23_i_14_n_0 : STD_LOGIC;
  signal W_45_23_i_15_n_0 : STD_LOGIC;
  signal W_45_23_i_16_n_0 : STD_LOGIC;
  signal W_45_23_i_17_n_0 : STD_LOGIC;
  signal W_45_23_i_2_n_0 : STD_LOGIC;
  signal W_45_23_i_3_n_0 : STD_LOGIC;
  signal W_45_23_i_4_n_0 : STD_LOGIC;
  signal W_45_23_i_5_n_0 : STD_LOGIC;
  signal W_45_23_i_6_n_0 : STD_LOGIC;
  signal W_45_23_i_7_n_0 : STD_LOGIC;
  signal W_45_23_i_8_n_0 : STD_LOGIC;
  signal W_45_23_i_9_n_0 : STD_LOGIC;
  signal W_45_27_i_10_n_0 : STD_LOGIC;
  signal W_45_27_i_11_n_0 : STD_LOGIC;
  signal W_45_27_i_12_n_0 : STD_LOGIC;
  signal W_45_27_i_13_n_0 : STD_LOGIC;
  signal W_45_27_i_14_n_0 : STD_LOGIC;
  signal W_45_27_i_15_n_0 : STD_LOGIC;
  signal W_45_27_i_16_n_0 : STD_LOGIC;
  signal W_45_27_i_17_n_0 : STD_LOGIC;
  signal W_45_27_i_2_n_0 : STD_LOGIC;
  signal W_45_27_i_3_n_0 : STD_LOGIC;
  signal W_45_27_i_4_n_0 : STD_LOGIC;
  signal W_45_27_i_5_n_0 : STD_LOGIC;
  signal W_45_27_i_6_n_0 : STD_LOGIC;
  signal W_45_27_i_7_n_0 : STD_LOGIC;
  signal W_45_27_i_8_n_0 : STD_LOGIC;
  signal W_45_27_i_9_n_0 : STD_LOGIC;
  signal W_45_31_i_10_n_0 : STD_LOGIC;
  signal W_45_31_i_11_n_0 : STD_LOGIC;
  signal W_45_31_i_12_n_0 : STD_LOGIC;
  signal W_45_31_i_13_n_0 : STD_LOGIC;
  signal W_45_31_i_14_n_0 : STD_LOGIC;
  signal W_45_31_i_15_n_0 : STD_LOGIC;
  signal W_45_31_i_17_n_0 : STD_LOGIC;
  signal W_45_31_i_19_n_0 : STD_LOGIC;
  signal W_45_31_i_2_n_0 : STD_LOGIC;
  signal W_45_31_i_3_n_0 : STD_LOGIC;
  signal W_45_31_i_4_n_0 : STD_LOGIC;
  signal W_45_31_i_5_n_0 : STD_LOGIC;
  signal W_45_31_i_6_n_0 : STD_LOGIC;
  signal W_45_31_i_7_n_0 : STD_LOGIC;
  signal W_45_31_i_8_n_0 : STD_LOGIC;
  signal W_45_31_i_9_n_0 : STD_LOGIC;
  signal W_45_3_i_10_n_0 : STD_LOGIC;
  signal W_45_3_i_11_n_0 : STD_LOGIC;
  signal W_45_3_i_15_n_0 : STD_LOGIC;
  signal W_45_3_i_2_n_0 : STD_LOGIC;
  signal W_45_3_i_3_n_0 : STD_LOGIC;
  signal W_45_3_i_4_n_0 : STD_LOGIC;
  signal W_45_3_i_5_n_0 : STD_LOGIC;
  signal W_45_3_i_6_n_0 : STD_LOGIC;
  signal W_45_3_i_7_n_0 : STD_LOGIC;
  signal W_45_3_i_8_n_0 : STD_LOGIC;
  signal W_45_3_i_9_n_0 : STD_LOGIC;
  signal W_45_7_i_10_n_0 : STD_LOGIC;
  signal W_45_7_i_11_n_0 : STD_LOGIC;
  signal W_45_7_i_12_n_0 : STD_LOGIC;
  signal W_45_7_i_13_n_0 : STD_LOGIC;
  signal W_45_7_i_14_n_0 : STD_LOGIC;
  signal W_45_7_i_15_n_0 : STD_LOGIC;
  signal W_45_7_i_16_n_0 : STD_LOGIC;
  signal W_45_7_i_17_n_0 : STD_LOGIC;
  signal W_45_7_i_2_n_0 : STD_LOGIC;
  signal W_45_7_i_3_n_0 : STD_LOGIC;
  signal W_45_7_i_4_n_0 : STD_LOGIC;
  signal W_45_7_i_5_n_0 : STD_LOGIC;
  signal W_45_7_i_6_n_0 : STD_LOGIC;
  signal W_45_7_i_7_n_0 : STD_LOGIC;
  signal W_45_7_i_8_n_0 : STD_LOGIC;
  signal W_45_7_i_9_n_0 : STD_LOGIC;
  signal W_46_11_i_10_n_0 : STD_LOGIC;
  signal W_46_11_i_11_n_0 : STD_LOGIC;
  signal W_46_11_i_12_n_0 : STD_LOGIC;
  signal W_46_11_i_13_n_0 : STD_LOGIC;
  signal W_46_11_i_14_n_0 : STD_LOGIC;
  signal W_46_11_i_15_n_0 : STD_LOGIC;
  signal W_46_11_i_16_n_0 : STD_LOGIC;
  signal W_46_11_i_17_n_0 : STD_LOGIC;
  signal W_46_11_i_2_n_0 : STD_LOGIC;
  signal W_46_11_i_3_n_0 : STD_LOGIC;
  signal W_46_11_i_4_n_0 : STD_LOGIC;
  signal W_46_11_i_5_n_0 : STD_LOGIC;
  signal W_46_11_i_6_n_0 : STD_LOGIC;
  signal W_46_11_i_7_n_0 : STD_LOGIC;
  signal W_46_11_i_8_n_0 : STD_LOGIC;
  signal W_46_11_i_9_n_0 : STD_LOGIC;
  signal W_46_15_i_10_n_0 : STD_LOGIC;
  signal W_46_15_i_11_n_0 : STD_LOGIC;
  signal W_46_15_i_12_n_0 : STD_LOGIC;
  signal W_46_15_i_13_n_0 : STD_LOGIC;
  signal W_46_15_i_14_n_0 : STD_LOGIC;
  signal W_46_15_i_15_n_0 : STD_LOGIC;
  signal W_46_15_i_16_n_0 : STD_LOGIC;
  signal W_46_15_i_17_n_0 : STD_LOGIC;
  signal W_46_15_i_2_n_0 : STD_LOGIC;
  signal W_46_15_i_3_n_0 : STD_LOGIC;
  signal W_46_15_i_4_n_0 : STD_LOGIC;
  signal W_46_15_i_5_n_0 : STD_LOGIC;
  signal W_46_15_i_6_n_0 : STD_LOGIC;
  signal W_46_15_i_7_n_0 : STD_LOGIC;
  signal W_46_15_i_8_n_0 : STD_LOGIC;
  signal W_46_15_i_9_n_0 : STD_LOGIC;
  signal W_46_19_i_10_n_0 : STD_LOGIC;
  signal W_46_19_i_11_n_0 : STD_LOGIC;
  signal W_46_19_i_12_n_0 : STD_LOGIC;
  signal W_46_19_i_13_n_0 : STD_LOGIC;
  signal W_46_19_i_14_n_0 : STD_LOGIC;
  signal W_46_19_i_15_n_0 : STD_LOGIC;
  signal W_46_19_i_16_n_0 : STD_LOGIC;
  signal W_46_19_i_17_n_0 : STD_LOGIC;
  signal W_46_19_i_2_n_0 : STD_LOGIC;
  signal W_46_19_i_3_n_0 : STD_LOGIC;
  signal W_46_19_i_4_n_0 : STD_LOGIC;
  signal W_46_19_i_5_n_0 : STD_LOGIC;
  signal W_46_19_i_6_n_0 : STD_LOGIC;
  signal W_46_19_i_7_n_0 : STD_LOGIC;
  signal W_46_19_i_8_n_0 : STD_LOGIC;
  signal W_46_19_i_9_n_0 : STD_LOGIC;
  signal W_46_23_i_10_n_0 : STD_LOGIC;
  signal W_46_23_i_11_n_0 : STD_LOGIC;
  signal W_46_23_i_12_n_0 : STD_LOGIC;
  signal W_46_23_i_13_n_0 : STD_LOGIC;
  signal W_46_23_i_14_n_0 : STD_LOGIC;
  signal W_46_23_i_15_n_0 : STD_LOGIC;
  signal W_46_23_i_16_n_0 : STD_LOGIC;
  signal W_46_23_i_17_n_0 : STD_LOGIC;
  signal W_46_23_i_2_n_0 : STD_LOGIC;
  signal W_46_23_i_3_n_0 : STD_LOGIC;
  signal W_46_23_i_4_n_0 : STD_LOGIC;
  signal W_46_23_i_5_n_0 : STD_LOGIC;
  signal W_46_23_i_6_n_0 : STD_LOGIC;
  signal W_46_23_i_7_n_0 : STD_LOGIC;
  signal W_46_23_i_8_n_0 : STD_LOGIC;
  signal W_46_23_i_9_n_0 : STD_LOGIC;
  signal W_46_27_i_10_n_0 : STD_LOGIC;
  signal W_46_27_i_11_n_0 : STD_LOGIC;
  signal W_46_27_i_12_n_0 : STD_LOGIC;
  signal W_46_27_i_13_n_0 : STD_LOGIC;
  signal W_46_27_i_14_n_0 : STD_LOGIC;
  signal W_46_27_i_15_n_0 : STD_LOGIC;
  signal W_46_27_i_16_n_0 : STD_LOGIC;
  signal W_46_27_i_17_n_0 : STD_LOGIC;
  signal W_46_27_i_2_n_0 : STD_LOGIC;
  signal W_46_27_i_3_n_0 : STD_LOGIC;
  signal W_46_27_i_4_n_0 : STD_LOGIC;
  signal W_46_27_i_5_n_0 : STD_LOGIC;
  signal W_46_27_i_6_n_0 : STD_LOGIC;
  signal W_46_27_i_7_n_0 : STD_LOGIC;
  signal W_46_27_i_8_n_0 : STD_LOGIC;
  signal W_46_27_i_9_n_0 : STD_LOGIC;
  signal W_46_31_i_10_n_0 : STD_LOGIC;
  signal W_46_31_i_11_n_0 : STD_LOGIC;
  signal W_46_31_i_12_n_0 : STD_LOGIC;
  signal W_46_31_i_13_n_0 : STD_LOGIC;
  signal W_46_31_i_14_n_0 : STD_LOGIC;
  signal W_46_31_i_15_n_0 : STD_LOGIC;
  signal W_46_31_i_17_n_0 : STD_LOGIC;
  signal W_46_31_i_19_n_0 : STD_LOGIC;
  signal W_46_31_i_2_n_0 : STD_LOGIC;
  signal W_46_31_i_3_n_0 : STD_LOGIC;
  signal W_46_31_i_4_n_0 : STD_LOGIC;
  signal W_46_31_i_5_n_0 : STD_LOGIC;
  signal W_46_31_i_6_n_0 : STD_LOGIC;
  signal W_46_31_i_7_n_0 : STD_LOGIC;
  signal W_46_31_i_8_n_0 : STD_LOGIC;
  signal W_46_31_i_9_n_0 : STD_LOGIC;
  signal W_46_3_i_10_n_0 : STD_LOGIC;
  signal W_46_3_i_11_n_0 : STD_LOGIC;
  signal W_46_3_i_15_n_0 : STD_LOGIC;
  signal W_46_3_i_2_n_0 : STD_LOGIC;
  signal W_46_3_i_3_n_0 : STD_LOGIC;
  signal W_46_3_i_4_n_0 : STD_LOGIC;
  signal W_46_3_i_5_n_0 : STD_LOGIC;
  signal W_46_3_i_6_n_0 : STD_LOGIC;
  signal W_46_3_i_7_n_0 : STD_LOGIC;
  signal W_46_3_i_8_n_0 : STD_LOGIC;
  signal W_46_3_i_9_n_0 : STD_LOGIC;
  signal W_46_7_i_10_n_0 : STD_LOGIC;
  signal W_46_7_i_11_n_0 : STD_LOGIC;
  signal W_46_7_i_12_n_0 : STD_LOGIC;
  signal W_46_7_i_13_n_0 : STD_LOGIC;
  signal W_46_7_i_14_n_0 : STD_LOGIC;
  signal W_46_7_i_15_n_0 : STD_LOGIC;
  signal W_46_7_i_16_n_0 : STD_LOGIC;
  signal W_46_7_i_17_n_0 : STD_LOGIC;
  signal W_46_7_i_2_n_0 : STD_LOGIC;
  signal W_46_7_i_3_n_0 : STD_LOGIC;
  signal W_46_7_i_4_n_0 : STD_LOGIC;
  signal W_46_7_i_5_n_0 : STD_LOGIC;
  signal W_46_7_i_6_n_0 : STD_LOGIC;
  signal W_46_7_i_7_n_0 : STD_LOGIC;
  signal W_46_7_i_8_n_0 : STD_LOGIC;
  signal W_46_7_i_9_n_0 : STD_LOGIC;
  signal W_47_11_i_10_n_0 : STD_LOGIC;
  signal W_47_11_i_11_n_0 : STD_LOGIC;
  signal W_47_11_i_12_n_0 : STD_LOGIC;
  signal W_47_11_i_13_n_0 : STD_LOGIC;
  signal W_47_11_i_14_n_0 : STD_LOGIC;
  signal W_47_11_i_15_n_0 : STD_LOGIC;
  signal W_47_11_i_16_n_0 : STD_LOGIC;
  signal W_47_11_i_17_n_0 : STD_LOGIC;
  signal W_47_11_i_2_n_0 : STD_LOGIC;
  signal W_47_11_i_3_n_0 : STD_LOGIC;
  signal W_47_11_i_4_n_0 : STD_LOGIC;
  signal W_47_11_i_5_n_0 : STD_LOGIC;
  signal W_47_11_i_6_n_0 : STD_LOGIC;
  signal W_47_11_i_7_n_0 : STD_LOGIC;
  signal W_47_11_i_8_n_0 : STD_LOGIC;
  signal W_47_11_i_9_n_0 : STD_LOGIC;
  signal W_47_15_i_10_n_0 : STD_LOGIC;
  signal W_47_15_i_11_n_0 : STD_LOGIC;
  signal W_47_15_i_12_n_0 : STD_LOGIC;
  signal W_47_15_i_13_n_0 : STD_LOGIC;
  signal W_47_15_i_14_n_0 : STD_LOGIC;
  signal W_47_15_i_15_n_0 : STD_LOGIC;
  signal W_47_15_i_16_n_0 : STD_LOGIC;
  signal W_47_15_i_17_n_0 : STD_LOGIC;
  signal W_47_15_i_2_n_0 : STD_LOGIC;
  signal W_47_15_i_3_n_0 : STD_LOGIC;
  signal W_47_15_i_4_n_0 : STD_LOGIC;
  signal W_47_15_i_5_n_0 : STD_LOGIC;
  signal W_47_15_i_6_n_0 : STD_LOGIC;
  signal W_47_15_i_7_n_0 : STD_LOGIC;
  signal W_47_15_i_8_n_0 : STD_LOGIC;
  signal W_47_15_i_9_n_0 : STD_LOGIC;
  signal W_47_19_i_10_n_0 : STD_LOGIC;
  signal W_47_19_i_11_n_0 : STD_LOGIC;
  signal W_47_19_i_12_n_0 : STD_LOGIC;
  signal W_47_19_i_13_n_0 : STD_LOGIC;
  signal W_47_19_i_14_n_0 : STD_LOGIC;
  signal W_47_19_i_15_n_0 : STD_LOGIC;
  signal W_47_19_i_16_n_0 : STD_LOGIC;
  signal W_47_19_i_17_n_0 : STD_LOGIC;
  signal W_47_19_i_2_n_0 : STD_LOGIC;
  signal W_47_19_i_3_n_0 : STD_LOGIC;
  signal W_47_19_i_4_n_0 : STD_LOGIC;
  signal W_47_19_i_5_n_0 : STD_LOGIC;
  signal W_47_19_i_6_n_0 : STD_LOGIC;
  signal W_47_19_i_7_n_0 : STD_LOGIC;
  signal W_47_19_i_8_n_0 : STD_LOGIC;
  signal W_47_19_i_9_n_0 : STD_LOGIC;
  signal W_47_23_i_10_n_0 : STD_LOGIC;
  signal W_47_23_i_11_n_0 : STD_LOGIC;
  signal W_47_23_i_12_n_0 : STD_LOGIC;
  signal W_47_23_i_13_n_0 : STD_LOGIC;
  signal W_47_23_i_14_n_0 : STD_LOGIC;
  signal W_47_23_i_15_n_0 : STD_LOGIC;
  signal W_47_23_i_16_n_0 : STD_LOGIC;
  signal W_47_23_i_17_n_0 : STD_LOGIC;
  signal W_47_23_i_2_n_0 : STD_LOGIC;
  signal W_47_23_i_3_n_0 : STD_LOGIC;
  signal W_47_23_i_4_n_0 : STD_LOGIC;
  signal W_47_23_i_5_n_0 : STD_LOGIC;
  signal W_47_23_i_6_n_0 : STD_LOGIC;
  signal W_47_23_i_7_n_0 : STD_LOGIC;
  signal W_47_23_i_8_n_0 : STD_LOGIC;
  signal W_47_23_i_9_n_0 : STD_LOGIC;
  signal W_47_27_i_10_n_0 : STD_LOGIC;
  signal W_47_27_i_11_n_0 : STD_LOGIC;
  signal W_47_27_i_12_n_0 : STD_LOGIC;
  signal W_47_27_i_13_n_0 : STD_LOGIC;
  signal W_47_27_i_14_n_0 : STD_LOGIC;
  signal W_47_27_i_15_n_0 : STD_LOGIC;
  signal W_47_27_i_16_n_0 : STD_LOGIC;
  signal W_47_27_i_17_n_0 : STD_LOGIC;
  signal W_47_27_i_2_n_0 : STD_LOGIC;
  signal W_47_27_i_3_n_0 : STD_LOGIC;
  signal W_47_27_i_4_n_0 : STD_LOGIC;
  signal W_47_27_i_5_n_0 : STD_LOGIC;
  signal W_47_27_i_6_n_0 : STD_LOGIC;
  signal W_47_27_i_7_n_0 : STD_LOGIC;
  signal W_47_27_i_8_n_0 : STD_LOGIC;
  signal W_47_27_i_9_n_0 : STD_LOGIC;
  signal W_47_31_i_10_n_0 : STD_LOGIC;
  signal W_47_31_i_11_n_0 : STD_LOGIC;
  signal W_47_31_i_12_n_0 : STD_LOGIC;
  signal W_47_31_i_13_n_0 : STD_LOGIC;
  signal W_47_31_i_14_n_0 : STD_LOGIC;
  signal W_47_31_i_15_n_0 : STD_LOGIC;
  signal W_47_31_i_17_n_0 : STD_LOGIC;
  signal W_47_31_i_19_n_0 : STD_LOGIC;
  signal W_47_31_i_2_n_0 : STD_LOGIC;
  signal W_47_31_i_3_n_0 : STD_LOGIC;
  signal W_47_31_i_4_n_0 : STD_LOGIC;
  signal W_47_31_i_5_n_0 : STD_LOGIC;
  signal W_47_31_i_6_n_0 : STD_LOGIC;
  signal W_47_31_i_7_n_0 : STD_LOGIC;
  signal W_47_31_i_8_n_0 : STD_LOGIC;
  signal W_47_31_i_9_n_0 : STD_LOGIC;
  signal W_47_3_i_10_n_0 : STD_LOGIC;
  signal W_47_3_i_11_n_0 : STD_LOGIC;
  signal W_47_3_i_15_n_0 : STD_LOGIC;
  signal W_47_3_i_2_n_0 : STD_LOGIC;
  signal W_47_3_i_3_n_0 : STD_LOGIC;
  signal W_47_3_i_4_n_0 : STD_LOGIC;
  signal W_47_3_i_5_n_0 : STD_LOGIC;
  signal W_47_3_i_6_n_0 : STD_LOGIC;
  signal W_47_3_i_7_n_0 : STD_LOGIC;
  signal W_47_3_i_8_n_0 : STD_LOGIC;
  signal W_47_3_i_9_n_0 : STD_LOGIC;
  signal W_47_7_i_10_n_0 : STD_LOGIC;
  signal W_47_7_i_11_n_0 : STD_LOGIC;
  signal W_47_7_i_12_n_0 : STD_LOGIC;
  signal W_47_7_i_13_n_0 : STD_LOGIC;
  signal W_47_7_i_14_n_0 : STD_LOGIC;
  signal W_47_7_i_15_n_0 : STD_LOGIC;
  signal W_47_7_i_16_n_0 : STD_LOGIC;
  signal W_47_7_i_17_n_0 : STD_LOGIC;
  signal W_47_7_i_2_n_0 : STD_LOGIC;
  signal W_47_7_i_3_n_0 : STD_LOGIC;
  signal W_47_7_i_4_n_0 : STD_LOGIC;
  signal W_47_7_i_5_n_0 : STD_LOGIC;
  signal W_47_7_i_6_n_0 : STD_LOGIC;
  signal W_47_7_i_7_n_0 : STD_LOGIC;
  signal W_47_7_i_8_n_0 : STD_LOGIC;
  signal W_47_7_i_9_n_0 : STD_LOGIC;
  signal W_48 : STD_LOGIC;
  signal W_48_11_i_10_n_0 : STD_LOGIC;
  signal W_48_11_i_11_n_0 : STD_LOGIC;
  signal W_48_11_i_12_n_0 : STD_LOGIC;
  signal W_48_11_i_13_n_0 : STD_LOGIC;
  signal W_48_11_i_14_n_0 : STD_LOGIC;
  signal W_48_11_i_15_n_0 : STD_LOGIC;
  signal W_48_11_i_16_n_0 : STD_LOGIC;
  signal W_48_11_i_17_n_0 : STD_LOGIC;
  signal W_48_11_i_2_n_0 : STD_LOGIC;
  signal W_48_11_i_3_n_0 : STD_LOGIC;
  signal W_48_11_i_4_n_0 : STD_LOGIC;
  signal W_48_11_i_5_n_0 : STD_LOGIC;
  signal W_48_11_i_6_n_0 : STD_LOGIC;
  signal W_48_11_i_7_n_0 : STD_LOGIC;
  signal W_48_11_i_8_n_0 : STD_LOGIC;
  signal W_48_11_i_9_n_0 : STD_LOGIC;
  signal W_48_15_i_10_n_0 : STD_LOGIC;
  signal W_48_15_i_11_n_0 : STD_LOGIC;
  signal W_48_15_i_12_n_0 : STD_LOGIC;
  signal W_48_15_i_13_n_0 : STD_LOGIC;
  signal W_48_15_i_14_n_0 : STD_LOGIC;
  signal W_48_15_i_15_n_0 : STD_LOGIC;
  signal W_48_15_i_16_n_0 : STD_LOGIC;
  signal W_48_15_i_17_n_0 : STD_LOGIC;
  signal W_48_15_i_2_n_0 : STD_LOGIC;
  signal W_48_15_i_3_n_0 : STD_LOGIC;
  signal W_48_15_i_4_n_0 : STD_LOGIC;
  signal W_48_15_i_5_n_0 : STD_LOGIC;
  signal W_48_15_i_6_n_0 : STD_LOGIC;
  signal W_48_15_i_7_n_0 : STD_LOGIC;
  signal W_48_15_i_8_n_0 : STD_LOGIC;
  signal W_48_15_i_9_n_0 : STD_LOGIC;
  signal W_48_19_i_10_n_0 : STD_LOGIC;
  signal W_48_19_i_11_n_0 : STD_LOGIC;
  signal W_48_19_i_12_n_0 : STD_LOGIC;
  signal W_48_19_i_13_n_0 : STD_LOGIC;
  signal W_48_19_i_14_n_0 : STD_LOGIC;
  signal W_48_19_i_15_n_0 : STD_LOGIC;
  signal W_48_19_i_16_n_0 : STD_LOGIC;
  signal W_48_19_i_17_n_0 : STD_LOGIC;
  signal W_48_19_i_2_n_0 : STD_LOGIC;
  signal W_48_19_i_3_n_0 : STD_LOGIC;
  signal W_48_19_i_4_n_0 : STD_LOGIC;
  signal W_48_19_i_5_n_0 : STD_LOGIC;
  signal W_48_19_i_6_n_0 : STD_LOGIC;
  signal W_48_19_i_7_n_0 : STD_LOGIC;
  signal W_48_19_i_8_n_0 : STD_LOGIC;
  signal W_48_19_i_9_n_0 : STD_LOGIC;
  signal W_48_23_i_10_n_0 : STD_LOGIC;
  signal W_48_23_i_11_n_0 : STD_LOGIC;
  signal W_48_23_i_12_n_0 : STD_LOGIC;
  signal W_48_23_i_13_n_0 : STD_LOGIC;
  signal W_48_23_i_14_n_0 : STD_LOGIC;
  signal W_48_23_i_15_n_0 : STD_LOGIC;
  signal W_48_23_i_16_n_0 : STD_LOGIC;
  signal W_48_23_i_17_n_0 : STD_LOGIC;
  signal W_48_23_i_2_n_0 : STD_LOGIC;
  signal W_48_23_i_3_n_0 : STD_LOGIC;
  signal W_48_23_i_4_n_0 : STD_LOGIC;
  signal W_48_23_i_5_n_0 : STD_LOGIC;
  signal W_48_23_i_6_n_0 : STD_LOGIC;
  signal W_48_23_i_7_n_0 : STD_LOGIC;
  signal W_48_23_i_8_n_0 : STD_LOGIC;
  signal W_48_23_i_9_n_0 : STD_LOGIC;
  signal W_48_27_i_10_n_0 : STD_LOGIC;
  signal W_48_27_i_11_n_0 : STD_LOGIC;
  signal W_48_27_i_12_n_0 : STD_LOGIC;
  signal W_48_27_i_13_n_0 : STD_LOGIC;
  signal W_48_27_i_14_n_0 : STD_LOGIC;
  signal W_48_27_i_15_n_0 : STD_LOGIC;
  signal W_48_27_i_16_n_0 : STD_LOGIC;
  signal W_48_27_i_17_n_0 : STD_LOGIC;
  signal W_48_27_i_2_n_0 : STD_LOGIC;
  signal W_48_27_i_3_n_0 : STD_LOGIC;
  signal W_48_27_i_4_n_0 : STD_LOGIC;
  signal W_48_27_i_5_n_0 : STD_LOGIC;
  signal W_48_27_i_6_n_0 : STD_LOGIC;
  signal W_48_27_i_7_n_0 : STD_LOGIC;
  signal W_48_27_i_8_n_0 : STD_LOGIC;
  signal W_48_27_i_9_n_0 : STD_LOGIC;
  signal W_48_31_i_10_n_0 : STD_LOGIC;
  signal W_48_31_i_11_n_0 : STD_LOGIC;
  signal W_48_31_i_12_n_0 : STD_LOGIC;
  signal W_48_31_i_13_n_0 : STD_LOGIC;
  signal W_48_31_i_14_n_0 : STD_LOGIC;
  signal W_48_31_i_15_n_0 : STD_LOGIC;
  signal W_48_31_i_16_n_0 : STD_LOGIC;
  signal W_48_31_i_18_n_0 : STD_LOGIC;
  signal W_48_31_i_20_n_0 : STD_LOGIC;
  signal W_48_31_i_3_n_0 : STD_LOGIC;
  signal W_48_31_i_4_n_0 : STD_LOGIC;
  signal W_48_31_i_5_n_0 : STD_LOGIC;
  signal W_48_31_i_6_n_0 : STD_LOGIC;
  signal W_48_31_i_7_n_0 : STD_LOGIC;
  signal W_48_31_i_8_n_0 : STD_LOGIC;
  signal W_48_31_i_9_n_0 : STD_LOGIC;
  signal W_48_3_i_10_n_0 : STD_LOGIC;
  signal W_48_3_i_11_n_0 : STD_LOGIC;
  signal W_48_3_i_15_n_0 : STD_LOGIC;
  signal W_48_3_i_2_n_0 : STD_LOGIC;
  signal W_48_3_i_3_n_0 : STD_LOGIC;
  signal W_48_3_i_4_n_0 : STD_LOGIC;
  signal W_48_3_i_5_n_0 : STD_LOGIC;
  signal W_48_3_i_6_n_0 : STD_LOGIC;
  signal W_48_3_i_7_n_0 : STD_LOGIC;
  signal W_48_3_i_8_n_0 : STD_LOGIC;
  signal W_48_3_i_9_n_0 : STD_LOGIC;
  signal W_48_7_i_10_n_0 : STD_LOGIC;
  signal W_48_7_i_11_n_0 : STD_LOGIC;
  signal W_48_7_i_12_n_0 : STD_LOGIC;
  signal W_48_7_i_13_n_0 : STD_LOGIC;
  signal W_48_7_i_14_n_0 : STD_LOGIC;
  signal W_48_7_i_15_n_0 : STD_LOGIC;
  signal W_48_7_i_16_n_0 : STD_LOGIC;
  signal W_48_7_i_17_n_0 : STD_LOGIC;
  signal W_48_7_i_2_n_0 : STD_LOGIC;
  signal W_48_7_i_3_n_0 : STD_LOGIC;
  signal W_48_7_i_4_n_0 : STD_LOGIC;
  signal W_48_7_i_5_n_0 : STD_LOGIC;
  signal W_48_7_i_6_n_0 : STD_LOGIC;
  signal W_48_7_i_7_n_0 : STD_LOGIC;
  signal W_48_7_i_8_n_0 : STD_LOGIC;
  signal W_48_7_i_9_n_0 : STD_LOGIC;
  signal W_49_11_i_10_n_0 : STD_LOGIC;
  signal W_49_11_i_11_n_0 : STD_LOGIC;
  signal W_49_11_i_12_n_0 : STD_LOGIC;
  signal W_49_11_i_13_n_0 : STD_LOGIC;
  signal W_49_11_i_14_n_0 : STD_LOGIC;
  signal W_49_11_i_15_n_0 : STD_LOGIC;
  signal W_49_11_i_16_n_0 : STD_LOGIC;
  signal W_49_11_i_17_n_0 : STD_LOGIC;
  signal W_49_11_i_2_n_0 : STD_LOGIC;
  signal W_49_11_i_3_n_0 : STD_LOGIC;
  signal W_49_11_i_4_n_0 : STD_LOGIC;
  signal W_49_11_i_5_n_0 : STD_LOGIC;
  signal W_49_11_i_6_n_0 : STD_LOGIC;
  signal W_49_11_i_7_n_0 : STD_LOGIC;
  signal W_49_11_i_8_n_0 : STD_LOGIC;
  signal W_49_11_i_9_n_0 : STD_LOGIC;
  signal W_49_15_i_10_n_0 : STD_LOGIC;
  signal W_49_15_i_11_n_0 : STD_LOGIC;
  signal W_49_15_i_12_n_0 : STD_LOGIC;
  signal W_49_15_i_13_n_0 : STD_LOGIC;
  signal W_49_15_i_14_n_0 : STD_LOGIC;
  signal W_49_15_i_15_n_0 : STD_LOGIC;
  signal W_49_15_i_16_n_0 : STD_LOGIC;
  signal W_49_15_i_17_n_0 : STD_LOGIC;
  signal W_49_15_i_2_n_0 : STD_LOGIC;
  signal W_49_15_i_3_n_0 : STD_LOGIC;
  signal W_49_15_i_4_n_0 : STD_LOGIC;
  signal W_49_15_i_5_n_0 : STD_LOGIC;
  signal W_49_15_i_6_n_0 : STD_LOGIC;
  signal W_49_15_i_7_n_0 : STD_LOGIC;
  signal W_49_15_i_8_n_0 : STD_LOGIC;
  signal W_49_15_i_9_n_0 : STD_LOGIC;
  signal W_49_19_i_10_n_0 : STD_LOGIC;
  signal W_49_19_i_11_n_0 : STD_LOGIC;
  signal W_49_19_i_12_n_0 : STD_LOGIC;
  signal W_49_19_i_13_n_0 : STD_LOGIC;
  signal W_49_19_i_14_n_0 : STD_LOGIC;
  signal W_49_19_i_15_n_0 : STD_LOGIC;
  signal W_49_19_i_16_n_0 : STD_LOGIC;
  signal W_49_19_i_17_n_0 : STD_LOGIC;
  signal W_49_19_i_2_n_0 : STD_LOGIC;
  signal W_49_19_i_3_n_0 : STD_LOGIC;
  signal W_49_19_i_4_n_0 : STD_LOGIC;
  signal W_49_19_i_5_n_0 : STD_LOGIC;
  signal W_49_19_i_6_n_0 : STD_LOGIC;
  signal W_49_19_i_7_n_0 : STD_LOGIC;
  signal W_49_19_i_8_n_0 : STD_LOGIC;
  signal W_49_19_i_9_n_0 : STD_LOGIC;
  signal W_49_23_i_10_n_0 : STD_LOGIC;
  signal W_49_23_i_11_n_0 : STD_LOGIC;
  signal W_49_23_i_12_n_0 : STD_LOGIC;
  signal W_49_23_i_13_n_0 : STD_LOGIC;
  signal W_49_23_i_14_n_0 : STD_LOGIC;
  signal W_49_23_i_15_n_0 : STD_LOGIC;
  signal W_49_23_i_16_n_0 : STD_LOGIC;
  signal W_49_23_i_17_n_0 : STD_LOGIC;
  signal W_49_23_i_2_n_0 : STD_LOGIC;
  signal W_49_23_i_3_n_0 : STD_LOGIC;
  signal W_49_23_i_4_n_0 : STD_LOGIC;
  signal W_49_23_i_5_n_0 : STD_LOGIC;
  signal W_49_23_i_6_n_0 : STD_LOGIC;
  signal W_49_23_i_7_n_0 : STD_LOGIC;
  signal W_49_23_i_8_n_0 : STD_LOGIC;
  signal W_49_23_i_9_n_0 : STD_LOGIC;
  signal W_49_27_i_10_n_0 : STD_LOGIC;
  signal W_49_27_i_11_n_0 : STD_LOGIC;
  signal W_49_27_i_12_n_0 : STD_LOGIC;
  signal W_49_27_i_13_n_0 : STD_LOGIC;
  signal W_49_27_i_14_n_0 : STD_LOGIC;
  signal W_49_27_i_15_n_0 : STD_LOGIC;
  signal W_49_27_i_16_n_0 : STD_LOGIC;
  signal W_49_27_i_17_n_0 : STD_LOGIC;
  signal W_49_27_i_2_n_0 : STD_LOGIC;
  signal W_49_27_i_3_n_0 : STD_LOGIC;
  signal W_49_27_i_4_n_0 : STD_LOGIC;
  signal W_49_27_i_5_n_0 : STD_LOGIC;
  signal W_49_27_i_6_n_0 : STD_LOGIC;
  signal W_49_27_i_7_n_0 : STD_LOGIC;
  signal W_49_27_i_8_n_0 : STD_LOGIC;
  signal W_49_27_i_9_n_0 : STD_LOGIC;
  signal W_49_31_i_10_n_0 : STD_LOGIC;
  signal W_49_31_i_11_n_0 : STD_LOGIC;
  signal W_49_31_i_12_n_0 : STD_LOGIC;
  signal W_49_31_i_13_n_0 : STD_LOGIC;
  signal W_49_31_i_14_n_0 : STD_LOGIC;
  signal W_49_31_i_15_n_0 : STD_LOGIC;
  signal W_49_31_i_17_n_0 : STD_LOGIC;
  signal W_49_31_i_19_n_0 : STD_LOGIC;
  signal W_49_31_i_2_n_0 : STD_LOGIC;
  signal W_49_31_i_3_n_0 : STD_LOGIC;
  signal W_49_31_i_4_n_0 : STD_LOGIC;
  signal W_49_31_i_5_n_0 : STD_LOGIC;
  signal W_49_31_i_6_n_0 : STD_LOGIC;
  signal W_49_31_i_7_n_0 : STD_LOGIC;
  signal W_49_31_i_8_n_0 : STD_LOGIC;
  signal W_49_31_i_9_n_0 : STD_LOGIC;
  signal W_49_3_i_10_n_0 : STD_LOGIC;
  signal W_49_3_i_11_n_0 : STD_LOGIC;
  signal W_49_3_i_15_n_0 : STD_LOGIC;
  signal W_49_3_i_2_n_0 : STD_LOGIC;
  signal W_49_3_i_3_n_0 : STD_LOGIC;
  signal W_49_3_i_4_n_0 : STD_LOGIC;
  signal W_49_3_i_5_n_0 : STD_LOGIC;
  signal W_49_3_i_6_n_0 : STD_LOGIC;
  signal W_49_3_i_7_n_0 : STD_LOGIC;
  signal W_49_3_i_8_n_0 : STD_LOGIC;
  signal W_49_3_i_9_n_0 : STD_LOGIC;
  signal W_49_7_i_10_n_0 : STD_LOGIC;
  signal W_49_7_i_11_n_0 : STD_LOGIC;
  signal W_49_7_i_12_n_0 : STD_LOGIC;
  signal W_49_7_i_13_n_0 : STD_LOGIC;
  signal W_49_7_i_14_n_0 : STD_LOGIC;
  signal W_49_7_i_15_n_0 : STD_LOGIC;
  signal W_49_7_i_16_n_0 : STD_LOGIC;
  signal W_49_7_i_17_n_0 : STD_LOGIC;
  signal W_49_7_i_2_n_0 : STD_LOGIC;
  signal W_49_7_i_3_n_0 : STD_LOGIC;
  signal W_49_7_i_4_n_0 : STD_LOGIC;
  signal W_49_7_i_5_n_0 : STD_LOGIC;
  signal W_49_7_i_6_n_0 : STD_LOGIC;
  signal W_49_7_i_7_n_0 : STD_LOGIC;
  signal W_49_7_i_8_n_0 : STD_LOGIC;
  signal W_49_7_i_9_n_0 : STD_LOGIC;
  signal W_50_11_i_10_n_0 : STD_LOGIC;
  signal W_50_11_i_11_n_0 : STD_LOGIC;
  signal W_50_11_i_12_n_0 : STD_LOGIC;
  signal W_50_11_i_13_n_0 : STD_LOGIC;
  signal W_50_11_i_14_n_0 : STD_LOGIC;
  signal W_50_11_i_15_n_0 : STD_LOGIC;
  signal W_50_11_i_16_n_0 : STD_LOGIC;
  signal W_50_11_i_17_n_0 : STD_LOGIC;
  signal W_50_11_i_2_n_0 : STD_LOGIC;
  signal W_50_11_i_3_n_0 : STD_LOGIC;
  signal W_50_11_i_4_n_0 : STD_LOGIC;
  signal W_50_11_i_5_n_0 : STD_LOGIC;
  signal W_50_11_i_6_n_0 : STD_LOGIC;
  signal W_50_11_i_7_n_0 : STD_LOGIC;
  signal W_50_11_i_8_n_0 : STD_LOGIC;
  signal W_50_11_i_9_n_0 : STD_LOGIC;
  signal W_50_15_i_10_n_0 : STD_LOGIC;
  signal W_50_15_i_11_n_0 : STD_LOGIC;
  signal W_50_15_i_12_n_0 : STD_LOGIC;
  signal W_50_15_i_13_n_0 : STD_LOGIC;
  signal W_50_15_i_14_n_0 : STD_LOGIC;
  signal W_50_15_i_15_n_0 : STD_LOGIC;
  signal W_50_15_i_16_n_0 : STD_LOGIC;
  signal W_50_15_i_17_n_0 : STD_LOGIC;
  signal W_50_15_i_2_n_0 : STD_LOGIC;
  signal W_50_15_i_3_n_0 : STD_LOGIC;
  signal W_50_15_i_4_n_0 : STD_LOGIC;
  signal W_50_15_i_5_n_0 : STD_LOGIC;
  signal W_50_15_i_6_n_0 : STD_LOGIC;
  signal W_50_15_i_7_n_0 : STD_LOGIC;
  signal W_50_15_i_8_n_0 : STD_LOGIC;
  signal W_50_15_i_9_n_0 : STD_LOGIC;
  signal W_50_19_i_10_n_0 : STD_LOGIC;
  signal W_50_19_i_11_n_0 : STD_LOGIC;
  signal W_50_19_i_12_n_0 : STD_LOGIC;
  signal W_50_19_i_13_n_0 : STD_LOGIC;
  signal W_50_19_i_14_n_0 : STD_LOGIC;
  signal W_50_19_i_15_n_0 : STD_LOGIC;
  signal W_50_19_i_16_n_0 : STD_LOGIC;
  signal W_50_19_i_17_n_0 : STD_LOGIC;
  signal W_50_19_i_2_n_0 : STD_LOGIC;
  signal W_50_19_i_3_n_0 : STD_LOGIC;
  signal W_50_19_i_4_n_0 : STD_LOGIC;
  signal W_50_19_i_5_n_0 : STD_LOGIC;
  signal W_50_19_i_6_n_0 : STD_LOGIC;
  signal W_50_19_i_7_n_0 : STD_LOGIC;
  signal W_50_19_i_8_n_0 : STD_LOGIC;
  signal W_50_19_i_9_n_0 : STD_LOGIC;
  signal W_50_23_i_10_n_0 : STD_LOGIC;
  signal W_50_23_i_11_n_0 : STD_LOGIC;
  signal W_50_23_i_12_n_0 : STD_LOGIC;
  signal W_50_23_i_13_n_0 : STD_LOGIC;
  signal W_50_23_i_14_n_0 : STD_LOGIC;
  signal W_50_23_i_15_n_0 : STD_LOGIC;
  signal W_50_23_i_16_n_0 : STD_LOGIC;
  signal W_50_23_i_17_n_0 : STD_LOGIC;
  signal W_50_23_i_2_n_0 : STD_LOGIC;
  signal W_50_23_i_3_n_0 : STD_LOGIC;
  signal W_50_23_i_4_n_0 : STD_LOGIC;
  signal W_50_23_i_5_n_0 : STD_LOGIC;
  signal W_50_23_i_6_n_0 : STD_LOGIC;
  signal W_50_23_i_7_n_0 : STD_LOGIC;
  signal W_50_23_i_8_n_0 : STD_LOGIC;
  signal W_50_23_i_9_n_0 : STD_LOGIC;
  signal W_50_27_i_10_n_0 : STD_LOGIC;
  signal W_50_27_i_11_n_0 : STD_LOGIC;
  signal W_50_27_i_12_n_0 : STD_LOGIC;
  signal W_50_27_i_13_n_0 : STD_LOGIC;
  signal W_50_27_i_14_n_0 : STD_LOGIC;
  signal W_50_27_i_15_n_0 : STD_LOGIC;
  signal W_50_27_i_16_n_0 : STD_LOGIC;
  signal W_50_27_i_17_n_0 : STD_LOGIC;
  signal W_50_27_i_2_n_0 : STD_LOGIC;
  signal W_50_27_i_3_n_0 : STD_LOGIC;
  signal W_50_27_i_4_n_0 : STD_LOGIC;
  signal W_50_27_i_5_n_0 : STD_LOGIC;
  signal W_50_27_i_6_n_0 : STD_LOGIC;
  signal W_50_27_i_7_n_0 : STD_LOGIC;
  signal W_50_27_i_8_n_0 : STD_LOGIC;
  signal W_50_27_i_9_n_0 : STD_LOGIC;
  signal W_50_31_i_10_n_0 : STD_LOGIC;
  signal W_50_31_i_11_n_0 : STD_LOGIC;
  signal W_50_31_i_12_n_0 : STD_LOGIC;
  signal W_50_31_i_13_n_0 : STD_LOGIC;
  signal W_50_31_i_14_n_0 : STD_LOGIC;
  signal W_50_31_i_15_n_0 : STD_LOGIC;
  signal W_50_31_i_17_n_0 : STD_LOGIC;
  signal W_50_31_i_19_n_0 : STD_LOGIC;
  signal W_50_31_i_2_n_0 : STD_LOGIC;
  signal W_50_31_i_3_n_0 : STD_LOGIC;
  signal W_50_31_i_4_n_0 : STD_LOGIC;
  signal W_50_31_i_5_n_0 : STD_LOGIC;
  signal W_50_31_i_6_n_0 : STD_LOGIC;
  signal W_50_31_i_7_n_0 : STD_LOGIC;
  signal W_50_31_i_8_n_0 : STD_LOGIC;
  signal W_50_31_i_9_n_0 : STD_LOGIC;
  signal W_50_3_i_10_n_0 : STD_LOGIC;
  signal W_50_3_i_11_n_0 : STD_LOGIC;
  signal W_50_3_i_15_n_0 : STD_LOGIC;
  signal W_50_3_i_2_n_0 : STD_LOGIC;
  signal W_50_3_i_3_n_0 : STD_LOGIC;
  signal W_50_3_i_4_n_0 : STD_LOGIC;
  signal W_50_3_i_5_n_0 : STD_LOGIC;
  signal W_50_3_i_6_n_0 : STD_LOGIC;
  signal W_50_3_i_7_n_0 : STD_LOGIC;
  signal W_50_3_i_8_n_0 : STD_LOGIC;
  signal W_50_3_i_9_n_0 : STD_LOGIC;
  signal W_50_7_i_10_n_0 : STD_LOGIC;
  signal W_50_7_i_11_n_0 : STD_LOGIC;
  signal W_50_7_i_12_n_0 : STD_LOGIC;
  signal W_50_7_i_13_n_0 : STD_LOGIC;
  signal W_50_7_i_14_n_0 : STD_LOGIC;
  signal W_50_7_i_15_n_0 : STD_LOGIC;
  signal W_50_7_i_16_n_0 : STD_LOGIC;
  signal W_50_7_i_17_n_0 : STD_LOGIC;
  signal W_50_7_i_2_n_0 : STD_LOGIC;
  signal W_50_7_i_3_n_0 : STD_LOGIC;
  signal W_50_7_i_4_n_0 : STD_LOGIC;
  signal W_50_7_i_5_n_0 : STD_LOGIC;
  signal W_50_7_i_6_n_0 : STD_LOGIC;
  signal W_50_7_i_7_n_0 : STD_LOGIC;
  signal W_50_7_i_8_n_0 : STD_LOGIC;
  signal W_50_7_i_9_n_0 : STD_LOGIC;
  signal W_51_11_i_10_n_0 : STD_LOGIC;
  signal W_51_11_i_11_n_0 : STD_LOGIC;
  signal W_51_11_i_12_n_0 : STD_LOGIC;
  signal W_51_11_i_13_n_0 : STD_LOGIC;
  signal W_51_11_i_14_n_0 : STD_LOGIC;
  signal W_51_11_i_15_n_0 : STD_LOGIC;
  signal W_51_11_i_16_n_0 : STD_LOGIC;
  signal W_51_11_i_17_n_0 : STD_LOGIC;
  signal W_51_11_i_2_n_0 : STD_LOGIC;
  signal W_51_11_i_3_n_0 : STD_LOGIC;
  signal W_51_11_i_4_n_0 : STD_LOGIC;
  signal W_51_11_i_5_n_0 : STD_LOGIC;
  signal W_51_11_i_6_n_0 : STD_LOGIC;
  signal W_51_11_i_7_n_0 : STD_LOGIC;
  signal W_51_11_i_8_n_0 : STD_LOGIC;
  signal W_51_11_i_9_n_0 : STD_LOGIC;
  signal W_51_15_i_10_n_0 : STD_LOGIC;
  signal W_51_15_i_11_n_0 : STD_LOGIC;
  signal W_51_15_i_12_n_0 : STD_LOGIC;
  signal W_51_15_i_13_n_0 : STD_LOGIC;
  signal W_51_15_i_14_n_0 : STD_LOGIC;
  signal W_51_15_i_15_n_0 : STD_LOGIC;
  signal W_51_15_i_16_n_0 : STD_LOGIC;
  signal W_51_15_i_17_n_0 : STD_LOGIC;
  signal W_51_15_i_2_n_0 : STD_LOGIC;
  signal W_51_15_i_3_n_0 : STD_LOGIC;
  signal W_51_15_i_4_n_0 : STD_LOGIC;
  signal W_51_15_i_5_n_0 : STD_LOGIC;
  signal W_51_15_i_6_n_0 : STD_LOGIC;
  signal W_51_15_i_7_n_0 : STD_LOGIC;
  signal W_51_15_i_8_n_0 : STD_LOGIC;
  signal W_51_15_i_9_n_0 : STD_LOGIC;
  signal W_51_19_i_10_n_0 : STD_LOGIC;
  signal W_51_19_i_11_n_0 : STD_LOGIC;
  signal W_51_19_i_12_n_0 : STD_LOGIC;
  signal W_51_19_i_13_n_0 : STD_LOGIC;
  signal W_51_19_i_14_n_0 : STD_LOGIC;
  signal W_51_19_i_15_n_0 : STD_LOGIC;
  signal W_51_19_i_16_n_0 : STD_LOGIC;
  signal W_51_19_i_17_n_0 : STD_LOGIC;
  signal W_51_19_i_2_n_0 : STD_LOGIC;
  signal W_51_19_i_3_n_0 : STD_LOGIC;
  signal W_51_19_i_4_n_0 : STD_LOGIC;
  signal W_51_19_i_5_n_0 : STD_LOGIC;
  signal W_51_19_i_6_n_0 : STD_LOGIC;
  signal W_51_19_i_7_n_0 : STD_LOGIC;
  signal W_51_19_i_8_n_0 : STD_LOGIC;
  signal W_51_19_i_9_n_0 : STD_LOGIC;
  signal W_51_23_i_10_n_0 : STD_LOGIC;
  signal W_51_23_i_11_n_0 : STD_LOGIC;
  signal W_51_23_i_12_n_0 : STD_LOGIC;
  signal W_51_23_i_13_n_0 : STD_LOGIC;
  signal W_51_23_i_14_n_0 : STD_LOGIC;
  signal W_51_23_i_15_n_0 : STD_LOGIC;
  signal W_51_23_i_16_n_0 : STD_LOGIC;
  signal W_51_23_i_17_n_0 : STD_LOGIC;
  signal W_51_23_i_2_n_0 : STD_LOGIC;
  signal W_51_23_i_3_n_0 : STD_LOGIC;
  signal W_51_23_i_4_n_0 : STD_LOGIC;
  signal W_51_23_i_5_n_0 : STD_LOGIC;
  signal W_51_23_i_6_n_0 : STD_LOGIC;
  signal W_51_23_i_7_n_0 : STD_LOGIC;
  signal W_51_23_i_8_n_0 : STD_LOGIC;
  signal W_51_23_i_9_n_0 : STD_LOGIC;
  signal W_51_27_i_10_n_0 : STD_LOGIC;
  signal W_51_27_i_11_n_0 : STD_LOGIC;
  signal W_51_27_i_12_n_0 : STD_LOGIC;
  signal W_51_27_i_13_n_0 : STD_LOGIC;
  signal W_51_27_i_14_n_0 : STD_LOGIC;
  signal W_51_27_i_15_n_0 : STD_LOGIC;
  signal W_51_27_i_16_n_0 : STD_LOGIC;
  signal W_51_27_i_17_n_0 : STD_LOGIC;
  signal W_51_27_i_2_n_0 : STD_LOGIC;
  signal W_51_27_i_3_n_0 : STD_LOGIC;
  signal W_51_27_i_4_n_0 : STD_LOGIC;
  signal W_51_27_i_5_n_0 : STD_LOGIC;
  signal W_51_27_i_6_n_0 : STD_LOGIC;
  signal W_51_27_i_7_n_0 : STD_LOGIC;
  signal W_51_27_i_8_n_0 : STD_LOGIC;
  signal W_51_27_i_9_n_0 : STD_LOGIC;
  signal W_51_31_i_10_n_0 : STD_LOGIC;
  signal W_51_31_i_11_n_0 : STD_LOGIC;
  signal W_51_31_i_12_n_0 : STD_LOGIC;
  signal W_51_31_i_13_n_0 : STD_LOGIC;
  signal W_51_31_i_14_n_0 : STD_LOGIC;
  signal W_51_31_i_15_n_0 : STD_LOGIC;
  signal W_51_31_i_17_n_0 : STD_LOGIC;
  signal W_51_31_i_19_n_0 : STD_LOGIC;
  signal W_51_31_i_2_n_0 : STD_LOGIC;
  signal W_51_31_i_3_n_0 : STD_LOGIC;
  signal W_51_31_i_4_n_0 : STD_LOGIC;
  signal W_51_31_i_5_n_0 : STD_LOGIC;
  signal W_51_31_i_6_n_0 : STD_LOGIC;
  signal W_51_31_i_7_n_0 : STD_LOGIC;
  signal W_51_31_i_8_n_0 : STD_LOGIC;
  signal W_51_31_i_9_n_0 : STD_LOGIC;
  signal W_51_3_i_10_n_0 : STD_LOGIC;
  signal W_51_3_i_11_n_0 : STD_LOGIC;
  signal W_51_3_i_15_n_0 : STD_LOGIC;
  signal W_51_3_i_2_n_0 : STD_LOGIC;
  signal W_51_3_i_3_n_0 : STD_LOGIC;
  signal W_51_3_i_4_n_0 : STD_LOGIC;
  signal W_51_3_i_5_n_0 : STD_LOGIC;
  signal W_51_3_i_6_n_0 : STD_LOGIC;
  signal W_51_3_i_7_n_0 : STD_LOGIC;
  signal W_51_3_i_8_n_0 : STD_LOGIC;
  signal W_51_3_i_9_n_0 : STD_LOGIC;
  signal W_51_7_i_10_n_0 : STD_LOGIC;
  signal W_51_7_i_11_n_0 : STD_LOGIC;
  signal W_51_7_i_12_n_0 : STD_LOGIC;
  signal W_51_7_i_13_n_0 : STD_LOGIC;
  signal W_51_7_i_14_n_0 : STD_LOGIC;
  signal W_51_7_i_15_n_0 : STD_LOGIC;
  signal W_51_7_i_16_n_0 : STD_LOGIC;
  signal W_51_7_i_17_n_0 : STD_LOGIC;
  signal W_51_7_i_2_n_0 : STD_LOGIC;
  signal W_51_7_i_3_n_0 : STD_LOGIC;
  signal W_51_7_i_4_n_0 : STD_LOGIC;
  signal W_51_7_i_5_n_0 : STD_LOGIC;
  signal W_51_7_i_6_n_0 : STD_LOGIC;
  signal W_51_7_i_7_n_0 : STD_LOGIC;
  signal W_51_7_i_8_n_0 : STD_LOGIC;
  signal W_51_7_i_9_n_0 : STD_LOGIC;
  signal W_52_11_i_10_n_0 : STD_LOGIC;
  signal W_52_11_i_11_n_0 : STD_LOGIC;
  signal W_52_11_i_12_n_0 : STD_LOGIC;
  signal W_52_11_i_13_n_0 : STD_LOGIC;
  signal W_52_11_i_14_n_0 : STD_LOGIC;
  signal W_52_11_i_15_n_0 : STD_LOGIC;
  signal W_52_11_i_16_n_0 : STD_LOGIC;
  signal W_52_11_i_17_n_0 : STD_LOGIC;
  signal W_52_11_i_2_n_0 : STD_LOGIC;
  signal W_52_11_i_3_n_0 : STD_LOGIC;
  signal W_52_11_i_4_n_0 : STD_LOGIC;
  signal W_52_11_i_5_n_0 : STD_LOGIC;
  signal W_52_11_i_6_n_0 : STD_LOGIC;
  signal W_52_11_i_7_n_0 : STD_LOGIC;
  signal W_52_11_i_8_n_0 : STD_LOGIC;
  signal W_52_11_i_9_n_0 : STD_LOGIC;
  signal W_52_15_i_10_n_0 : STD_LOGIC;
  signal W_52_15_i_11_n_0 : STD_LOGIC;
  signal W_52_15_i_12_n_0 : STD_LOGIC;
  signal W_52_15_i_13_n_0 : STD_LOGIC;
  signal W_52_15_i_14_n_0 : STD_LOGIC;
  signal W_52_15_i_15_n_0 : STD_LOGIC;
  signal W_52_15_i_16_n_0 : STD_LOGIC;
  signal W_52_15_i_17_n_0 : STD_LOGIC;
  signal W_52_15_i_2_n_0 : STD_LOGIC;
  signal W_52_15_i_3_n_0 : STD_LOGIC;
  signal W_52_15_i_4_n_0 : STD_LOGIC;
  signal W_52_15_i_5_n_0 : STD_LOGIC;
  signal W_52_15_i_6_n_0 : STD_LOGIC;
  signal W_52_15_i_7_n_0 : STD_LOGIC;
  signal W_52_15_i_8_n_0 : STD_LOGIC;
  signal W_52_15_i_9_n_0 : STD_LOGIC;
  signal W_52_19_i_10_n_0 : STD_LOGIC;
  signal W_52_19_i_11_n_0 : STD_LOGIC;
  signal W_52_19_i_12_n_0 : STD_LOGIC;
  signal W_52_19_i_13_n_0 : STD_LOGIC;
  signal W_52_19_i_14_n_0 : STD_LOGIC;
  signal W_52_19_i_15_n_0 : STD_LOGIC;
  signal W_52_19_i_16_n_0 : STD_LOGIC;
  signal W_52_19_i_17_n_0 : STD_LOGIC;
  signal W_52_19_i_2_n_0 : STD_LOGIC;
  signal W_52_19_i_3_n_0 : STD_LOGIC;
  signal W_52_19_i_4_n_0 : STD_LOGIC;
  signal W_52_19_i_5_n_0 : STD_LOGIC;
  signal W_52_19_i_6_n_0 : STD_LOGIC;
  signal W_52_19_i_7_n_0 : STD_LOGIC;
  signal W_52_19_i_8_n_0 : STD_LOGIC;
  signal W_52_19_i_9_n_0 : STD_LOGIC;
  signal W_52_23_i_10_n_0 : STD_LOGIC;
  signal W_52_23_i_11_n_0 : STD_LOGIC;
  signal W_52_23_i_12_n_0 : STD_LOGIC;
  signal W_52_23_i_13_n_0 : STD_LOGIC;
  signal W_52_23_i_14_n_0 : STD_LOGIC;
  signal W_52_23_i_15_n_0 : STD_LOGIC;
  signal W_52_23_i_16_n_0 : STD_LOGIC;
  signal W_52_23_i_17_n_0 : STD_LOGIC;
  signal W_52_23_i_2_n_0 : STD_LOGIC;
  signal W_52_23_i_3_n_0 : STD_LOGIC;
  signal W_52_23_i_4_n_0 : STD_LOGIC;
  signal W_52_23_i_5_n_0 : STD_LOGIC;
  signal W_52_23_i_6_n_0 : STD_LOGIC;
  signal W_52_23_i_7_n_0 : STD_LOGIC;
  signal W_52_23_i_8_n_0 : STD_LOGIC;
  signal W_52_23_i_9_n_0 : STD_LOGIC;
  signal W_52_27_i_10_n_0 : STD_LOGIC;
  signal W_52_27_i_11_n_0 : STD_LOGIC;
  signal W_52_27_i_12_n_0 : STD_LOGIC;
  signal W_52_27_i_13_n_0 : STD_LOGIC;
  signal W_52_27_i_14_n_0 : STD_LOGIC;
  signal W_52_27_i_15_n_0 : STD_LOGIC;
  signal W_52_27_i_16_n_0 : STD_LOGIC;
  signal W_52_27_i_17_n_0 : STD_LOGIC;
  signal W_52_27_i_2_n_0 : STD_LOGIC;
  signal W_52_27_i_3_n_0 : STD_LOGIC;
  signal W_52_27_i_4_n_0 : STD_LOGIC;
  signal W_52_27_i_5_n_0 : STD_LOGIC;
  signal W_52_27_i_6_n_0 : STD_LOGIC;
  signal W_52_27_i_7_n_0 : STD_LOGIC;
  signal W_52_27_i_8_n_0 : STD_LOGIC;
  signal W_52_27_i_9_n_0 : STD_LOGIC;
  signal W_52_31_i_10_n_0 : STD_LOGIC;
  signal W_52_31_i_11_n_0 : STD_LOGIC;
  signal W_52_31_i_12_n_0 : STD_LOGIC;
  signal W_52_31_i_13_n_0 : STD_LOGIC;
  signal W_52_31_i_14_n_0 : STD_LOGIC;
  signal W_52_31_i_15_n_0 : STD_LOGIC;
  signal W_52_31_i_17_n_0 : STD_LOGIC;
  signal W_52_31_i_19_n_0 : STD_LOGIC;
  signal W_52_31_i_2_n_0 : STD_LOGIC;
  signal W_52_31_i_3_n_0 : STD_LOGIC;
  signal W_52_31_i_4_n_0 : STD_LOGIC;
  signal W_52_31_i_5_n_0 : STD_LOGIC;
  signal W_52_31_i_6_n_0 : STD_LOGIC;
  signal W_52_31_i_7_n_0 : STD_LOGIC;
  signal W_52_31_i_8_n_0 : STD_LOGIC;
  signal W_52_31_i_9_n_0 : STD_LOGIC;
  signal W_52_3_i_10_n_0 : STD_LOGIC;
  signal W_52_3_i_11_n_0 : STD_LOGIC;
  signal W_52_3_i_15_n_0 : STD_LOGIC;
  signal W_52_3_i_2_n_0 : STD_LOGIC;
  signal W_52_3_i_3_n_0 : STD_LOGIC;
  signal W_52_3_i_4_n_0 : STD_LOGIC;
  signal W_52_3_i_5_n_0 : STD_LOGIC;
  signal W_52_3_i_6_n_0 : STD_LOGIC;
  signal W_52_3_i_7_n_0 : STD_LOGIC;
  signal W_52_3_i_8_n_0 : STD_LOGIC;
  signal W_52_3_i_9_n_0 : STD_LOGIC;
  signal W_52_7_i_10_n_0 : STD_LOGIC;
  signal W_52_7_i_11_n_0 : STD_LOGIC;
  signal W_52_7_i_12_n_0 : STD_LOGIC;
  signal W_52_7_i_13_n_0 : STD_LOGIC;
  signal W_52_7_i_14_n_0 : STD_LOGIC;
  signal W_52_7_i_15_n_0 : STD_LOGIC;
  signal W_52_7_i_16_n_0 : STD_LOGIC;
  signal W_52_7_i_17_n_0 : STD_LOGIC;
  signal W_52_7_i_2_n_0 : STD_LOGIC;
  signal W_52_7_i_3_n_0 : STD_LOGIC;
  signal W_52_7_i_4_n_0 : STD_LOGIC;
  signal W_52_7_i_5_n_0 : STD_LOGIC;
  signal W_52_7_i_6_n_0 : STD_LOGIC;
  signal W_52_7_i_7_n_0 : STD_LOGIC;
  signal W_52_7_i_8_n_0 : STD_LOGIC;
  signal W_52_7_i_9_n_0 : STD_LOGIC;
  signal W_53_11_i_10_n_0 : STD_LOGIC;
  signal W_53_11_i_11_n_0 : STD_LOGIC;
  signal W_53_11_i_12_n_0 : STD_LOGIC;
  signal W_53_11_i_13_n_0 : STD_LOGIC;
  signal W_53_11_i_14_n_0 : STD_LOGIC;
  signal W_53_11_i_15_n_0 : STD_LOGIC;
  signal W_53_11_i_16_n_0 : STD_LOGIC;
  signal W_53_11_i_17_n_0 : STD_LOGIC;
  signal W_53_11_i_2_n_0 : STD_LOGIC;
  signal W_53_11_i_3_n_0 : STD_LOGIC;
  signal W_53_11_i_4_n_0 : STD_LOGIC;
  signal W_53_11_i_5_n_0 : STD_LOGIC;
  signal W_53_11_i_6_n_0 : STD_LOGIC;
  signal W_53_11_i_7_n_0 : STD_LOGIC;
  signal W_53_11_i_8_n_0 : STD_LOGIC;
  signal W_53_11_i_9_n_0 : STD_LOGIC;
  signal W_53_15_i_10_n_0 : STD_LOGIC;
  signal W_53_15_i_11_n_0 : STD_LOGIC;
  signal W_53_15_i_12_n_0 : STD_LOGIC;
  signal W_53_15_i_13_n_0 : STD_LOGIC;
  signal W_53_15_i_14_n_0 : STD_LOGIC;
  signal W_53_15_i_15_n_0 : STD_LOGIC;
  signal W_53_15_i_16_n_0 : STD_LOGIC;
  signal W_53_15_i_17_n_0 : STD_LOGIC;
  signal W_53_15_i_2_n_0 : STD_LOGIC;
  signal W_53_15_i_3_n_0 : STD_LOGIC;
  signal W_53_15_i_4_n_0 : STD_LOGIC;
  signal W_53_15_i_5_n_0 : STD_LOGIC;
  signal W_53_15_i_6_n_0 : STD_LOGIC;
  signal W_53_15_i_7_n_0 : STD_LOGIC;
  signal W_53_15_i_8_n_0 : STD_LOGIC;
  signal W_53_15_i_9_n_0 : STD_LOGIC;
  signal W_53_19_i_10_n_0 : STD_LOGIC;
  signal W_53_19_i_11_n_0 : STD_LOGIC;
  signal W_53_19_i_12_n_0 : STD_LOGIC;
  signal W_53_19_i_13_n_0 : STD_LOGIC;
  signal W_53_19_i_14_n_0 : STD_LOGIC;
  signal W_53_19_i_15_n_0 : STD_LOGIC;
  signal W_53_19_i_16_n_0 : STD_LOGIC;
  signal W_53_19_i_17_n_0 : STD_LOGIC;
  signal W_53_19_i_2_n_0 : STD_LOGIC;
  signal W_53_19_i_3_n_0 : STD_LOGIC;
  signal W_53_19_i_4_n_0 : STD_LOGIC;
  signal W_53_19_i_5_n_0 : STD_LOGIC;
  signal W_53_19_i_6_n_0 : STD_LOGIC;
  signal W_53_19_i_7_n_0 : STD_LOGIC;
  signal W_53_19_i_8_n_0 : STD_LOGIC;
  signal W_53_19_i_9_n_0 : STD_LOGIC;
  signal W_53_23_i_10_n_0 : STD_LOGIC;
  signal W_53_23_i_11_n_0 : STD_LOGIC;
  signal W_53_23_i_12_n_0 : STD_LOGIC;
  signal W_53_23_i_13_n_0 : STD_LOGIC;
  signal W_53_23_i_14_n_0 : STD_LOGIC;
  signal W_53_23_i_15_n_0 : STD_LOGIC;
  signal W_53_23_i_16_n_0 : STD_LOGIC;
  signal W_53_23_i_17_n_0 : STD_LOGIC;
  signal W_53_23_i_2_n_0 : STD_LOGIC;
  signal W_53_23_i_3_n_0 : STD_LOGIC;
  signal W_53_23_i_4_n_0 : STD_LOGIC;
  signal W_53_23_i_5_n_0 : STD_LOGIC;
  signal W_53_23_i_6_n_0 : STD_LOGIC;
  signal W_53_23_i_7_n_0 : STD_LOGIC;
  signal W_53_23_i_8_n_0 : STD_LOGIC;
  signal W_53_23_i_9_n_0 : STD_LOGIC;
  signal W_53_27_i_10_n_0 : STD_LOGIC;
  signal W_53_27_i_11_n_0 : STD_LOGIC;
  signal W_53_27_i_12_n_0 : STD_LOGIC;
  signal W_53_27_i_13_n_0 : STD_LOGIC;
  signal W_53_27_i_14_n_0 : STD_LOGIC;
  signal W_53_27_i_15_n_0 : STD_LOGIC;
  signal W_53_27_i_16_n_0 : STD_LOGIC;
  signal W_53_27_i_17_n_0 : STD_LOGIC;
  signal W_53_27_i_2_n_0 : STD_LOGIC;
  signal W_53_27_i_3_n_0 : STD_LOGIC;
  signal W_53_27_i_4_n_0 : STD_LOGIC;
  signal W_53_27_i_5_n_0 : STD_LOGIC;
  signal W_53_27_i_6_n_0 : STD_LOGIC;
  signal W_53_27_i_7_n_0 : STD_LOGIC;
  signal W_53_27_i_8_n_0 : STD_LOGIC;
  signal W_53_27_i_9_n_0 : STD_LOGIC;
  signal W_53_31_i_10_n_0 : STD_LOGIC;
  signal W_53_31_i_11_n_0 : STD_LOGIC;
  signal W_53_31_i_12_n_0 : STD_LOGIC;
  signal W_53_31_i_13_n_0 : STD_LOGIC;
  signal W_53_31_i_14_n_0 : STD_LOGIC;
  signal W_53_31_i_15_n_0 : STD_LOGIC;
  signal W_53_31_i_17_n_0 : STD_LOGIC;
  signal W_53_31_i_19_n_0 : STD_LOGIC;
  signal W_53_31_i_2_n_0 : STD_LOGIC;
  signal W_53_31_i_3_n_0 : STD_LOGIC;
  signal W_53_31_i_4_n_0 : STD_LOGIC;
  signal W_53_31_i_5_n_0 : STD_LOGIC;
  signal W_53_31_i_6_n_0 : STD_LOGIC;
  signal W_53_31_i_7_n_0 : STD_LOGIC;
  signal W_53_31_i_8_n_0 : STD_LOGIC;
  signal W_53_31_i_9_n_0 : STD_LOGIC;
  signal W_53_3_i_10_n_0 : STD_LOGIC;
  signal W_53_3_i_11_n_0 : STD_LOGIC;
  signal W_53_3_i_15_n_0 : STD_LOGIC;
  signal W_53_3_i_2_n_0 : STD_LOGIC;
  signal W_53_3_i_3_n_0 : STD_LOGIC;
  signal W_53_3_i_4_n_0 : STD_LOGIC;
  signal W_53_3_i_5_n_0 : STD_LOGIC;
  signal W_53_3_i_6_n_0 : STD_LOGIC;
  signal W_53_3_i_7_n_0 : STD_LOGIC;
  signal W_53_3_i_8_n_0 : STD_LOGIC;
  signal W_53_3_i_9_n_0 : STD_LOGIC;
  signal W_53_7_i_10_n_0 : STD_LOGIC;
  signal W_53_7_i_11_n_0 : STD_LOGIC;
  signal W_53_7_i_12_n_0 : STD_LOGIC;
  signal W_53_7_i_13_n_0 : STD_LOGIC;
  signal W_53_7_i_14_n_0 : STD_LOGIC;
  signal W_53_7_i_15_n_0 : STD_LOGIC;
  signal W_53_7_i_16_n_0 : STD_LOGIC;
  signal W_53_7_i_17_n_0 : STD_LOGIC;
  signal W_53_7_i_2_n_0 : STD_LOGIC;
  signal W_53_7_i_3_n_0 : STD_LOGIC;
  signal W_53_7_i_4_n_0 : STD_LOGIC;
  signal W_53_7_i_5_n_0 : STD_LOGIC;
  signal W_53_7_i_6_n_0 : STD_LOGIC;
  signal W_53_7_i_7_n_0 : STD_LOGIC;
  signal W_53_7_i_8_n_0 : STD_LOGIC;
  signal W_53_7_i_9_n_0 : STD_LOGIC;
  signal W_54_11_i_10_n_0 : STD_LOGIC;
  signal W_54_11_i_11_n_0 : STD_LOGIC;
  signal W_54_11_i_12_n_0 : STD_LOGIC;
  signal W_54_11_i_13_n_0 : STD_LOGIC;
  signal W_54_11_i_14_n_0 : STD_LOGIC;
  signal W_54_11_i_15_n_0 : STD_LOGIC;
  signal W_54_11_i_16_n_0 : STD_LOGIC;
  signal W_54_11_i_17_n_0 : STD_LOGIC;
  signal W_54_11_i_2_n_0 : STD_LOGIC;
  signal W_54_11_i_3_n_0 : STD_LOGIC;
  signal W_54_11_i_4_n_0 : STD_LOGIC;
  signal W_54_11_i_5_n_0 : STD_LOGIC;
  signal W_54_11_i_6_n_0 : STD_LOGIC;
  signal W_54_11_i_7_n_0 : STD_LOGIC;
  signal W_54_11_i_8_n_0 : STD_LOGIC;
  signal W_54_11_i_9_n_0 : STD_LOGIC;
  signal W_54_15_i_10_n_0 : STD_LOGIC;
  signal W_54_15_i_11_n_0 : STD_LOGIC;
  signal W_54_15_i_12_n_0 : STD_LOGIC;
  signal W_54_15_i_13_n_0 : STD_LOGIC;
  signal W_54_15_i_14_n_0 : STD_LOGIC;
  signal W_54_15_i_15_n_0 : STD_LOGIC;
  signal W_54_15_i_16_n_0 : STD_LOGIC;
  signal W_54_15_i_17_n_0 : STD_LOGIC;
  signal W_54_15_i_2_n_0 : STD_LOGIC;
  signal W_54_15_i_3_n_0 : STD_LOGIC;
  signal W_54_15_i_4_n_0 : STD_LOGIC;
  signal W_54_15_i_5_n_0 : STD_LOGIC;
  signal W_54_15_i_6_n_0 : STD_LOGIC;
  signal W_54_15_i_7_n_0 : STD_LOGIC;
  signal W_54_15_i_8_n_0 : STD_LOGIC;
  signal W_54_15_i_9_n_0 : STD_LOGIC;
  signal W_54_19_i_10_n_0 : STD_LOGIC;
  signal W_54_19_i_11_n_0 : STD_LOGIC;
  signal W_54_19_i_12_n_0 : STD_LOGIC;
  signal W_54_19_i_13_n_0 : STD_LOGIC;
  signal W_54_19_i_14_n_0 : STD_LOGIC;
  signal W_54_19_i_15_n_0 : STD_LOGIC;
  signal W_54_19_i_16_n_0 : STD_LOGIC;
  signal W_54_19_i_17_n_0 : STD_LOGIC;
  signal W_54_19_i_2_n_0 : STD_LOGIC;
  signal W_54_19_i_3_n_0 : STD_LOGIC;
  signal W_54_19_i_4_n_0 : STD_LOGIC;
  signal W_54_19_i_5_n_0 : STD_LOGIC;
  signal W_54_19_i_6_n_0 : STD_LOGIC;
  signal W_54_19_i_7_n_0 : STD_LOGIC;
  signal W_54_19_i_8_n_0 : STD_LOGIC;
  signal W_54_19_i_9_n_0 : STD_LOGIC;
  signal W_54_23_i_10_n_0 : STD_LOGIC;
  signal W_54_23_i_11_n_0 : STD_LOGIC;
  signal W_54_23_i_12_n_0 : STD_LOGIC;
  signal W_54_23_i_13_n_0 : STD_LOGIC;
  signal W_54_23_i_14_n_0 : STD_LOGIC;
  signal W_54_23_i_15_n_0 : STD_LOGIC;
  signal W_54_23_i_16_n_0 : STD_LOGIC;
  signal W_54_23_i_17_n_0 : STD_LOGIC;
  signal W_54_23_i_2_n_0 : STD_LOGIC;
  signal W_54_23_i_3_n_0 : STD_LOGIC;
  signal W_54_23_i_4_n_0 : STD_LOGIC;
  signal W_54_23_i_5_n_0 : STD_LOGIC;
  signal W_54_23_i_6_n_0 : STD_LOGIC;
  signal W_54_23_i_7_n_0 : STD_LOGIC;
  signal W_54_23_i_8_n_0 : STD_LOGIC;
  signal W_54_23_i_9_n_0 : STD_LOGIC;
  signal W_54_27_i_10_n_0 : STD_LOGIC;
  signal W_54_27_i_11_n_0 : STD_LOGIC;
  signal W_54_27_i_12_n_0 : STD_LOGIC;
  signal W_54_27_i_13_n_0 : STD_LOGIC;
  signal W_54_27_i_14_n_0 : STD_LOGIC;
  signal W_54_27_i_15_n_0 : STD_LOGIC;
  signal W_54_27_i_16_n_0 : STD_LOGIC;
  signal W_54_27_i_17_n_0 : STD_LOGIC;
  signal W_54_27_i_2_n_0 : STD_LOGIC;
  signal W_54_27_i_3_n_0 : STD_LOGIC;
  signal W_54_27_i_4_n_0 : STD_LOGIC;
  signal W_54_27_i_5_n_0 : STD_LOGIC;
  signal W_54_27_i_6_n_0 : STD_LOGIC;
  signal W_54_27_i_7_n_0 : STD_LOGIC;
  signal W_54_27_i_8_n_0 : STD_LOGIC;
  signal W_54_27_i_9_n_0 : STD_LOGIC;
  signal W_54_31_i_10_n_0 : STD_LOGIC;
  signal W_54_31_i_11_n_0 : STD_LOGIC;
  signal W_54_31_i_12_n_0 : STD_LOGIC;
  signal W_54_31_i_13_n_0 : STD_LOGIC;
  signal W_54_31_i_14_n_0 : STD_LOGIC;
  signal W_54_31_i_15_n_0 : STD_LOGIC;
  signal W_54_31_i_17_n_0 : STD_LOGIC;
  signal W_54_31_i_19_n_0 : STD_LOGIC;
  signal W_54_31_i_2_n_0 : STD_LOGIC;
  signal W_54_31_i_3_n_0 : STD_LOGIC;
  signal W_54_31_i_4_n_0 : STD_LOGIC;
  signal W_54_31_i_5_n_0 : STD_LOGIC;
  signal W_54_31_i_6_n_0 : STD_LOGIC;
  signal W_54_31_i_7_n_0 : STD_LOGIC;
  signal W_54_31_i_8_n_0 : STD_LOGIC;
  signal W_54_31_i_9_n_0 : STD_LOGIC;
  signal W_54_3_i_10_n_0 : STD_LOGIC;
  signal W_54_3_i_11_n_0 : STD_LOGIC;
  signal W_54_3_i_15_n_0 : STD_LOGIC;
  signal W_54_3_i_2_n_0 : STD_LOGIC;
  signal W_54_3_i_3_n_0 : STD_LOGIC;
  signal W_54_3_i_4_n_0 : STD_LOGIC;
  signal W_54_3_i_5_n_0 : STD_LOGIC;
  signal W_54_3_i_6_n_0 : STD_LOGIC;
  signal W_54_3_i_7_n_0 : STD_LOGIC;
  signal W_54_3_i_8_n_0 : STD_LOGIC;
  signal W_54_3_i_9_n_0 : STD_LOGIC;
  signal W_54_7_i_10_n_0 : STD_LOGIC;
  signal W_54_7_i_11_n_0 : STD_LOGIC;
  signal W_54_7_i_12_n_0 : STD_LOGIC;
  signal W_54_7_i_13_n_0 : STD_LOGIC;
  signal W_54_7_i_14_n_0 : STD_LOGIC;
  signal W_54_7_i_15_n_0 : STD_LOGIC;
  signal W_54_7_i_16_n_0 : STD_LOGIC;
  signal W_54_7_i_17_n_0 : STD_LOGIC;
  signal W_54_7_i_2_n_0 : STD_LOGIC;
  signal W_54_7_i_3_n_0 : STD_LOGIC;
  signal W_54_7_i_4_n_0 : STD_LOGIC;
  signal W_54_7_i_5_n_0 : STD_LOGIC;
  signal W_54_7_i_6_n_0 : STD_LOGIC;
  signal W_54_7_i_7_n_0 : STD_LOGIC;
  signal W_54_7_i_8_n_0 : STD_LOGIC;
  signal W_54_7_i_9_n_0 : STD_LOGIC;
  signal W_55_11_i_10_n_0 : STD_LOGIC;
  signal W_55_11_i_11_n_0 : STD_LOGIC;
  signal W_55_11_i_12_n_0 : STD_LOGIC;
  signal W_55_11_i_13_n_0 : STD_LOGIC;
  signal W_55_11_i_14_n_0 : STD_LOGIC;
  signal W_55_11_i_15_n_0 : STD_LOGIC;
  signal W_55_11_i_16_n_0 : STD_LOGIC;
  signal W_55_11_i_17_n_0 : STD_LOGIC;
  signal W_55_11_i_2_n_0 : STD_LOGIC;
  signal W_55_11_i_3_n_0 : STD_LOGIC;
  signal W_55_11_i_4_n_0 : STD_LOGIC;
  signal W_55_11_i_5_n_0 : STD_LOGIC;
  signal W_55_11_i_6_n_0 : STD_LOGIC;
  signal W_55_11_i_7_n_0 : STD_LOGIC;
  signal W_55_11_i_8_n_0 : STD_LOGIC;
  signal W_55_11_i_9_n_0 : STD_LOGIC;
  signal W_55_15_i_10_n_0 : STD_LOGIC;
  signal W_55_15_i_11_n_0 : STD_LOGIC;
  signal W_55_15_i_12_n_0 : STD_LOGIC;
  signal W_55_15_i_13_n_0 : STD_LOGIC;
  signal W_55_15_i_14_n_0 : STD_LOGIC;
  signal W_55_15_i_15_n_0 : STD_LOGIC;
  signal W_55_15_i_16_n_0 : STD_LOGIC;
  signal W_55_15_i_17_n_0 : STD_LOGIC;
  signal W_55_15_i_2_n_0 : STD_LOGIC;
  signal W_55_15_i_3_n_0 : STD_LOGIC;
  signal W_55_15_i_4_n_0 : STD_LOGIC;
  signal W_55_15_i_5_n_0 : STD_LOGIC;
  signal W_55_15_i_6_n_0 : STD_LOGIC;
  signal W_55_15_i_7_n_0 : STD_LOGIC;
  signal W_55_15_i_8_n_0 : STD_LOGIC;
  signal W_55_15_i_9_n_0 : STD_LOGIC;
  signal W_55_19_i_10_n_0 : STD_LOGIC;
  signal W_55_19_i_11_n_0 : STD_LOGIC;
  signal W_55_19_i_12_n_0 : STD_LOGIC;
  signal W_55_19_i_13_n_0 : STD_LOGIC;
  signal W_55_19_i_14_n_0 : STD_LOGIC;
  signal W_55_19_i_15_n_0 : STD_LOGIC;
  signal W_55_19_i_16_n_0 : STD_LOGIC;
  signal W_55_19_i_17_n_0 : STD_LOGIC;
  signal W_55_19_i_2_n_0 : STD_LOGIC;
  signal W_55_19_i_3_n_0 : STD_LOGIC;
  signal W_55_19_i_4_n_0 : STD_LOGIC;
  signal W_55_19_i_5_n_0 : STD_LOGIC;
  signal W_55_19_i_6_n_0 : STD_LOGIC;
  signal W_55_19_i_7_n_0 : STD_LOGIC;
  signal W_55_19_i_8_n_0 : STD_LOGIC;
  signal W_55_19_i_9_n_0 : STD_LOGIC;
  signal W_55_23_i_10_n_0 : STD_LOGIC;
  signal W_55_23_i_11_n_0 : STD_LOGIC;
  signal W_55_23_i_12_n_0 : STD_LOGIC;
  signal W_55_23_i_13_n_0 : STD_LOGIC;
  signal W_55_23_i_14_n_0 : STD_LOGIC;
  signal W_55_23_i_15_n_0 : STD_LOGIC;
  signal W_55_23_i_16_n_0 : STD_LOGIC;
  signal W_55_23_i_17_n_0 : STD_LOGIC;
  signal W_55_23_i_2_n_0 : STD_LOGIC;
  signal W_55_23_i_3_n_0 : STD_LOGIC;
  signal W_55_23_i_4_n_0 : STD_LOGIC;
  signal W_55_23_i_5_n_0 : STD_LOGIC;
  signal W_55_23_i_6_n_0 : STD_LOGIC;
  signal W_55_23_i_7_n_0 : STD_LOGIC;
  signal W_55_23_i_8_n_0 : STD_LOGIC;
  signal W_55_23_i_9_n_0 : STD_LOGIC;
  signal W_55_27_i_10_n_0 : STD_LOGIC;
  signal W_55_27_i_11_n_0 : STD_LOGIC;
  signal W_55_27_i_12_n_0 : STD_LOGIC;
  signal W_55_27_i_13_n_0 : STD_LOGIC;
  signal W_55_27_i_14_n_0 : STD_LOGIC;
  signal W_55_27_i_15_n_0 : STD_LOGIC;
  signal W_55_27_i_16_n_0 : STD_LOGIC;
  signal W_55_27_i_17_n_0 : STD_LOGIC;
  signal W_55_27_i_2_n_0 : STD_LOGIC;
  signal W_55_27_i_3_n_0 : STD_LOGIC;
  signal W_55_27_i_4_n_0 : STD_LOGIC;
  signal W_55_27_i_5_n_0 : STD_LOGIC;
  signal W_55_27_i_6_n_0 : STD_LOGIC;
  signal W_55_27_i_7_n_0 : STD_LOGIC;
  signal W_55_27_i_8_n_0 : STD_LOGIC;
  signal W_55_27_i_9_n_0 : STD_LOGIC;
  signal W_55_31_i_10_n_0 : STD_LOGIC;
  signal W_55_31_i_11_n_0 : STD_LOGIC;
  signal W_55_31_i_12_n_0 : STD_LOGIC;
  signal W_55_31_i_13_n_0 : STD_LOGIC;
  signal W_55_31_i_14_n_0 : STD_LOGIC;
  signal W_55_31_i_15_n_0 : STD_LOGIC;
  signal W_55_31_i_17_n_0 : STD_LOGIC;
  signal W_55_31_i_19_n_0 : STD_LOGIC;
  signal W_55_31_i_2_n_0 : STD_LOGIC;
  signal W_55_31_i_3_n_0 : STD_LOGIC;
  signal W_55_31_i_4_n_0 : STD_LOGIC;
  signal W_55_31_i_5_n_0 : STD_LOGIC;
  signal W_55_31_i_6_n_0 : STD_LOGIC;
  signal W_55_31_i_7_n_0 : STD_LOGIC;
  signal W_55_31_i_8_n_0 : STD_LOGIC;
  signal W_55_31_i_9_n_0 : STD_LOGIC;
  signal W_55_3_i_10_n_0 : STD_LOGIC;
  signal W_55_3_i_11_n_0 : STD_LOGIC;
  signal W_55_3_i_15_n_0 : STD_LOGIC;
  signal W_55_3_i_2_n_0 : STD_LOGIC;
  signal W_55_3_i_3_n_0 : STD_LOGIC;
  signal W_55_3_i_4_n_0 : STD_LOGIC;
  signal W_55_3_i_5_n_0 : STD_LOGIC;
  signal W_55_3_i_6_n_0 : STD_LOGIC;
  signal W_55_3_i_7_n_0 : STD_LOGIC;
  signal W_55_3_i_8_n_0 : STD_LOGIC;
  signal W_55_3_i_9_n_0 : STD_LOGIC;
  signal W_55_7_i_10_n_0 : STD_LOGIC;
  signal W_55_7_i_11_n_0 : STD_LOGIC;
  signal W_55_7_i_12_n_0 : STD_LOGIC;
  signal W_55_7_i_13_n_0 : STD_LOGIC;
  signal W_55_7_i_14_n_0 : STD_LOGIC;
  signal W_55_7_i_15_n_0 : STD_LOGIC;
  signal W_55_7_i_16_n_0 : STD_LOGIC;
  signal W_55_7_i_17_n_0 : STD_LOGIC;
  signal W_55_7_i_2_n_0 : STD_LOGIC;
  signal W_55_7_i_3_n_0 : STD_LOGIC;
  signal W_55_7_i_4_n_0 : STD_LOGIC;
  signal W_55_7_i_5_n_0 : STD_LOGIC;
  signal W_55_7_i_6_n_0 : STD_LOGIC;
  signal W_55_7_i_7_n_0 : STD_LOGIC;
  signal W_55_7_i_8_n_0 : STD_LOGIC;
  signal W_55_7_i_9_n_0 : STD_LOGIC;
  signal W_56_11_i_10_n_0 : STD_LOGIC;
  signal W_56_11_i_11_n_0 : STD_LOGIC;
  signal W_56_11_i_12_n_0 : STD_LOGIC;
  signal W_56_11_i_13_n_0 : STD_LOGIC;
  signal W_56_11_i_14_n_0 : STD_LOGIC;
  signal W_56_11_i_15_n_0 : STD_LOGIC;
  signal W_56_11_i_16_n_0 : STD_LOGIC;
  signal W_56_11_i_17_n_0 : STD_LOGIC;
  signal W_56_11_i_2_n_0 : STD_LOGIC;
  signal W_56_11_i_3_n_0 : STD_LOGIC;
  signal W_56_11_i_4_n_0 : STD_LOGIC;
  signal W_56_11_i_5_n_0 : STD_LOGIC;
  signal W_56_11_i_6_n_0 : STD_LOGIC;
  signal W_56_11_i_7_n_0 : STD_LOGIC;
  signal W_56_11_i_8_n_0 : STD_LOGIC;
  signal W_56_11_i_9_n_0 : STD_LOGIC;
  signal W_56_15_i_10_n_0 : STD_LOGIC;
  signal W_56_15_i_11_n_0 : STD_LOGIC;
  signal W_56_15_i_12_n_0 : STD_LOGIC;
  signal W_56_15_i_13_n_0 : STD_LOGIC;
  signal W_56_15_i_14_n_0 : STD_LOGIC;
  signal W_56_15_i_15_n_0 : STD_LOGIC;
  signal W_56_15_i_16_n_0 : STD_LOGIC;
  signal W_56_15_i_17_n_0 : STD_LOGIC;
  signal W_56_15_i_2_n_0 : STD_LOGIC;
  signal W_56_15_i_3_n_0 : STD_LOGIC;
  signal W_56_15_i_4_n_0 : STD_LOGIC;
  signal W_56_15_i_5_n_0 : STD_LOGIC;
  signal W_56_15_i_6_n_0 : STD_LOGIC;
  signal W_56_15_i_7_n_0 : STD_LOGIC;
  signal W_56_15_i_8_n_0 : STD_LOGIC;
  signal W_56_15_i_9_n_0 : STD_LOGIC;
  signal W_56_19_i_10_n_0 : STD_LOGIC;
  signal W_56_19_i_11_n_0 : STD_LOGIC;
  signal W_56_19_i_12_n_0 : STD_LOGIC;
  signal W_56_19_i_13_n_0 : STD_LOGIC;
  signal W_56_19_i_14_n_0 : STD_LOGIC;
  signal W_56_19_i_15_n_0 : STD_LOGIC;
  signal W_56_19_i_16_n_0 : STD_LOGIC;
  signal W_56_19_i_17_n_0 : STD_LOGIC;
  signal W_56_19_i_2_n_0 : STD_LOGIC;
  signal W_56_19_i_3_n_0 : STD_LOGIC;
  signal W_56_19_i_4_n_0 : STD_LOGIC;
  signal W_56_19_i_5_n_0 : STD_LOGIC;
  signal W_56_19_i_6_n_0 : STD_LOGIC;
  signal W_56_19_i_7_n_0 : STD_LOGIC;
  signal W_56_19_i_8_n_0 : STD_LOGIC;
  signal W_56_19_i_9_n_0 : STD_LOGIC;
  signal W_56_23_i_10_n_0 : STD_LOGIC;
  signal W_56_23_i_11_n_0 : STD_LOGIC;
  signal W_56_23_i_12_n_0 : STD_LOGIC;
  signal W_56_23_i_13_n_0 : STD_LOGIC;
  signal W_56_23_i_14_n_0 : STD_LOGIC;
  signal W_56_23_i_15_n_0 : STD_LOGIC;
  signal W_56_23_i_16_n_0 : STD_LOGIC;
  signal W_56_23_i_17_n_0 : STD_LOGIC;
  signal W_56_23_i_2_n_0 : STD_LOGIC;
  signal W_56_23_i_3_n_0 : STD_LOGIC;
  signal W_56_23_i_4_n_0 : STD_LOGIC;
  signal W_56_23_i_5_n_0 : STD_LOGIC;
  signal W_56_23_i_6_n_0 : STD_LOGIC;
  signal W_56_23_i_7_n_0 : STD_LOGIC;
  signal W_56_23_i_8_n_0 : STD_LOGIC;
  signal W_56_23_i_9_n_0 : STD_LOGIC;
  signal W_56_27_i_10_n_0 : STD_LOGIC;
  signal W_56_27_i_11_n_0 : STD_LOGIC;
  signal W_56_27_i_12_n_0 : STD_LOGIC;
  signal W_56_27_i_13_n_0 : STD_LOGIC;
  signal W_56_27_i_14_n_0 : STD_LOGIC;
  signal W_56_27_i_15_n_0 : STD_LOGIC;
  signal W_56_27_i_16_n_0 : STD_LOGIC;
  signal W_56_27_i_17_n_0 : STD_LOGIC;
  signal W_56_27_i_2_n_0 : STD_LOGIC;
  signal W_56_27_i_3_n_0 : STD_LOGIC;
  signal W_56_27_i_4_n_0 : STD_LOGIC;
  signal W_56_27_i_5_n_0 : STD_LOGIC;
  signal W_56_27_i_6_n_0 : STD_LOGIC;
  signal W_56_27_i_7_n_0 : STD_LOGIC;
  signal W_56_27_i_8_n_0 : STD_LOGIC;
  signal W_56_27_i_9_n_0 : STD_LOGIC;
  signal W_56_31_i_10_n_0 : STD_LOGIC;
  signal W_56_31_i_11_n_0 : STD_LOGIC;
  signal W_56_31_i_12_n_0 : STD_LOGIC;
  signal W_56_31_i_13_n_0 : STD_LOGIC;
  signal W_56_31_i_14_n_0 : STD_LOGIC;
  signal W_56_31_i_15_n_0 : STD_LOGIC;
  signal W_56_31_i_17_n_0 : STD_LOGIC;
  signal W_56_31_i_19_n_0 : STD_LOGIC;
  signal W_56_31_i_2_n_0 : STD_LOGIC;
  signal W_56_31_i_3_n_0 : STD_LOGIC;
  signal W_56_31_i_4_n_0 : STD_LOGIC;
  signal W_56_31_i_5_n_0 : STD_LOGIC;
  signal W_56_31_i_6_n_0 : STD_LOGIC;
  signal W_56_31_i_7_n_0 : STD_LOGIC;
  signal W_56_31_i_8_n_0 : STD_LOGIC;
  signal W_56_31_i_9_n_0 : STD_LOGIC;
  signal W_56_3_i_10_n_0 : STD_LOGIC;
  signal W_56_3_i_11_n_0 : STD_LOGIC;
  signal W_56_3_i_15_n_0 : STD_LOGIC;
  signal W_56_3_i_2_n_0 : STD_LOGIC;
  signal W_56_3_i_3_n_0 : STD_LOGIC;
  signal W_56_3_i_4_n_0 : STD_LOGIC;
  signal W_56_3_i_5_n_0 : STD_LOGIC;
  signal W_56_3_i_6_n_0 : STD_LOGIC;
  signal W_56_3_i_7_n_0 : STD_LOGIC;
  signal W_56_3_i_8_n_0 : STD_LOGIC;
  signal W_56_3_i_9_n_0 : STD_LOGIC;
  signal W_56_7_i_10_n_0 : STD_LOGIC;
  signal W_56_7_i_11_n_0 : STD_LOGIC;
  signal W_56_7_i_12_n_0 : STD_LOGIC;
  signal W_56_7_i_13_n_0 : STD_LOGIC;
  signal W_56_7_i_14_n_0 : STD_LOGIC;
  signal W_56_7_i_15_n_0 : STD_LOGIC;
  signal W_56_7_i_16_n_0 : STD_LOGIC;
  signal W_56_7_i_17_n_0 : STD_LOGIC;
  signal W_56_7_i_2_n_0 : STD_LOGIC;
  signal W_56_7_i_3_n_0 : STD_LOGIC;
  signal W_56_7_i_4_n_0 : STD_LOGIC;
  signal W_56_7_i_5_n_0 : STD_LOGIC;
  signal W_56_7_i_6_n_0 : STD_LOGIC;
  signal W_56_7_i_7_n_0 : STD_LOGIC;
  signal W_56_7_i_8_n_0 : STD_LOGIC;
  signal W_56_7_i_9_n_0 : STD_LOGIC;
  signal W_57_11_i_10_n_0 : STD_LOGIC;
  signal W_57_11_i_11_n_0 : STD_LOGIC;
  signal W_57_11_i_12_n_0 : STD_LOGIC;
  signal W_57_11_i_13_n_0 : STD_LOGIC;
  signal W_57_11_i_14_n_0 : STD_LOGIC;
  signal W_57_11_i_15_n_0 : STD_LOGIC;
  signal W_57_11_i_16_n_0 : STD_LOGIC;
  signal W_57_11_i_17_n_0 : STD_LOGIC;
  signal W_57_11_i_2_n_0 : STD_LOGIC;
  signal W_57_11_i_3_n_0 : STD_LOGIC;
  signal W_57_11_i_4_n_0 : STD_LOGIC;
  signal W_57_11_i_5_n_0 : STD_LOGIC;
  signal W_57_11_i_6_n_0 : STD_LOGIC;
  signal W_57_11_i_7_n_0 : STD_LOGIC;
  signal W_57_11_i_8_n_0 : STD_LOGIC;
  signal W_57_11_i_9_n_0 : STD_LOGIC;
  signal W_57_15_i_10_n_0 : STD_LOGIC;
  signal W_57_15_i_11_n_0 : STD_LOGIC;
  signal W_57_15_i_12_n_0 : STD_LOGIC;
  signal W_57_15_i_13_n_0 : STD_LOGIC;
  signal W_57_15_i_14_n_0 : STD_LOGIC;
  signal W_57_15_i_15_n_0 : STD_LOGIC;
  signal W_57_15_i_16_n_0 : STD_LOGIC;
  signal W_57_15_i_17_n_0 : STD_LOGIC;
  signal W_57_15_i_2_n_0 : STD_LOGIC;
  signal W_57_15_i_3_n_0 : STD_LOGIC;
  signal W_57_15_i_4_n_0 : STD_LOGIC;
  signal W_57_15_i_5_n_0 : STD_LOGIC;
  signal W_57_15_i_6_n_0 : STD_LOGIC;
  signal W_57_15_i_7_n_0 : STD_LOGIC;
  signal W_57_15_i_8_n_0 : STD_LOGIC;
  signal W_57_15_i_9_n_0 : STD_LOGIC;
  signal W_57_19_i_10_n_0 : STD_LOGIC;
  signal W_57_19_i_11_n_0 : STD_LOGIC;
  signal W_57_19_i_12_n_0 : STD_LOGIC;
  signal W_57_19_i_13_n_0 : STD_LOGIC;
  signal W_57_19_i_14_n_0 : STD_LOGIC;
  signal W_57_19_i_15_n_0 : STD_LOGIC;
  signal W_57_19_i_16_n_0 : STD_LOGIC;
  signal W_57_19_i_17_n_0 : STD_LOGIC;
  signal W_57_19_i_2_n_0 : STD_LOGIC;
  signal W_57_19_i_3_n_0 : STD_LOGIC;
  signal W_57_19_i_4_n_0 : STD_LOGIC;
  signal W_57_19_i_5_n_0 : STD_LOGIC;
  signal W_57_19_i_6_n_0 : STD_LOGIC;
  signal W_57_19_i_7_n_0 : STD_LOGIC;
  signal W_57_19_i_8_n_0 : STD_LOGIC;
  signal W_57_19_i_9_n_0 : STD_LOGIC;
  signal W_57_23_i_10_n_0 : STD_LOGIC;
  signal W_57_23_i_11_n_0 : STD_LOGIC;
  signal W_57_23_i_12_n_0 : STD_LOGIC;
  signal W_57_23_i_13_n_0 : STD_LOGIC;
  signal W_57_23_i_14_n_0 : STD_LOGIC;
  signal W_57_23_i_15_n_0 : STD_LOGIC;
  signal W_57_23_i_16_n_0 : STD_LOGIC;
  signal W_57_23_i_17_n_0 : STD_LOGIC;
  signal W_57_23_i_2_n_0 : STD_LOGIC;
  signal W_57_23_i_3_n_0 : STD_LOGIC;
  signal W_57_23_i_4_n_0 : STD_LOGIC;
  signal W_57_23_i_5_n_0 : STD_LOGIC;
  signal W_57_23_i_6_n_0 : STD_LOGIC;
  signal W_57_23_i_7_n_0 : STD_LOGIC;
  signal W_57_23_i_8_n_0 : STD_LOGIC;
  signal W_57_23_i_9_n_0 : STD_LOGIC;
  signal W_57_27_i_10_n_0 : STD_LOGIC;
  signal W_57_27_i_11_n_0 : STD_LOGIC;
  signal W_57_27_i_12_n_0 : STD_LOGIC;
  signal W_57_27_i_13_n_0 : STD_LOGIC;
  signal W_57_27_i_14_n_0 : STD_LOGIC;
  signal W_57_27_i_15_n_0 : STD_LOGIC;
  signal W_57_27_i_16_n_0 : STD_LOGIC;
  signal W_57_27_i_17_n_0 : STD_LOGIC;
  signal W_57_27_i_2_n_0 : STD_LOGIC;
  signal W_57_27_i_3_n_0 : STD_LOGIC;
  signal W_57_27_i_4_n_0 : STD_LOGIC;
  signal W_57_27_i_5_n_0 : STD_LOGIC;
  signal W_57_27_i_6_n_0 : STD_LOGIC;
  signal W_57_27_i_7_n_0 : STD_LOGIC;
  signal W_57_27_i_8_n_0 : STD_LOGIC;
  signal W_57_27_i_9_n_0 : STD_LOGIC;
  signal W_57_31_i_10_n_0 : STD_LOGIC;
  signal W_57_31_i_11_n_0 : STD_LOGIC;
  signal W_57_31_i_12_n_0 : STD_LOGIC;
  signal W_57_31_i_13_n_0 : STD_LOGIC;
  signal W_57_31_i_14_n_0 : STD_LOGIC;
  signal W_57_31_i_15_n_0 : STD_LOGIC;
  signal W_57_31_i_17_n_0 : STD_LOGIC;
  signal W_57_31_i_19_n_0 : STD_LOGIC;
  signal W_57_31_i_2_n_0 : STD_LOGIC;
  signal W_57_31_i_3_n_0 : STD_LOGIC;
  signal W_57_31_i_4_n_0 : STD_LOGIC;
  signal W_57_31_i_5_n_0 : STD_LOGIC;
  signal W_57_31_i_6_n_0 : STD_LOGIC;
  signal W_57_31_i_7_n_0 : STD_LOGIC;
  signal W_57_31_i_8_n_0 : STD_LOGIC;
  signal W_57_31_i_9_n_0 : STD_LOGIC;
  signal W_57_3_i_10_n_0 : STD_LOGIC;
  signal W_57_3_i_11_n_0 : STD_LOGIC;
  signal W_57_3_i_15_n_0 : STD_LOGIC;
  signal W_57_3_i_2_n_0 : STD_LOGIC;
  signal W_57_3_i_3_n_0 : STD_LOGIC;
  signal W_57_3_i_4_n_0 : STD_LOGIC;
  signal W_57_3_i_5_n_0 : STD_LOGIC;
  signal W_57_3_i_6_n_0 : STD_LOGIC;
  signal W_57_3_i_7_n_0 : STD_LOGIC;
  signal W_57_3_i_8_n_0 : STD_LOGIC;
  signal W_57_3_i_9_n_0 : STD_LOGIC;
  signal W_57_7_i_10_n_0 : STD_LOGIC;
  signal W_57_7_i_11_n_0 : STD_LOGIC;
  signal W_57_7_i_12_n_0 : STD_LOGIC;
  signal W_57_7_i_13_n_0 : STD_LOGIC;
  signal W_57_7_i_14_n_0 : STD_LOGIC;
  signal W_57_7_i_15_n_0 : STD_LOGIC;
  signal W_57_7_i_16_n_0 : STD_LOGIC;
  signal W_57_7_i_17_n_0 : STD_LOGIC;
  signal W_57_7_i_2_n_0 : STD_LOGIC;
  signal W_57_7_i_3_n_0 : STD_LOGIC;
  signal W_57_7_i_4_n_0 : STD_LOGIC;
  signal W_57_7_i_5_n_0 : STD_LOGIC;
  signal W_57_7_i_6_n_0 : STD_LOGIC;
  signal W_57_7_i_7_n_0 : STD_LOGIC;
  signal W_57_7_i_8_n_0 : STD_LOGIC;
  signal W_57_7_i_9_n_0 : STD_LOGIC;
  signal W_58_11_i_10_n_0 : STD_LOGIC;
  signal W_58_11_i_11_n_0 : STD_LOGIC;
  signal W_58_11_i_12_n_0 : STD_LOGIC;
  signal W_58_11_i_13_n_0 : STD_LOGIC;
  signal W_58_11_i_14_n_0 : STD_LOGIC;
  signal W_58_11_i_15_n_0 : STD_LOGIC;
  signal W_58_11_i_16_n_0 : STD_LOGIC;
  signal W_58_11_i_17_n_0 : STD_LOGIC;
  signal W_58_11_i_2_n_0 : STD_LOGIC;
  signal W_58_11_i_3_n_0 : STD_LOGIC;
  signal W_58_11_i_4_n_0 : STD_LOGIC;
  signal W_58_11_i_5_n_0 : STD_LOGIC;
  signal W_58_11_i_6_n_0 : STD_LOGIC;
  signal W_58_11_i_7_n_0 : STD_LOGIC;
  signal W_58_11_i_8_n_0 : STD_LOGIC;
  signal W_58_11_i_9_n_0 : STD_LOGIC;
  signal W_58_15_i_10_n_0 : STD_LOGIC;
  signal W_58_15_i_11_n_0 : STD_LOGIC;
  signal W_58_15_i_12_n_0 : STD_LOGIC;
  signal W_58_15_i_13_n_0 : STD_LOGIC;
  signal W_58_15_i_14_n_0 : STD_LOGIC;
  signal W_58_15_i_15_n_0 : STD_LOGIC;
  signal W_58_15_i_16_n_0 : STD_LOGIC;
  signal W_58_15_i_17_n_0 : STD_LOGIC;
  signal W_58_15_i_2_n_0 : STD_LOGIC;
  signal W_58_15_i_3_n_0 : STD_LOGIC;
  signal W_58_15_i_4_n_0 : STD_LOGIC;
  signal W_58_15_i_5_n_0 : STD_LOGIC;
  signal W_58_15_i_6_n_0 : STD_LOGIC;
  signal W_58_15_i_7_n_0 : STD_LOGIC;
  signal W_58_15_i_8_n_0 : STD_LOGIC;
  signal W_58_15_i_9_n_0 : STD_LOGIC;
  signal W_58_19_i_10_n_0 : STD_LOGIC;
  signal W_58_19_i_11_n_0 : STD_LOGIC;
  signal W_58_19_i_12_n_0 : STD_LOGIC;
  signal W_58_19_i_13_n_0 : STD_LOGIC;
  signal W_58_19_i_14_n_0 : STD_LOGIC;
  signal W_58_19_i_15_n_0 : STD_LOGIC;
  signal W_58_19_i_16_n_0 : STD_LOGIC;
  signal W_58_19_i_17_n_0 : STD_LOGIC;
  signal W_58_19_i_2_n_0 : STD_LOGIC;
  signal W_58_19_i_3_n_0 : STD_LOGIC;
  signal W_58_19_i_4_n_0 : STD_LOGIC;
  signal W_58_19_i_5_n_0 : STD_LOGIC;
  signal W_58_19_i_6_n_0 : STD_LOGIC;
  signal W_58_19_i_7_n_0 : STD_LOGIC;
  signal W_58_19_i_8_n_0 : STD_LOGIC;
  signal W_58_19_i_9_n_0 : STD_LOGIC;
  signal W_58_23_i_10_n_0 : STD_LOGIC;
  signal W_58_23_i_11_n_0 : STD_LOGIC;
  signal W_58_23_i_12_n_0 : STD_LOGIC;
  signal W_58_23_i_13_n_0 : STD_LOGIC;
  signal W_58_23_i_14_n_0 : STD_LOGIC;
  signal W_58_23_i_15_n_0 : STD_LOGIC;
  signal W_58_23_i_16_n_0 : STD_LOGIC;
  signal W_58_23_i_17_n_0 : STD_LOGIC;
  signal W_58_23_i_2_n_0 : STD_LOGIC;
  signal W_58_23_i_3_n_0 : STD_LOGIC;
  signal W_58_23_i_4_n_0 : STD_LOGIC;
  signal W_58_23_i_5_n_0 : STD_LOGIC;
  signal W_58_23_i_6_n_0 : STD_LOGIC;
  signal W_58_23_i_7_n_0 : STD_LOGIC;
  signal W_58_23_i_8_n_0 : STD_LOGIC;
  signal W_58_23_i_9_n_0 : STD_LOGIC;
  signal W_58_27_i_10_n_0 : STD_LOGIC;
  signal W_58_27_i_11_n_0 : STD_LOGIC;
  signal W_58_27_i_12_n_0 : STD_LOGIC;
  signal W_58_27_i_13_n_0 : STD_LOGIC;
  signal W_58_27_i_14_n_0 : STD_LOGIC;
  signal W_58_27_i_15_n_0 : STD_LOGIC;
  signal W_58_27_i_16_n_0 : STD_LOGIC;
  signal W_58_27_i_17_n_0 : STD_LOGIC;
  signal W_58_27_i_2_n_0 : STD_LOGIC;
  signal W_58_27_i_3_n_0 : STD_LOGIC;
  signal W_58_27_i_4_n_0 : STD_LOGIC;
  signal W_58_27_i_5_n_0 : STD_LOGIC;
  signal W_58_27_i_6_n_0 : STD_LOGIC;
  signal W_58_27_i_7_n_0 : STD_LOGIC;
  signal W_58_27_i_8_n_0 : STD_LOGIC;
  signal W_58_27_i_9_n_0 : STD_LOGIC;
  signal W_58_31_i_10_n_0 : STD_LOGIC;
  signal W_58_31_i_11_n_0 : STD_LOGIC;
  signal W_58_31_i_12_n_0 : STD_LOGIC;
  signal W_58_31_i_13_n_0 : STD_LOGIC;
  signal W_58_31_i_14_n_0 : STD_LOGIC;
  signal W_58_31_i_15_n_0 : STD_LOGIC;
  signal W_58_31_i_17_n_0 : STD_LOGIC;
  signal W_58_31_i_19_n_0 : STD_LOGIC;
  signal W_58_31_i_2_n_0 : STD_LOGIC;
  signal W_58_31_i_3_n_0 : STD_LOGIC;
  signal W_58_31_i_4_n_0 : STD_LOGIC;
  signal W_58_31_i_5_n_0 : STD_LOGIC;
  signal W_58_31_i_6_n_0 : STD_LOGIC;
  signal W_58_31_i_7_n_0 : STD_LOGIC;
  signal W_58_31_i_8_n_0 : STD_LOGIC;
  signal W_58_31_i_9_n_0 : STD_LOGIC;
  signal W_58_3_i_10_n_0 : STD_LOGIC;
  signal W_58_3_i_11_n_0 : STD_LOGIC;
  signal W_58_3_i_15_n_0 : STD_LOGIC;
  signal W_58_3_i_2_n_0 : STD_LOGIC;
  signal W_58_3_i_3_n_0 : STD_LOGIC;
  signal W_58_3_i_4_n_0 : STD_LOGIC;
  signal W_58_3_i_5_n_0 : STD_LOGIC;
  signal W_58_3_i_6_n_0 : STD_LOGIC;
  signal W_58_3_i_7_n_0 : STD_LOGIC;
  signal W_58_3_i_8_n_0 : STD_LOGIC;
  signal W_58_3_i_9_n_0 : STD_LOGIC;
  signal W_58_7_i_10_n_0 : STD_LOGIC;
  signal W_58_7_i_11_n_0 : STD_LOGIC;
  signal W_58_7_i_12_n_0 : STD_LOGIC;
  signal W_58_7_i_13_n_0 : STD_LOGIC;
  signal W_58_7_i_14_n_0 : STD_LOGIC;
  signal W_58_7_i_15_n_0 : STD_LOGIC;
  signal W_58_7_i_16_n_0 : STD_LOGIC;
  signal W_58_7_i_17_n_0 : STD_LOGIC;
  signal W_58_7_i_2_n_0 : STD_LOGIC;
  signal W_58_7_i_3_n_0 : STD_LOGIC;
  signal W_58_7_i_4_n_0 : STD_LOGIC;
  signal W_58_7_i_5_n_0 : STD_LOGIC;
  signal W_58_7_i_6_n_0 : STD_LOGIC;
  signal W_58_7_i_7_n_0 : STD_LOGIC;
  signal W_58_7_i_8_n_0 : STD_LOGIC;
  signal W_58_7_i_9_n_0 : STD_LOGIC;
  signal W_59_11_i_10_n_0 : STD_LOGIC;
  signal W_59_11_i_11_n_0 : STD_LOGIC;
  signal W_59_11_i_12_n_0 : STD_LOGIC;
  signal W_59_11_i_13_n_0 : STD_LOGIC;
  signal W_59_11_i_14_n_0 : STD_LOGIC;
  signal W_59_11_i_15_n_0 : STD_LOGIC;
  signal W_59_11_i_16_n_0 : STD_LOGIC;
  signal W_59_11_i_17_n_0 : STD_LOGIC;
  signal W_59_11_i_2_n_0 : STD_LOGIC;
  signal W_59_11_i_3_n_0 : STD_LOGIC;
  signal W_59_11_i_4_n_0 : STD_LOGIC;
  signal W_59_11_i_5_n_0 : STD_LOGIC;
  signal W_59_11_i_6_n_0 : STD_LOGIC;
  signal W_59_11_i_7_n_0 : STD_LOGIC;
  signal W_59_11_i_8_n_0 : STD_LOGIC;
  signal W_59_11_i_9_n_0 : STD_LOGIC;
  signal W_59_15_i_10_n_0 : STD_LOGIC;
  signal W_59_15_i_11_n_0 : STD_LOGIC;
  signal W_59_15_i_12_n_0 : STD_LOGIC;
  signal W_59_15_i_13_n_0 : STD_LOGIC;
  signal W_59_15_i_14_n_0 : STD_LOGIC;
  signal W_59_15_i_15_n_0 : STD_LOGIC;
  signal W_59_15_i_16_n_0 : STD_LOGIC;
  signal W_59_15_i_17_n_0 : STD_LOGIC;
  signal W_59_15_i_2_n_0 : STD_LOGIC;
  signal W_59_15_i_3_n_0 : STD_LOGIC;
  signal W_59_15_i_4_n_0 : STD_LOGIC;
  signal W_59_15_i_5_n_0 : STD_LOGIC;
  signal W_59_15_i_6_n_0 : STD_LOGIC;
  signal W_59_15_i_7_n_0 : STD_LOGIC;
  signal W_59_15_i_8_n_0 : STD_LOGIC;
  signal W_59_15_i_9_n_0 : STD_LOGIC;
  signal W_59_19_i_10_n_0 : STD_LOGIC;
  signal W_59_19_i_11_n_0 : STD_LOGIC;
  signal W_59_19_i_12_n_0 : STD_LOGIC;
  signal W_59_19_i_13_n_0 : STD_LOGIC;
  signal W_59_19_i_14_n_0 : STD_LOGIC;
  signal W_59_19_i_15_n_0 : STD_LOGIC;
  signal W_59_19_i_16_n_0 : STD_LOGIC;
  signal W_59_19_i_17_n_0 : STD_LOGIC;
  signal W_59_19_i_2_n_0 : STD_LOGIC;
  signal W_59_19_i_3_n_0 : STD_LOGIC;
  signal W_59_19_i_4_n_0 : STD_LOGIC;
  signal W_59_19_i_5_n_0 : STD_LOGIC;
  signal W_59_19_i_6_n_0 : STD_LOGIC;
  signal W_59_19_i_7_n_0 : STD_LOGIC;
  signal W_59_19_i_8_n_0 : STD_LOGIC;
  signal W_59_19_i_9_n_0 : STD_LOGIC;
  signal W_59_23_i_10_n_0 : STD_LOGIC;
  signal W_59_23_i_11_n_0 : STD_LOGIC;
  signal W_59_23_i_12_n_0 : STD_LOGIC;
  signal W_59_23_i_13_n_0 : STD_LOGIC;
  signal W_59_23_i_14_n_0 : STD_LOGIC;
  signal W_59_23_i_15_n_0 : STD_LOGIC;
  signal W_59_23_i_16_n_0 : STD_LOGIC;
  signal W_59_23_i_17_n_0 : STD_LOGIC;
  signal W_59_23_i_2_n_0 : STD_LOGIC;
  signal W_59_23_i_3_n_0 : STD_LOGIC;
  signal W_59_23_i_4_n_0 : STD_LOGIC;
  signal W_59_23_i_5_n_0 : STD_LOGIC;
  signal W_59_23_i_6_n_0 : STD_LOGIC;
  signal W_59_23_i_7_n_0 : STD_LOGIC;
  signal W_59_23_i_8_n_0 : STD_LOGIC;
  signal W_59_23_i_9_n_0 : STD_LOGIC;
  signal W_59_27_i_10_n_0 : STD_LOGIC;
  signal W_59_27_i_11_n_0 : STD_LOGIC;
  signal W_59_27_i_12_n_0 : STD_LOGIC;
  signal W_59_27_i_13_n_0 : STD_LOGIC;
  signal W_59_27_i_14_n_0 : STD_LOGIC;
  signal W_59_27_i_15_n_0 : STD_LOGIC;
  signal W_59_27_i_16_n_0 : STD_LOGIC;
  signal W_59_27_i_17_n_0 : STD_LOGIC;
  signal W_59_27_i_2_n_0 : STD_LOGIC;
  signal W_59_27_i_3_n_0 : STD_LOGIC;
  signal W_59_27_i_4_n_0 : STD_LOGIC;
  signal W_59_27_i_5_n_0 : STD_LOGIC;
  signal W_59_27_i_6_n_0 : STD_LOGIC;
  signal W_59_27_i_7_n_0 : STD_LOGIC;
  signal W_59_27_i_8_n_0 : STD_LOGIC;
  signal W_59_27_i_9_n_0 : STD_LOGIC;
  signal W_59_31_i_10_n_0 : STD_LOGIC;
  signal W_59_31_i_11_n_0 : STD_LOGIC;
  signal W_59_31_i_12_n_0 : STD_LOGIC;
  signal W_59_31_i_13_n_0 : STD_LOGIC;
  signal W_59_31_i_14_n_0 : STD_LOGIC;
  signal W_59_31_i_15_n_0 : STD_LOGIC;
  signal W_59_31_i_17_n_0 : STD_LOGIC;
  signal W_59_31_i_19_n_0 : STD_LOGIC;
  signal W_59_31_i_2_n_0 : STD_LOGIC;
  signal W_59_31_i_3_n_0 : STD_LOGIC;
  signal W_59_31_i_4_n_0 : STD_LOGIC;
  signal W_59_31_i_5_n_0 : STD_LOGIC;
  signal W_59_31_i_6_n_0 : STD_LOGIC;
  signal W_59_31_i_7_n_0 : STD_LOGIC;
  signal W_59_31_i_8_n_0 : STD_LOGIC;
  signal W_59_31_i_9_n_0 : STD_LOGIC;
  signal W_59_3_i_10_n_0 : STD_LOGIC;
  signal W_59_3_i_11_n_0 : STD_LOGIC;
  signal W_59_3_i_15_n_0 : STD_LOGIC;
  signal W_59_3_i_2_n_0 : STD_LOGIC;
  signal W_59_3_i_3_n_0 : STD_LOGIC;
  signal W_59_3_i_4_n_0 : STD_LOGIC;
  signal W_59_3_i_5_n_0 : STD_LOGIC;
  signal W_59_3_i_6_n_0 : STD_LOGIC;
  signal W_59_3_i_7_n_0 : STD_LOGIC;
  signal W_59_3_i_8_n_0 : STD_LOGIC;
  signal W_59_3_i_9_n_0 : STD_LOGIC;
  signal W_59_7_i_10_n_0 : STD_LOGIC;
  signal W_59_7_i_11_n_0 : STD_LOGIC;
  signal W_59_7_i_12_n_0 : STD_LOGIC;
  signal W_59_7_i_13_n_0 : STD_LOGIC;
  signal W_59_7_i_14_n_0 : STD_LOGIC;
  signal W_59_7_i_15_n_0 : STD_LOGIC;
  signal W_59_7_i_16_n_0 : STD_LOGIC;
  signal W_59_7_i_17_n_0 : STD_LOGIC;
  signal W_59_7_i_2_n_0 : STD_LOGIC;
  signal W_59_7_i_3_n_0 : STD_LOGIC;
  signal W_59_7_i_4_n_0 : STD_LOGIC;
  signal W_59_7_i_5_n_0 : STD_LOGIC;
  signal W_59_7_i_6_n_0 : STD_LOGIC;
  signal W_59_7_i_7_n_0 : STD_LOGIC;
  signal W_59_7_i_8_n_0 : STD_LOGIC;
  signal W_59_7_i_9_n_0 : STD_LOGIC;
  signal W_60_11_i_10_n_0 : STD_LOGIC;
  signal W_60_11_i_11_n_0 : STD_LOGIC;
  signal W_60_11_i_12_n_0 : STD_LOGIC;
  signal W_60_11_i_13_n_0 : STD_LOGIC;
  signal W_60_11_i_14_n_0 : STD_LOGIC;
  signal W_60_11_i_15_n_0 : STD_LOGIC;
  signal W_60_11_i_16_n_0 : STD_LOGIC;
  signal W_60_11_i_17_n_0 : STD_LOGIC;
  signal W_60_11_i_2_n_0 : STD_LOGIC;
  signal W_60_11_i_3_n_0 : STD_LOGIC;
  signal W_60_11_i_4_n_0 : STD_LOGIC;
  signal W_60_11_i_5_n_0 : STD_LOGIC;
  signal W_60_11_i_6_n_0 : STD_LOGIC;
  signal W_60_11_i_7_n_0 : STD_LOGIC;
  signal W_60_11_i_8_n_0 : STD_LOGIC;
  signal W_60_11_i_9_n_0 : STD_LOGIC;
  signal W_60_15_i_10_n_0 : STD_LOGIC;
  signal W_60_15_i_11_n_0 : STD_LOGIC;
  signal W_60_15_i_12_n_0 : STD_LOGIC;
  signal W_60_15_i_13_n_0 : STD_LOGIC;
  signal W_60_15_i_14_n_0 : STD_LOGIC;
  signal W_60_15_i_15_n_0 : STD_LOGIC;
  signal W_60_15_i_16_n_0 : STD_LOGIC;
  signal W_60_15_i_17_n_0 : STD_LOGIC;
  signal W_60_15_i_2_n_0 : STD_LOGIC;
  signal W_60_15_i_3_n_0 : STD_LOGIC;
  signal W_60_15_i_4_n_0 : STD_LOGIC;
  signal W_60_15_i_5_n_0 : STD_LOGIC;
  signal W_60_15_i_6_n_0 : STD_LOGIC;
  signal W_60_15_i_7_n_0 : STD_LOGIC;
  signal W_60_15_i_8_n_0 : STD_LOGIC;
  signal W_60_15_i_9_n_0 : STD_LOGIC;
  signal W_60_19_i_10_n_0 : STD_LOGIC;
  signal W_60_19_i_11_n_0 : STD_LOGIC;
  signal W_60_19_i_12_n_0 : STD_LOGIC;
  signal W_60_19_i_13_n_0 : STD_LOGIC;
  signal W_60_19_i_14_n_0 : STD_LOGIC;
  signal W_60_19_i_15_n_0 : STD_LOGIC;
  signal W_60_19_i_16_n_0 : STD_LOGIC;
  signal W_60_19_i_17_n_0 : STD_LOGIC;
  signal W_60_19_i_2_n_0 : STD_LOGIC;
  signal W_60_19_i_3_n_0 : STD_LOGIC;
  signal W_60_19_i_4_n_0 : STD_LOGIC;
  signal W_60_19_i_5_n_0 : STD_LOGIC;
  signal W_60_19_i_6_n_0 : STD_LOGIC;
  signal W_60_19_i_7_n_0 : STD_LOGIC;
  signal W_60_19_i_8_n_0 : STD_LOGIC;
  signal W_60_19_i_9_n_0 : STD_LOGIC;
  signal W_60_23_i_10_n_0 : STD_LOGIC;
  signal W_60_23_i_11_n_0 : STD_LOGIC;
  signal W_60_23_i_12_n_0 : STD_LOGIC;
  signal W_60_23_i_13_n_0 : STD_LOGIC;
  signal W_60_23_i_14_n_0 : STD_LOGIC;
  signal W_60_23_i_15_n_0 : STD_LOGIC;
  signal W_60_23_i_16_n_0 : STD_LOGIC;
  signal W_60_23_i_17_n_0 : STD_LOGIC;
  signal W_60_23_i_2_n_0 : STD_LOGIC;
  signal W_60_23_i_3_n_0 : STD_LOGIC;
  signal W_60_23_i_4_n_0 : STD_LOGIC;
  signal W_60_23_i_5_n_0 : STD_LOGIC;
  signal W_60_23_i_6_n_0 : STD_LOGIC;
  signal W_60_23_i_7_n_0 : STD_LOGIC;
  signal W_60_23_i_8_n_0 : STD_LOGIC;
  signal W_60_23_i_9_n_0 : STD_LOGIC;
  signal W_60_27_i_10_n_0 : STD_LOGIC;
  signal W_60_27_i_11_n_0 : STD_LOGIC;
  signal W_60_27_i_12_n_0 : STD_LOGIC;
  signal W_60_27_i_13_n_0 : STD_LOGIC;
  signal W_60_27_i_14_n_0 : STD_LOGIC;
  signal W_60_27_i_15_n_0 : STD_LOGIC;
  signal W_60_27_i_16_n_0 : STD_LOGIC;
  signal W_60_27_i_17_n_0 : STD_LOGIC;
  signal W_60_27_i_2_n_0 : STD_LOGIC;
  signal W_60_27_i_3_n_0 : STD_LOGIC;
  signal W_60_27_i_4_n_0 : STD_LOGIC;
  signal W_60_27_i_5_n_0 : STD_LOGIC;
  signal W_60_27_i_6_n_0 : STD_LOGIC;
  signal W_60_27_i_7_n_0 : STD_LOGIC;
  signal W_60_27_i_8_n_0 : STD_LOGIC;
  signal W_60_27_i_9_n_0 : STD_LOGIC;
  signal W_60_31_i_10_n_0 : STD_LOGIC;
  signal W_60_31_i_11_n_0 : STD_LOGIC;
  signal W_60_31_i_12_n_0 : STD_LOGIC;
  signal W_60_31_i_13_n_0 : STD_LOGIC;
  signal W_60_31_i_14_n_0 : STD_LOGIC;
  signal W_60_31_i_15_n_0 : STD_LOGIC;
  signal W_60_31_i_17_n_0 : STD_LOGIC;
  signal W_60_31_i_19_n_0 : STD_LOGIC;
  signal W_60_31_i_2_n_0 : STD_LOGIC;
  signal W_60_31_i_3_n_0 : STD_LOGIC;
  signal W_60_31_i_4_n_0 : STD_LOGIC;
  signal W_60_31_i_5_n_0 : STD_LOGIC;
  signal W_60_31_i_6_n_0 : STD_LOGIC;
  signal W_60_31_i_7_n_0 : STD_LOGIC;
  signal W_60_31_i_8_n_0 : STD_LOGIC;
  signal W_60_31_i_9_n_0 : STD_LOGIC;
  signal W_60_3_i_10_n_0 : STD_LOGIC;
  signal W_60_3_i_11_n_0 : STD_LOGIC;
  signal W_60_3_i_15_n_0 : STD_LOGIC;
  signal W_60_3_i_2_n_0 : STD_LOGIC;
  signal W_60_3_i_3_n_0 : STD_LOGIC;
  signal W_60_3_i_4_n_0 : STD_LOGIC;
  signal W_60_3_i_5_n_0 : STD_LOGIC;
  signal W_60_3_i_6_n_0 : STD_LOGIC;
  signal W_60_3_i_7_n_0 : STD_LOGIC;
  signal W_60_3_i_8_n_0 : STD_LOGIC;
  signal W_60_3_i_9_n_0 : STD_LOGIC;
  signal W_60_7_i_10_n_0 : STD_LOGIC;
  signal W_60_7_i_11_n_0 : STD_LOGIC;
  signal W_60_7_i_12_n_0 : STD_LOGIC;
  signal W_60_7_i_13_n_0 : STD_LOGIC;
  signal W_60_7_i_14_n_0 : STD_LOGIC;
  signal W_60_7_i_15_n_0 : STD_LOGIC;
  signal W_60_7_i_16_n_0 : STD_LOGIC;
  signal W_60_7_i_17_n_0 : STD_LOGIC;
  signal W_60_7_i_2_n_0 : STD_LOGIC;
  signal W_60_7_i_3_n_0 : STD_LOGIC;
  signal W_60_7_i_4_n_0 : STD_LOGIC;
  signal W_60_7_i_5_n_0 : STD_LOGIC;
  signal W_60_7_i_6_n_0 : STD_LOGIC;
  signal W_60_7_i_7_n_0 : STD_LOGIC;
  signal W_60_7_i_8_n_0 : STD_LOGIC;
  signal W_60_7_i_9_n_0 : STD_LOGIC;
  signal W_61_11_i_10_n_0 : STD_LOGIC;
  signal W_61_11_i_11_n_0 : STD_LOGIC;
  signal W_61_11_i_12_n_0 : STD_LOGIC;
  signal W_61_11_i_13_n_0 : STD_LOGIC;
  signal W_61_11_i_14_n_0 : STD_LOGIC;
  signal W_61_11_i_15_n_0 : STD_LOGIC;
  signal W_61_11_i_16_n_0 : STD_LOGIC;
  signal W_61_11_i_17_n_0 : STD_LOGIC;
  signal W_61_11_i_2_n_0 : STD_LOGIC;
  signal W_61_11_i_3_n_0 : STD_LOGIC;
  signal W_61_11_i_4_n_0 : STD_LOGIC;
  signal W_61_11_i_5_n_0 : STD_LOGIC;
  signal W_61_11_i_6_n_0 : STD_LOGIC;
  signal W_61_11_i_7_n_0 : STD_LOGIC;
  signal W_61_11_i_8_n_0 : STD_LOGIC;
  signal W_61_11_i_9_n_0 : STD_LOGIC;
  signal W_61_15_i_10_n_0 : STD_LOGIC;
  signal W_61_15_i_11_n_0 : STD_LOGIC;
  signal W_61_15_i_12_n_0 : STD_LOGIC;
  signal W_61_15_i_13_n_0 : STD_LOGIC;
  signal W_61_15_i_14_n_0 : STD_LOGIC;
  signal W_61_15_i_15_n_0 : STD_LOGIC;
  signal W_61_15_i_16_n_0 : STD_LOGIC;
  signal W_61_15_i_17_n_0 : STD_LOGIC;
  signal W_61_15_i_2_n_0 : STD_LOGIC;
  signal W_61_15_i_3_n_0 : STD_LOGIC;
  signal W_61_15_i_4_n_0 : STD_LOGIC;
  signal W_61_15_i_5_n_0 : STD_LOGIC;
  signal W_61_15_i_6_n_0 : STD_LOGIC;
  signal W_61_15_i_7_n_0 : STD_LOGIC;
  signal W_61_15_i_8_n_0 : STD_LOGIC;
  signal W_61_15_i_9_n_0 : STD_LOGIC;
  signal W_61_19_i_10_n_0 : STD_LOGIC;
  signal W_61_19_i_11_n_0 : STD_LOGIC;
  signal W_61_19_i_12_n_0 : STD_LOGIC;
  signal W_61_19_i_13_n_0 : STD_LOGIC;
  signal W_61_19_i_14_n_0 : STD_LOGIC;
  signal W_61_19_i_15_n_0 : STD_LOGIC;
  signal W_61_19_i_16_n_0 : STD_LOGIC;
  signal W_61_19_i_17_n_0 : STD_LOGIC;
  signal W_61_19_i_2_n_0 : STD_LOGIC;
  signal W_61_19_i_3_n_0 : STD_LOGIC;
  signal W_61_19_i_4_n_0 : STD_LOGIC;
  signal W_61_19_i_5_n_0 : STD_LOGIC;
  signal W_61_19_i_6_n_0 : STD_LOGIC;
  signal W_61_19_i_7_n_0 : STD_LOGIC;
  signal W_61_19_i_8_n_0 : STD_LOGIC;
  signal W_61_19_i_9_n_0 : STD_LOGIC;
  signal W_61_23_i_10_n_0 : STD_LOGIC;
  signal W_61_23_i_11_n_0 : STD_LOGIC;
  signal W_61_23_i_12_n_0 : STD_LOGIC;
  signal W_61_23_i_13_n_0 : STD_LOGIC;
  signal W_61_23_i_14_n_0 : STD_LOGIC;
  signal W_61_23_i_15_n_0 : STD_LOGIC;
  signal W_61_23_i_16_n_0 : STD_LOGIC;
  signal W_61_23_i_17_n_0 : STD_LOGIC;
  signal W_61_23_i_2_n_0 : STD_LOGIC;
  signal W_61_23_i_3_n_0 : STD_LOGIC;
  signal W_61_23_i_4_n_0 : STD_LOGIC;
  signal W_61_23_i_5_n_0 : STD_LOGIC;
  signal W_61_23_i_6_n_0 : STD_LOGIC;
  signal W_61_23_i_7_n_0 : STD_LOGIC;
  signal W_61_23_i_8_n_0 : STD_LOGIC;
  signal W_61_23_i_9_n_0 : STD_LOGIC;
  signal W_61_27_i_10_n_0 : STD_LOGIC;
  signal W_61_27_i_11_n_0 : STD_LOGIC;
  signal W_61_27_i_12_n_0 : STD_LOGIC;
  signal W_61_27_i_13_n_0 : STD_LOGIC;
  signal W_61_27_i_14_n_0 : STD_LOGIC;
  signal W_61_27_i_15_n_0 : STD_LOGIC;
  signal W_61_27_i_16_n_0 : STD_LOGIC;
  signal W_61_27_i_17_n_0 : STD_LOGIC;
  signal W_61_27_i_2_n_0 : STD_LOGIC;
  signal W_61_27_i_3_n_0 : STD_LOGIC;
  signal W_61_27_i_4_n_0 : STD_LOGIC;
  signal W_61_27_i_5_n_0 : STD_LOGIC;
  signal W_61_27_i_6_n_0 : STD_LOGIC;
  signal W_61_27_i_7_n_0 : STD_LOGIC;
  signal W_61_27_i_8_n_0 : STD_LOGIC;
  signal W_61_27_i_9_n_0 : STD_LOGIC;
  signal W_61_31_i_10_n_0 : STD_LOGIC;
  signal W_61_31_i_11_n_0 : STD_LOGIC;
  signal W_61_31_i_12_n_0 : STD_LOGIC;
  signal W_61_31_i_13_n_0 : STD_LOGIC;
  signal W_61_31_i_14_n_0 : STD_LOGIC;
  signal W_61_31_i_15_n_0 : STD_LOGIC;
  signal W_61_31_i_17_n_0 : STD_LOGIC;
  signal W_61_31_i_19_n_0 : STD_LOGIC;
  signal W_61_31_i_2_n_0 : STD_LOGIC;
  signal W_61_31_i_3_n_0 : STD_LOGIC;
  signal W_61_31_i_4_n_0 : STD_LOGIC;
  signal W_61_31_i_5_n_0 : STD_LOGIC;
  signal W_61_31_i_6_n_0 : STD_LOGIC;
  signal W_61_31_i_7_n_0 : STD_LOGIC;
  signal W_61_31_i_8_n_0 : STD_LOGIC;
  signal W_61_31_i_9_n_0 : STD_LOGIC;
  signal W_61_3_i_10_n_0 : STD_LOGIC;
  signal W_61_3_i_11_n_0 : STD_LOGIC;
  signal W_61_3_i_15_n_0 : STD_LOGIC;
  signal W_61_3_i_2_n_0 : STD_LOGIC;
  signal W_61_3_i_3_n_0 : STD_LOGIC;
  signal W_61_3_i_4_n_0 : STD_LOGIC;
  signal W_61_3_i_5_n_0 : STD_LOGIC;
  signal W_61_3_i_6_n_0 : STD_LOGIC;
  signal W_61_3_i_7_n_0 : STD_LOGIC;
  signal W_61_3_i_8_n_0 : STD_LOGIC;
  signal W_61_3_i_9_n_0 : STD_LOGIC;
  signal W_61_7_i_10_n_0 : STD_LOGIC;
  signal W_61_7_i_11_n_0 : STD_LOGIC;
  signal W_61_7_i_12_n_0 : STD_LOGIC;
  signal W_61_7_i_13_n_0 : STD_LOGIC;
  signal W_61_7_i_14_n_0 : STD_LOGIC;
  signal W_61_7_i_15_n_0 : STD_LOGIC;
  signal W_61_7_i_16_n_0 : STD_LOGIC;
  signal W_61_7_i_17_n_0 : STD_LOGIC;
  signal W_61_7_i_2_n_0 : STD_LOGIC;
  signal W_61_7_i_3_n_0 : STD_LOGIC;
  signal W_61_7_i_4_n_0 : STD_LOGIC;
  signal W_61_7_i_5_n_0 : STD_LOGIC;
  signal W_61_7_i_6_n_0 : STD_LOGIC;
  signal W_61_7_i_7_n_0 : STD_LOGIC;
  signal W_61_7_i_8_n_0 : STD_LOGIC;
  signal W_61_7_i_9_n_0 : STD_LOGIC;
  signal W_62_11_i_10_n_0 : STD_LOGIC;
  signal W_62_11_i_11_n_0 : STD_LOGIC;
  signal W_62_11_i_12_n_0 : STD_LOGIC;
  signal W_62_11_i_13_n_0 : STD_LOGIC;
  signal W_62_11_i_14_n_0 : STD_LOGIC;
  signal W_62_11_i_15_n_0 : STD_LOGIC;
  signal W_62_11_i_16_n_0 : STD_LOGIC;
  signal W_62_11_i_17_n_0 : STD_LOGIC;
  signal W_62_11_i_2_n_0 : STD_LOGIC;
  signal W_62_11_i_3_n_0 : STD_LOGIC;
  signal W_62_11_i_4_n_0 : STD_LOGIC;
  signal W_62_11_i_5_n_0 : STD_LOGIC;
  signal W_62_11_i_6_n_0 : STD_LOGIC;
  signal W_62_11_i_7_n_0 : STD_LOGIC;
  signal W_62_11_i_8_n_0 : STD_LOGIC;
  signal W_62_11_i_9_n_0 : STD_LOGIC;
  signal W_62_15_i_10_n_0 : STD_LOGIC;
  signal W_62_15_i_11_n_0 : STD_LOGIC;
  signal W_62_15_i_12_n_0 : STD_LOGIC;
  signal W_62_15_i_13_n_0 : STD_LOGIC;
  signal W_62_15_i_14_n_0 : STD_LOGIC;
  signal W_62_15_i_15_n_0 : STD_LOGIC;
  signal W_62_15_i_16_n_0 : STD_LOGIC;
  signal W_62_15_i_17_n_0 : STD_LOGIC;
  signal W_62_15_i_2_n_0 : STD_LOGIC;
  signal W_62_15_i_3_n_0 : STD_LOGIC;
  signal W_62_15_i_4_n_0 : STD_LOGIC;
  signal W_62_15_i_5_n_0 : STD_LOGIC;
  signal W_62_15_i_6_n_0 : STD_LOGIC;
  signal W_62_15_i_7_n_0 : STD_LOGIC;
  signal W_62_15_i_8_n_0 : STD_LOGIC;
  signal W_62_15_i_9_n_0 : STD_LOGIC;
  signal W_62_19_i_10_n_0 : STD_LOGIC;
  signal W_62_19_i_11_n_0 : STD_LOGIC;
  signal W_62_19_i_12_n_0 : STD_LOGIC;
  signal W_62_19_i_13_n_0 : STD_LOGIC;
  signal W_62_19_i_14_n_0 : STD_LOGIC;
  signal W_62_19_i_15_n_0 : STD_LOGIC;
  signal W_62_19_i_16_n_0 : STD_LOGIC;
  signal W_62_19_i_17_n_0 : STD_LOGIC;
  signal W_62_19_i_2_n_0 : STD_LOGIC;
  signal W_62_19_i_3_n_0 : STD_LOGIC;
  signal W_62_19_i_4_n_0 : STD_LOGIC;
  signal W_62_19_i_5_n_0 : STD_LOGIC;
  signal W_62_19_i_6_n_0 : STD_LOGIC;
  signal W_62_19_i_7_n_0 : STD_LOGIC;
  signal W_62_19_i_8_n_0 : STD_LOGIC;
  signal W_62_19_i_9_n_0 : STD_LOGIC;
  signal W_62_23_i_10_n_0 : STD_LOGIC;
  signal W_62_23_i_11_n_0 : STD_LOGIC;
  signal W_62_23_i_12_n_0 : STD_LOGIC;
  signal W_62_23_i_13_n_0 : STD_LOGIC;
  signal W_62_23_i_14_n_0 : STD_LOGIC;
  signal W_62_23_i_15_n_0 : STD_LOGIC;
  signal W_62_23_i_16_n_0 : STD_LOGIC;
  signal W_62_23_i_17_n_0 : STD_LOGIC;
  signal W_62_23_i_2_n_0 : STD_LOGIC;
  signal W_62_23_i_3_n_0 : STD_LOGIC;
  signal W_62_23_i_4_n_0 : STD_LOGIC;
  signal W_62_23_i_5_n_0 : STD_LOGIC;
  signal W_62_23_i_6_n_0 : STD_LOGIC;
  signal W_62_23_i_7_n_0 : STD_LOGIC;
  signal W_62_23_i_8_n_0 : STD_LOGIC;
  signal W_62_23_i_9_n_0 : STD_LOGIC;
  signal W_62_27_i_10_n_0 : STD_LOGIC;
  signal W_62_27_i_11_n_0 : STD_LOGIC;
  signal W_62_27_i_12_n_0 : STD_LOGIC;
  signal W_62_27_i_13_n_0 : STD_LOGIC;
  signal W_62_27_i_14_n_0 : STD_LOGIC;
  signal W_62_27_i_15_n_0 : STD_LOGIC;
  signal W_62_27_i_16_n_0 : STD_LOGIC;
  signal W_62_27_i_17_n_0 : STD_LOGIC;
  signal W_62_27_i_2_n_0 : STD_LOGIC;
  signal W_62_27_i_3_n_0 : STD_LOGIC;
  signal W_62_27_i_4_n_0 : STD_LOGIC;
  signal W_62_27_i_5_n_0 : STD_LOGIC;
  signal W_62_27_i_6_n_0 : STD_LOGIC;
  signal W_62_27_i_7_n_0 : STD_LOGIC;
  signal W_62_27_i_8_n_0 : STD_LOGIC;
  signal W_62_27_i_9_n_0 : STD_LOGIC;
  signal W_62_31_i_10_n_0 : STD_LOGIC;
  signal W_62_31_i_11_n_0 : STD_LOGIC;
  signal W_62_31_i_12_n_0 : STD_LOGIC;
  signal W_62_31_i_13_n_0 : STD_LOGIC;
  signal W_62_31_i_14_n_0 : STD_LOGIC;
  signal W_62_31_i_15_n_0 : STD_LOGIC;
  signal W_62_31_i_17_n_0 : STD_LOGIC;
  signal W_62_31_i_19_n_0 : STD_LOGIC;
  signal W_62_31_i_2_n_0 : STD_LOGIC;
  signal W_62_31_i_3_n_0 : STD_LOGIC;
  signal W_62_31_i_4_n_0 : STD_LOGIC;
  signal W_62_31_i_5_n_0 : STD_LOGIC;
  signal W_62_31_i_6_n_0 : STD_LOGIC;
  signal W_62_31_i_7_n_0 : STD_LOGIC;
  signal W_62_31_i_8_n_0 : STD_LOGIC;
  signal W_62_31_i_9_n_0 : STD_LOGIC;
  signal W_62_3_i_10_n_0 : STD_LOGIC;
  signal W_62_3_i_11_n_0 : STD_LOGIC;
  signal W_62_3_i_15_n_0 : STD_LOGIC;
  signal W_62_3_i_2_n_0 : STD_LOGIC;
  signal W_62_3_i_3_n_0 : STD_LOGIC;
  signal W_62_3_i_4_n_0 : STD_LOGIC;
  signal W_62_3_i_5_n_0 : STD_LOGIC;
  signal W_62_3_i_6_n_0 : STD_LOGIC;
  signal W_62_3_i_7_n_0 : STD_LOGIC;
  signal W_62_3_i_8_n_0 : STD_LOGIC;
  signal W_62_3_i_9_n_0 : STD_LOGIC;
  signal W_62_7_i_10_n_0 : STD_LOGIC;
  signal W_62_7_i_11_n_0 : STD_LOGIC;
  signal W_62_7_i_12_n_0 : STD_LOGIC;
  signal W_62_7_i_13_n_0 : STD_LOGIC;
  signal W_62_7_i_14_n_0 : STD_LOGIC;
  signal W_62_7_i_15_n_0 : STD_LOGIC;
  signal W_62_7_i_16_n_0 : STD_LOGIC;
  signal W_62_7_i_17_n_0 : STD_LOGIC;
  signal W_62_7_i_2_n_0 : STD_LOGIC;
  signal W_62_7_i_3_n_0 : STD_LOGIC;
  signal W_62_7_i_4_n_0 : STD_LOGIC;
  signal W_62_7_i_5_n_0 : STD_LOGIC;
  signal W_62_7_i_6_n_0 : STD_LOGIC;
  signal W_62_7_i_7_n_0 : STD_LOGIC;
  signal W_62_7_i_8_n_0 : STD_LOGIC;
  signal W_62_7_i_9_n_0 : STD_LOGIC;
  signal W_63_11_i_10_n_0 : STD_LOGIC;
  signal W_63_11_i_11_n_0 : STD_LOGIC;
  signal W_63_11_i_12_n_0 : STD_LOGIC;
  signal W_63_11_i_13_n_0 : STD_LOGIC;
  signal W_63_11_i_14_n_0 : STD_LOGIC;
  signal W_63_11_i_15_n_0 : STD_LOGIC;
  signal W_63_11_i_16_n_0 : STD_LOGIC;
  signal W_63_11_i_17_n_0 : STD_LOGIC;
  signal W_63_11_i_2_n_0 : STD_LOGIC;
  signal W_63_11_i_3_n_0 : STD_LOGIC;
  signal W_63_11_i_4_n_0 : STD_LOGIC;
  signal W_63_11_i_5_n_0 : STD_LOGIC;
  signal W_63_11_i_6_n_0 : STD_LOGIC;
  signal W_63_11_i_7_n_0 : STD_LOGIC;
  signal W_63_11_i_8_n_0 : STD_LOGIC;
  signal W_63_11_i_9_n_0 : STD_LOGIC;
  signal W_63_15_i_10_n_0 : STD_LOGIC;
  signal W_63_15_i_11_n_0 : STD_LOGIC;
  signal W_63_15_i_12_n_0 : STD_LOGIC;
  signal W_63_15_i_13_n_0 : STD_LOGIC;
  signal W_63_15_i_14_n_0 : STD_LOGIC;
  signal W_63_15_i_15_n_0 : STD_LOGIC;
  signal W_63_15_i_16_n_0 : STD_LOGIC;
  signal W_63_15_i_17_n_0 : STD_LOGIC;
  signal W_63_15_i_2_n_0 : STD_LOGIC;
  signal W_63_15_i_3_n_0 : STD_LOGIC;
  signal W_63_15_i_4_n_0 : STD_LOGIC;
  signal W_63_15_i_5_n_0 : STD_LOGIC;
  signal W_63_15_i_6_n_0 : STD_LOGIC;
  signal W_63_15_i_7_n_0 : STD_LOGIC;
  signal W_63_15_i_8_n_0 : STD_LOGIC;
  signal W_63_15_i_9_n_0 : STD_LOGIC;
  signal W_63_19_i_10_n_0 : STD_LOGIC;
  signal W_63_19_i_11_n_0 : STD_LOGIC;
  signal W_63_19_i_12_n_0 : STD_LOGIC;
  signal W_63_19_i_13_n_0 : STD_LOGIC;
  signal W_63_19_i_14_n_0 : STD_LOGIC;
  signal W_63_19_i_15_n_0 : STD_LOGIC;
  signal W_63_19_i_16_n_0 : STD_LOGIC;
  signal W_63_19_i_17_n_0 : STD_LOGIC;
  signal W_63_19_i_2_n_0 : STD_LOGIC;
  signal W_63_19_i_3_n_0 : STD_LOGIC;
  signal W_63_19_i_4_n_0 : STD_LOGIC;
  signal W_63_19_i_5_n_0 : STD_LOGIC;
  signal W_63_19_i_6_n_0 : STD_LOGIC;
  signal W_63_19_i_7_n_0 : STD_LOGIC;
  signal W_63_19_i_8_n_0 : STD_LOGIC;
  signal W_63_19_i_9_n_0 : STD_LOGIC;
  signal W_63_23_i_10_n_0 : STD_LOGIC;
  signal W_63_23_i_11_n_0 : STD_LOGIC;
  signal W_63_23_i_12_n_0 : STD_LOGIC;
  signal W_63_23_i_13_n_0 : STD_LOGIC;
  signal W_63_23_i_14_n_0 : STD_LOGIC;
  signal W_63_23_i_15_n_0 : STD_LOGIC;
  signal W_63_23_i_16_n_0 : STD_LOGIC;
  signal W_63_23_i_17_n_0 : STD_LOGIC;
  signal W_63_23_i_2_n_0 : STD_LOGIC;
  signal W_63_23_i_3_n_0 : STD_LOGIC;
  signal W_63_23_i_4_n_0 : STD_LOGIC;
  signal W_63_23_i_5_n_0 : STD_LOGIC;
  signal W_63_23_i_6_n_0 : STD_LOGIC;
  signal W_63_23_i_7_n_0 : STD_LOGIC;
  signal W_63_23_i_8_n_0 : STD_LOGIC;
  signal W_63_23_i_9_n_0 : STD_LOGIC;
  signal W_63_27_i_10_n_0 : STD_LOGIC;
  signal W_63_27_i_11_n_0 : STD_LOGIC;
  signal W_63_27_i_12_n_0 : STD_LOGIC;
  signal W_63_27_i_13_n_0 : STD_LOGIC;
  signal W_63_27_i_14_n_0 : STD_LOGIC;
  signal W_63_27_i_15_n_0 : STD_LOGIC;
  signal W_63_27_i_16_n_0 : STD_LOGIC;
  signal W_63_27_i_17_n_0 : STD_LOGIC;
  signal W_63_27_i_2_n_0 : STD_LOGIC;
  signal W_63_27_i_3_n_0 : STD_LOGIC;
  signal W_63_27_i_4_n_0 : STD_LOGIC;
  signal W_63_27_i_5_n_0 : STD_LOGIC;
  signal W_63_27_i_6_n_0 : STD_LOGIC;
  signal W_63_27_i_7_n_0 : STD_LOGIC;
  signal W_63_27_i_8_n_0 : STD_LOGIC;
  signal W_63_27_i_9_n_0 : STD_LOGIC;
  signal W_63_31_i_10_n_0 : STD_LOGIC;
  signal W_63_31_i_11_n_0 : STD_LOGIC;
  signal W_63_31_i_12_n_0 : STD_LOGIC;
  signal W_63_31_i_13_n_0 : STD_LOGIC;
  signal W_63_31_i_14_n_0 : STD_LOGIC;
  signal W_63_31_i_15_n_0 : STD_LOGIC;
  signal W_63_31_i_17_n_0 : STD_LOGIC;
  signal W_63_31_i_19_n_0 : STD_LOGIC;
  signal W_63_31_i_2_n_0 : STD_LOGIC;
  signal W_63_31_i_3_n_0 : STD_LOGIC;
  signal W_63_31_i_4_n_0 : STD_LOGIC;
  signal W_63_31_i_5_n_0 : STD_LOGIC;
  signal W_63_31_i_6_n_0 : STD_LOGIC;
  signal W_63_31_i_7_n_0 : STD_LOGIC;
  signal W_63_31_i_8_n_0 : STD_LOGIC;
  signal W_63_31_i_9_n_0 : STD_LOGIC;
  signal W_63_3_i_10_n_0 : STD_LOGIC;
  signal W_63_3_i_11_n_0 : STD_LOGIC;
  signal W_63_3_i_15_n_0 : STD_LOGIC;
  signal W_63_3_i_2_n_0 : STD_LOGIC;
  signal W_63_3_i_3_n_0 : STD_LOGIC;
  signal W_63_3_i_4_n_0 : STD_LOGIC;
  signal W_63_3_i_5_n_0 : STD_LOGIC;
  signal W_63_3_i_6_n_0 : STD_LOGIC;
  signal W_63_3_i_7_n_0 : STD_LOGIC;
  signal W_63_3_i_8_n_0 : STD_LOGIC;
  signal W_63_3_i_9_n_0 : STD_LOGIC;
  signal W_63_7_i_10_n_0 : STD_LOGIC;
  signal W_63_7_i_11_n_0 : STD_LOGIC;
  signal W_63_7_i_12_n_0 : STD_LOGIC;
  signal W_63_7_i_13_n_0 : STD_LOGIC;
  signal W_63_7_i_14_n_0 : STD_LOGIC;
  signal W_63_7_i_15_n_0 : STD_LOGIC;
  signal W_63_7_i_16_n_0 : STD_LOGIC;
  signal W_63_7_i_17_n_0 : STD_LOGIC;
  signal W_63_7_i_2_n_0 : STD_LOGIC;
  signal W_63_7_i_3_n_0 : STD_LOGIC;
  signal W_63_7_i_4_n_0 : STD_LOGIC;
  signal W_63_7_i_5_n_0 : STD_LOGIC;
  signal W_63_7_i_6_n_0 : STD_LOGIC;
  signal W_63_7_i_7_n_0 : STD_LOGIC;
  signal W_63_7_i_8_n_0 : STD_LOGIC;
  signal W_63_7_i_9_n_0 : STD_LOGIC;
  signal W_INT_62_31 : STD_LOGIC;
  signal W_INT_62_30 : STD_LOGIC;
  signal W_INT_62_29 : STD_LOGIC;
  signal W_INT_62_28 : STD_LOGIC;
  signal W_INT_62_27 : STD_LOGIC;
  signal W_INT_62_26 : STD_LOGIC;
  signal W_INT_62_25 : STD_LOGIC;
  signal W_INT_62_24 : STD_LOGIC;
  signal W_INT_62_23 : STD_LOGIC;
  signal W_INT_62_22 : STD_LOGIC;
  signal W_INT_62_21 : STD_LOGIC;
  signal W_INT_62_20 : STD_LOGIC;
  signal W_INT_62_19 : STD_LOGIC;
  signal W_INT_62_18 : STD_LOGIC;
  signal W_INT_62_17 : STD_LOGIC;
  signal W_INT_62_16 : STD_LOGIC;
  signal W_INT_62_15 : STD_LOGIC;
  signal W_INT_62_14 : STD_LOGIC;
  signal W_INT_62_13 : STD_LOGIC;
  signal W_INT_62_12 : STD_LOGIC;
  signal W_INT_62_11 : STD_LOGIC;
  signal W_INT_62_10 : STD_LOGIC;
  signal W_INT_62_9 : STD_LOGIC;
  signal W_INT_62_8 : STD_LOGIC;
  signal W_INT_62_7 : STD_LOGIC;
  signal W_INT_62_6 : STD_LOGIC;
  signal W_INT_62_5 : STD_LOGIC;
  signal W_INT_62_4 : STD_LOGIC;
  signal W_INT_62_3 : STD_LOGIC;
  signal W_INT_62_2 : STD_LOGIC;
  signal W_INT_62_1 : STD_LOGIC;
  signal W_INT_62_0 : STD_LOGIC;
  signal W_INT_63_31 : STD_LOGIC;
  signal W_INT_63_30 : STD_LOGIC;
  signal W_INT_63_29 : STD_LOGIC;
  signal W_INT_63_28 : STD_LOGIC;
  signal W_INT_63_27 : STD_LOGIC;
  signal W_INT_63_26 : STD_LOGIC;
  signal W_INT_63_25 : STD_LOGIC;
  signal W_INT_63_24 : STD_LOGIC;
  signal W_INT_63_23 : STD_LOGIC;
  signal W_INT_63_22 : STD_LOGIC;
  signal W_INT_63_21 : STD_LOGIC;
  signal W_INT_63_20 : STD_LOGIC;
  signal W_INT_63_19 : STD_LOGIC;
  signal W_INT_63_18 : STD_LOGIC;
  signal W_INT_63_17 : STD_LOGIC;
  signal W_INT_63_16 : STD_LOGIC;
  signal W_INT_63_15 : STD_LOGIC;
  signal W_INT_63_14 : STD_LOGIC;
  signal W_INT_63_13 : STD_LOGIC;
  signal W_INT_63_12 : STD_LOGIC;
  signal W_INT_63_11 : STD_LOGIC;
  signal W_INT_63_10 : STD_LOGIC;
  signal W_INT_63_9 : STD_LOGIC;
  signal W_INT_63_8 : STD_LOGIC;
  signal W_INT_63_7 : STD_LOGIC;
  signal W_INT_63_6 : STD_LOGIC;
  signal W_INT_63_5 : STD_LOGIC;
  signal W_INT_63_4 : STD_LOGIC;
  signal W_INT_63_3 : STD_LOGIC;
  signal W_INT_63_2 : STD_LOGIC;
  signal W_INT_63_1 : STD_LOGIC;
  signal W_INT_63_0 : STD_LOGIC;
  signal W_reg_0_31 : STD_LOGIC;
  signal W_reg_0_30 : STD_LOGIC;
  signal W_reg_0_29 : STD_LOGIC;
  signal W_reg_0_28 : STD_LOGIC;
  signal W_reg_0_27 : STD_LOGIC;
  signal W_reg_0_26 : STD_LOGIC;
  signal W_reg_0_25 : STD_LOGIC;
  signal W_reg_0_24 : STD_LOGIC;
  signal W_reg_0_23 : STD_LOGIC;
  signal W_reg_0_22 : STD_LOGIC;
  signal W_reg_0_21 : STD_LOGIC;
  signal W_reg_0_20 : STD_LOGIC;
  signal W_reg_0_19 : STD_LOGIC;
  signal W_reg_0_18 : STD_LOGIC;
  signal W_reg_0_17 : STD_LOGIC;
  signal W_reg_0_16 : STD_LOGIC;
  signal W_reg_0_15 : STD_LOGIC;
  signal W_reg_0_14 : STD_LOGIC;
  signal W_reg_0_13 : STD_LOGIC;
  signal W_reg_0_12 : STD_LOGIC;
  signal W_reg_0_11 : STD_LOGIC;
  signal W_reg_0_10 : STD_LOGIC;
  signal W_reg_0_9 : STD_LOGIC;
  signal W_reg_0_8 : STD_LOGIC;
  signal W_reg_0_7 : STD_LOGIC;
  signal W_reg_0_6 : STD_LOGIC;
  signal W_reg_0_5 : STD_LOGIC;
  signal W_reg_0_4 : STD_LOGIC;
  signal W_reg_0_3 : STD_LOGIC;
  signal W_reg_0_2 : STD_LOGIC;
  signal W_reg_0_1 : STD_LOGIC;
  signal W_reg_0_0 : STD_LOGIC;
  signal W_reg_10_31 : STD_LOGIC;
  signal W_reg_10_30 : STD_LOGIC;
  signal W_reg_10_29 : STD_LOGIC;
  signal W_reg_10_28 : STD_LOGIC;
  signal W_reg_10_27 : STD_LOGIC;
  signal W_reg_10_26 : STD_LOGIC;
  signal W_reg_10_25 : STD_LOGIC;
  signal W_reg_10_24 : STD_LOGIC;
  signal W_reg_10_23 : STD_LOGIC;
  signal W_reg_10_22 : STD_LOGIC;
  signal W_reg_10_21 : STD_LOGIC;
  signal W_reg_10_20 : STD_LOGIC;
  signal W_reg_10_19 : STD_LOGIC;
  signal W_reg_10_18 : STD_LOGIC;
  signal W_reg_10_17 : STD_LOGIC;
  signal W_reg_10_16 : STD_LOGIC;
  signal W_reg_10_15 : STD_LOGIC;
  signal W_reg_10_14 : STD_LOGIC;
  signal W_reg_10_13 : STD_LOGIC;
  signal W_reg_10_12 : STD_LOGIC;
  signal W_reg_10_11 : STD_LOGIC;
  signal W_reg_10_10 : STD_LOGIC;
  signal W_reg_10_9 : STD_LOGIC;
  signal W_reg_10_8 : STD_LOGIC;
  signal W_reg_10_7 : STD_LOGIC;
  signal W_reg_10_6 : STD_LOGIC;
  signal W_reg_10_5 : STD_LOGIC;
  signal W_reg_10_4 : STD_LOGIC;
  signal W_reg_10_3 : STD_LOGIC;
  signal W_reg_10_2 : STD_LOGIC;
  signal W_reg_10_1 : STD_LOGIC;
  signal W_reg_10_0 : STD_LOGIC;
  signal W_reg_11_31 : STD_LOGIC;
  signal W_reg_11_30 : STD_LOGIC;
  signal W_reg_11_29 : STD_LOGIC;
  signal W_reg_11_28 : STD_LOGIC;
  signal W_reg_11_27 : STD_LOGIC;
  signal W_reg_11_26 : STD_LOGIC;
  signal W_reg_11_25 : STD_LOGIC;
  signal W_reg_11_24 : STD_LOGIC;
  signal W_reg_11_23 : STD_LOGIC;
  signal W_reg_11_22 : STD_LOGIC;
  signal W_reg_11_21 : STD_LOGIC;
  signal W_reg_11_20 : STD_LOGIC;
  signal W_reg_11_19 : STD_LOGIC;
  signal W_reg_11_18 : STD_LOGIC;
  signal W_reg_11_17 : STD_LOGIC;
  signal W_reg_11_16 : STD_LOGIC;
  signal W_reg_11_15 : STD_LOGIC;
  signal W_reg_11_14 : STD_LOGIC;
  signal W_reg_11_13 : STD_LOGIC;
  signal W_reg_11_12 : STD_LOGIC;
  signal W_reg_11_11 : STD_LOGIC;
  signal W_reg_11_10 : STD_LOGIC;
  signal W_reg_11_9 : STD_LOGIC;
  signal W_reg_11_8 : STD_LOGIC;
  signal W_reg_11_7 : STD_LOGIC;
  signal W_reg_11_6 : STD_LOGIC;
  signal W_reg_11_5 : STD_LOGIC;
  signal W_reg_11_4 : STD_LOGIC;
  signal W_reg_11_3 : STD_LOGIC;
  signal W_reg_11_2 : STD_LOGIC;
  signal W_reg_11_1 : STD_LOGIC;
  signal W_reg_11_0 : STD_LOGIC;
  signal W_reg_12_31 : STD_LOGIC;
  signal W_reg_12_30 : STD_LOGIC;
  signal W_reg_12_29 : STD_LOGIC;
  signal W_reg_12_28 : STD_LOGIC;
  signal W_reg_12_27 : STD_LOGIC;
  signal W_reg_12_26 : STD_LOGIC;
  signal W_reg_12_25 : STD_LOGIC;
  signal W_reg_12_24 : STD_LOGIC;
  signal W_reg_12_23 : STD_LOGIC;
  signal W_reg_12_22 : STD_LOGIC;
  signal W_reg_12_21 : STD_LOGIC;
  signal W_reg_12_20 : STD_LOGIC;
  signal W_reg_12_19 : STD_LOGIC;
  signal W_reg_12_18 : STD_LOGIC;
  signal W_reg_12_17 : STD_LOGIC;
  signal W_reg_12_16 : STD_LOGIC;
  signal W_reg_12_15 : STD_LOGIC;
  signal W_reg_12_14 : STD_LOGIC;
  signal W_reg_12_13 : STD_LOGIC;
  signal W_reg_12_12 : STD_LOGIC;
  signal W_reg_12_11 : STD_LOGIC;
  signal W_reg_12_10 : STD_LOGIC;
  signal W_reg_12_9 : STD_LOGIC;
  signal W_reg_12_8 : STD_LOGIC;
  signal W_reg_12_7 : STD_LOGIC;
  signal W_reg_12_6 : STD_LOGIC;
  signal W_reg_12_5 : STD_LOGIC;
  signal W_reg_12_4 : STD_LOGIC;
  signal W_reg_12_3 : STD_LOGIC;
  signal W_reg_12_2 : STD_LOGIC;
  signal W_reg_12_1 : STD_LOGIC;
  signal W_reg_12_0 : STD_LOGIC;
  signal W_reg_13_31 : STD_LOGIC;
  signal W_reg_13_30 : STD_LOGIC;
  signal W_reg_13_29 : STD_LOGIC;
  signal W_reg_13_28 : STD_LOGIC;
  signal W_reg_13_27 : STD_LOGIC;
  signal W_reg_13_26 : STD_LOGIC;
  signal W_reg_13_25 : STD_LOGIC;
  signal W_reg_13_24 : STD_LOGIC;
  signal W_reg_13_23 : STD_LOGIC;
  signal W_reg_13_22 : STD_LOGIC;
  signal W_reg_13_21 : STD_LOGIC;
  signal W_reg_13_20 : STD_LOGIC;
  signal W_reg_13_19 : STD_LOGIC;
  signal W_reg_13_18 : STD_LOGIC;
  signal W_reg_13_17 : STD_LOGIC;
  signal W_reg_13_16 : STD_LOGIC;
  signal W_reg_13_15 : STD_LOGIC;
  signal W_reg_13_14 : STD_LOGIC;
  signal W_reg_13_13 : STD_LOGIC;
  signal W_reg_13_12 : STD_LOGIC;
  signal W_reg_13_11 : STD_LOGIC;
  signal W_reg_13_10 : STD_LOGIC;
  signal W_reg_13_9 : STD_LOGIC;
  signal W_reg_13_8 : STD_LOGIC;
  signal W_reg_13_7 : STD_LOGIC;
  signal W_reg_13_6 : STD_LOGIC;
  signal W_reg_13_5 : STD_LOGIC;
  signal W_reg_13_4 : STD_LOGIC;
  signal W_reg_13_3 : STD_LOGIC;
  signal W_reg_13_2 : STD_LOGIC;
  signal W_reg_13_1 : STD_LOGIC;
  signal W_reg_13_0 : STD_LOGIC;
  signal W_reg_14_31 : STD_LOGIC;
  signal W_reg_14_30 : STD_LOGIC;
  signal W_reg_14_29 : STD_LOGIC;
  signal W_reg_14_28 : STD_LOGIC;
  signal W_reg_14_27 : STD_LOGIC;
  signal W_reg_14_26 : STD_LOGIC;
  signal W_reg_14_25 : STD_LOGIC;
  signal W_reg_14_24 : STD_LOGIC;
  signal W_reg_14_23 : STD_LOGIC;
  signal W_reg_14_22 : STD_LOGIC;
  signal W_reg_14_21 : STD_LOGIC;
  signal W_reg_14_20 : STD_LOGIC;
  signal W_reg_14_19 : STD_LOGIC;
  signal W_reg_14_18 : STD_LOGIC;
  signal W_reg_14_17 : STD_LOGIC;
  signal W_reg_14_16 : STD_LOGIC;
  signal W_reg_14_15 : STD_LOGIC;
  signal W_reg_14_14 : STD_LOGIC;
  signal W_reg_14_13 : STD_LOGIC;
  signal W_reg_14_12 : STD_LOGIC;
  signal W_reg_14_11 : STD_LOGIC;
  signal W_reg_14_10 : STD_LOGIC;
  signal W_reg_14_9 : STD_LOGIC;
  signal W_reg_14_8 : STD_LOGIC;
  signal W_reg_14_7 : STD_LOGIC;
  signal W_reg_14_6 : STD_LOGIC;
  signal W_reg_14_5 : STD_LOGIC;
  signal W_reg_14_4 : STD_LOGIC;
  signal W_reg_14_3 : STD_LOGIC;
  signal W_reg_14_2 : STD_LOGIC;
  signal W_reg_14_1 : STD_LOGIC;
  signal W_reg_14_0 : STD_LOGIC;
  signal W_reg_15_31 : STD_LOGIC;
  signal W_reg_15_30 : STD_LOGIC;
  signal W_reg_15_29 : STD_LOGIC;
  signal W_reg_15_28 : STD_LOGIC;
  signal W_reg_15_27 : STD_LOGIC;
  signal W_reg_15_26 : STD_LOGIC;
  signal W_reg_15_25 : STD_LOGIC;
  signal W_reg_15_24 : STD_LOGIC;
  signal W_reg_15_23 : STD_LOGIC;
  signal W_reg_15_22 : STD_LOGIC;
  signal W_reg_15_21 : STD_LOGIC;
  signal W_reg_15_20 : STD_LOGIC;
  signal W_reg_15_19 : STD_LOGIC;
  signal W_reg_15_18 : STD_LOGIC;
  signal W_reg_15_17 : STD_LOGIC;
  signal W_reg_15_16 : STD_LOGIC;
  signal W_reg_15_15 : STD_LOGIC;
  signal W_reg_15_14 : STD_LOGIC;
  signal W_reg_15_13 : STD_LOGIC;
  signal W_reg_15_12 : STD_LOGIC;
  signal W_reg_15_11 : STD_LOGIC;
  signal W_reg_15_10 : STD_LOGIC;
  signal W_reg_15_9 : STD_LOGIC;
  signal W_reg_15_8 : STD_LOGIC;
  signal W_reg_15_7 : STD_LOGIC;
  signal W_reg_15_6 : STD_LOGIC;
  signal W_reg_15_5 : STD_LOGIC;
  signal W_reg_15_4 : STD_LOGIC;
  signal W_reg_15_3 : STD_LOGIC;
  signal W_reg_15_2 : STD_LOGIC;
  signal W_reg_15_1 : STD_LOGIC;
  signal W_reg_15_0 : STD_LOGIC;
  signal W_reg_16_31 : STD_LOGIC;
  signal W_reg_16_30 : STD_LOGIC;
  signal W_reg_16_29 : STD_LOGIC;
  signal W_reg_16_28 : STD_LOGIC;
  signal W_reg_16_27 : STD_LOGIC;
  signal W_reg_16_26 : STD_LOGIC;
  signal W_reg_16_25 : STD_LOGIC;
  signal W_reg_16_24 : STD_LOGIC;
  signal W_reg_16_23 : STD_LOGIC;
  signal W_reg_16_22 : STD_LOGIC;
  signal W_reg_16_21 : STD_LOGIC;
  signal W_reg_16_20 : STD_LOGIC;
  signal W_reg_16_19 : STD_LOGIC;
  signal W_reg_16_18 : STD_LOGIC;
  signal W_reg_16_17 : STD_LOGIC;
  signal W_reg_16_16 : STD_LOGIC;
  signal W_reg_16_15 : STD_LOGIC;
  signal W_reg_16_14 : STD_LOGIC;
  signal W_reg_16_13 : STD_LOGIC;
  signal W_reg_16_12 : STD_LOGIC;
  signal W_reg_16_11 : STD_LOGIC;
  signal W_reg_16_10 : STD_LOGIC;
  signal W_reg_16_9 : STD_LOGIC;
  signal W_reg_16_8 : STD_LOGIC;
  signal W_reg_16_7 : STD_LOGIC;
  signal W_reg_16_6 : STD_LOGIC;
  signal W_reg_16_5 : STD_LOGIC;
  signal W_reg_16_4 : STD_LOGIC;
  signal W_reg_16_3 : STD_LOGIC;
  signal W_reg_16_2 : STD_LOGIC;
  signal W_reg_16_1 : STD_LOGIC;
  signal W_reg_16_0 : STD_LOGIC;
  signal W_reg_16_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_16_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_16_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_16_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_16_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_16_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_16_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_16_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_16_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_16_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_16_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_16_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_16_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_16_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_16_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_16_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_16_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_16_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_16_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_16_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_16_31_i_2_n_1 : STD_LOGIC;
  signal W_reg_16_31_i_2_n_2 : STD_LOGIC;
  signal W_reg_16_31_i_2_n_3 : STD_LOGIC;
  signal W_reg_16_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_16_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_16_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_16_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_16_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_16_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_16_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_16_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_17_31 : STD_LOGIC;
  signal W_reg_17_30 : STD_LOGIC;
  signal W_reg_17_29 : STD_LOGIC;
  signal W_reg_17_28 : STD_LOGIC;
  signal W_reg_17_27 : STD_LOGIC;
  signal W_reg_17_26 : STD_LOGIC;
  signal W_reg_17_25 : STD_LOGIC;
  signal W_reg_17_24 : STD_LOGIC;
  signal W_reg_17_23 : STD_LOGIC;
  signal W_reg_17_22 : STD_LOGIC;
  signal W_reg_17_21 : STD_LOGIC;
  signal W_reg_17_20 : STD_LOGIC;
  signal W_reg_17_19 : STD_LOGIC;
  signal W_reg_17_18 : STD_LOGIC;
  signal W_reg_17_17 : STD_LOGIC;
  signal W_reg_17_16 : STD_LOGIC;
  signal W_reg_17_15 : STD_LOGIC;
  signal W_reg_17_14 : STD_LOGIC;
  signal W_reg_17_13 : STD_LOGIC;
  signal W_reg_17_12 : STD_LOGIC;
  signal W_reg_17_11 : STD_LOGIC;
  signal W_reg_17_10 : STD_LOGIC;
  signal W_reg_17_9 : STD_LOGIC;
  signal W_reg_17_8 : STD_LOGIC;
  signal W_reg_17_7 : STD_LOGIC;
  signal W_reg_17_6 : STD_LOGIC;
  signal W_reg_17_5 : STD_LOGIC;
  signal W_reg_17_4 : STD_LOGIC;
  signal W_reg_17_3 : STD_LOGIC;
  signal W_reg_17_2 : STD_LOGIC;
  signal W_reg_17_1 : STD_LOGIC;
  signal W_reg_17_0 : STD_LOGIC;
  signal W_reg_17_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_17_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_17_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_17_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_17_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_17_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_17_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_17_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_17_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_17_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_17_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_17_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_17_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_17_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_17_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_17_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_17_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_17_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_17_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_17_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_17_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_17_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_17_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_17_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_17_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_17_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_17_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_17_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_17_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_17_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_17_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_18_31 : STD_LOGIC;
  signal W_reg_18_30 : STD_LOGIC;
  signal W_reg_18_29 : STD_LOGIC;
  signal W_reg_18_28 : STD_LOGIC;
  signal W_reg_18_27 : STD_LOGIC;
  signal W_reg_18_26 : STD_LOGIC;
  signal W_reg_18_25 : STD_LOGIC;
  signal W_reg_18_24 : STD_LOGIC;
  signal W_reg_18_23 : STD_LOGIC;
  signal W_reg_18_22 : STD_LOGIC;
  signal W_reg_18_21 : STD_LOGIC;
  signal W_reg_18_20 : STD_LOGIC;
  signal W_reg_18_19 : STD_LOGIC;
  signal W_reg_18_18 : STD_LOGIC;
  signal W_reg_18_17 : STD_LOGIC;
  signal W_reg_18_16 : STD_LOGIC;
  signal W_reg_18_15 : STD_LOGIC;
  signal W_reg_18_14 : STD_LOGIC;
  signal W_reg_18_13 : STD_LOGIC;
  signal W_reg_18_12 : STD_LOGIC;
  signal W_reg_18_11 : STD_LOGIC;
  signal W_reg_18_10 : STD_LOGIC;
  signal W_reg_18_9 : STD_LOGIC;
  signal W_reg_18_8 : STD_LOGIC;
  signal W_reg_18_7 : STD_LOGIC;
  signal W_reg_18_6 : STD_LOGIC;
  signal W_reg_18_5 : STD_LOGIC;
  signal W_reg_18_4 : STD_LOGIC;
  signal W_reg_18_3 : STD_LOGIC;
  signal W_reg_18_2 : STD_LOGIC;
  signal W_reg_18_1 : STD_LOGIC;
  signal W_reg_18_0 : STD_LOGIC;
  signal W_reg_18_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_18_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_18_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_18_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_18_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_18_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_18_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_18_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_18_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_18_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_18_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_18_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_18_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_18_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_18_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_18_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_18_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_18_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_18_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_18_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_18_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_18_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_18_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_18_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_18_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_18_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_18_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_18_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_18_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_18_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_18_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_19_31 : STD_LOGIC;
  signal W_reg_19_30 : STD_LOGIC;
  signal W_reg_19_29 : STD_LOGIC;
  signal W_reg_19_28 : STD_LOGIC;
  signal W_reg_19_27 : STD_LOGIC;
  signal W_reg_19_26 : STD_LOGIC;
  signal W_reg_19_25 : STD_LOGIC;
  signal W_reg_19_24 : STD_LOGIC;
  signal W_reg_19_23 : STD_LOGIC;
  signal W_reg_19_22 : STD_LOGIC;
  signal W_reg_19_21 : STD_LOGIC;
  signal W_reg_19_20 : STD_LOGIC;
  signal W_reg_19_19 : STD_LOGIC;
  signal W_reg_19_18 : STD_LOGIC;
  signal W_reg_19_17 : STD_LOGIC;
  signal W_reg_19_16 : STD_LOGIC;
  signal W_reg_19_15 : STD_LOGIC;
  signal W_reg_19_14 : STD_LOGIC;
  signal W_reg_19_13 : STD_LOGIC;
  signal W_reg_19_12 : STD_LOGIC;
  signal W_reg_19_11 : STD_LOGIC;
  signal W_reg_19_10 : STD_LOGIC;
  signal W_reg_19_9 : STD_LOGIC;
  signal W_reg_19_8 : STD_LOGIC;
  signal W_reg_19_7 : STD_LOGIC;
  signal W_reg_19_6 : STD_LOGIC;
  signal W_reg_19_5 : STD_LOGIC;
  signal W_reg_19_4 : STD_LOGIC;
  signal W_reg_19_3 : STD_LOGIC;
  signal W_reg_19_2 : STD_LOGIC;
  signal W_reg_19_1 : STD_LOGIC;
  signal W_reg_19_0 : STD_LOGIC;
  signal W_reg_19_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_19_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_19_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_19_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_19_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_19_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_19_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_19_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_19_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_19_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_19_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_19_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_19_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_19_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_19_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_19_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_19_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_19_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_19_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_19_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_19_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_19_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_19_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_19_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_19_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_19_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_19_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_19_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_19_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_19_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_19_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_1_31 : STD_LOGIC;
  signal W_reg_1_30 : STD_LOGIC;
  signal W_reg_1_29 : STD_LOGIC;
  signal W_reg_1_28 : STD_LOGIC;
  signal W_reg_1_27 : STD_LOGIC;
  signal W_reg_1_26 : STD_LOGIC;
  signal W_reg_1_25 : STD_LOGIC;
  signal W_reg_1_24 : STD_LOGIC;
  signal W_reg_1_23 : STD_LOGIC;
  signal W_reg_1_22 : STD_LOGIC;
  signal W_reg_1_21 : STD_LOGIC;
  signal W_reg_1_20 : STD_LOGIC;
  signal W_reg_1_19 : STD_LOGIC;
  signal W_reg_1_18 : STD_LOGIC;
  signal W_reg_1_17 : STD_LOGIC;
  signal W_reg_1_16 : STD_LOGIC;
  signal W_reg_1_15 : STD_LOGIC;
  signal W_reg_1_14 : STD_LOGIC;
  signal W_reg_1_13 : STD_LOGIC;
  signal W_reg_1_12 : STD_LOGIC;
  signal W_reg_1_11 : STD_LOGIC;
  signal W_reg_1_10 : STD_LOGIC;
  signal W_reg_1_9 : STD_LOGIC;
  signal W_reg_1_8 : STD_LOGIC;
  signal W_reg_1_7 : STD_LOGIC;
  signal W_reg_1_6 : STD_LOGIC;
  signal W_reg_1_5 : STD_LOGIC;
  signal W_reg_1_4 : STD_LOGIC;
  signal W_reg_1_3 : STD_LOGIC;
  signal W_reg_1_2 : STD_LOGIC;
  signal W_reg_1_1 : STD_LOGIC;
  signal W_reg_1_0 : STD_LOGIC;
  signal W_reg_20_31 : STD_LOGIC;
  signal W_reg_20_30 : STD_LOGIC;
  signal W_reg_20_29 : STD_LOGIC;
  signal W_reg_20_28 : STD_LOGIC;
  signal W_reg_20_27 : STD_LOGIC;
  signal W_reg_20_26 : STD_LOGIC;
  signal W_reg_20_25 : STD_LOGIC;
  signal W_reg_20_24 : STD_LOGIC;
  signal W_reg_20_23 : STD_LOGIC;
  signal W_reg_20_22 : STD_LOGIC;
  signal W_reg_20_21 : STD_LOGIC;
  signal W_reg_20_20 : STD_LOGIC;
  signal W_reg_20_19 : STD_LOGIC;
  signal W_reg_20_18 : STD_LOGIC;
  signal W_reg_20_17 : STD_LOGIC;
  signal W_reg_20_16 : STD_LOGIC;
  signal W_reg_20_15 : STD_LOGIC;
  signal W_reg_20_14 : STD_LOGIC;
  signal W_reg_20_13 : STD_LOGIC;
  signal W_reg_20_12 : STD_LOGIC;
  signal W_reg_20_11 : STD_LOGIC;
  signal W_reg_20_10 : STD_LOGIC;
  signal W_reg_20_9 : STD_LOGIC;
  signal W_reg_20_8 : STD_LOGIC;
  signal W_reg_20_7 : STD_LOGIC;
  signal W_reg_20_6 : STD_LOGIC;
  signal W_reg_20_5 : STD_LOGIC;
  signal W_reg_20_4 : STD_LOGIC;
  signal W_reg_20_3 : STD_LOGIC;
  signal W_reg_20_2 : STD_LOGIC;
  signal W_reg_20_1 : STD_LOGIC;
  signal W_reg_20_0 : STD_LOGIC;
  signal W_reg_20_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_20_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_20_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_20_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_20_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_20_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_20_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_20_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_20_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_20_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_20_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_20_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_20_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_20_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_20_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_20_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_20_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_20_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_20_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_20_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_20_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_20_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_20_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_20_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_20_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_20_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_20_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_20_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_20_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_20_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_20_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_21_31 : STD_LOGIC;
  signal W_reg_21_30 : STD_LOGIC;
  signal W_reg_21_29 : STD_LOGIC;
  signal W_reg_21_28 : STD_LOGIC;
  signal W_reg_21_27 : STD_LOGIC;
  signal W_reg_21_26 : STD_LOGIC;
  signal W_reg_21_25 : STD_LOGIC;
  signal W_reg_21_24 : STD_LOGIC;
  signal W_reg_21_23 : STD_LOGIC;
  signal W_reg_21_22 : STD_LOGIC;
  signal W_reg_21_21 : STD_LOGIC;
  signal W_reg_21_20 : STD_LOGIC;
  signal W_reg_21_19 : STD_LOGIC;
  signal W_reg_21_18 : STD_LOGIC;
  signal W_reg_21_17 : STD_LOGIC;
  signal W_reg_21_16 : STD_LOGIC;
  signal W_reg_21_15 : STD_LOGIC;
  signal W_reg_21_14 : STD_LOGIC;
  signal W_reg_21_13 : STD_LOGIC;
  signal W_reg_21_12 : STD_LOGIC;
  signal W_reg_21_11 : STD_LOGIC;
  signal W_reg_21_10 : STD_LOGIC;
  signal W_reg_21_9 : STD_LOGIC;
  signal W_reg_21_8 : STD_LOGIC;
  signal W_reg_21_7 : STD_LOGIC;
  signal W_reg_21_6 : STD_LOGIC;
  signal W_reg_21_5 : STD_LOGIC;
  signal W_reg_21_4 : STD_LOGIC;
  signal W_reg_21_3 : STD_LOGIC;
  signal W_reg_21_2 : STD_LOGIC;
  signal W_reg_21_1 : STD_LOGIC;
  signal W_reg_21_0 : STD_LOGIC;
  signal W_reg_21_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_21_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_21_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_21_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_21_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_21_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_21_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_21_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_21_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_21_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_21_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_21_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_21_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_21_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_21_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_21_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_21_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_21_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_21_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_21_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_21_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_21_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_21_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_21_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_21_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_21_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_21_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_21_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_21_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_21_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_21_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_22_31 : STD_LOGIC;
  signal W_reg_22_30 : STD_LOGIC;
  signal W_reg_22_29 : STD_LOGIC;
  signal W_reg_22_28 : STD_LOGIC;
  signal W_reg_22_27 : STD_LOGIC;
  signal W_reg_22_26 : STD_LOGIC;
  signal W_reg_22_25 : STD_LOGIC;
  signal W_reg_22_24 : STD_LOGIC;
  signal W_reg_22_23 : STD_LOGIC;
  signal W_reg_22_22 : STD_LOGIC;
  signal W_reg_22_21 : STD_LOGIC;
  signal W_reg_22_20 : STD_LOGIC;
  signal W_reg_22_19 : STD_LOGIC;
  signal W_reg_22_18 : STD_LOGIC;
  signal W_reg_22_17 : STD_LOGIC;
  signal W_reg_22_16 : STD_LOGIC;
  signal W_reg_22_15 : STD_LOGIC;
  signal W_reg_22_14 : STD_LOGIC;
  signal W_reg_22_13 : STD_LOGIC;
  signal W_reg_22_12 : STD_LOGIC;
  signal W_reg_22_11 : STD_LOGIC;
  signal W_reg_22_10 : STD_LOGIC;
  signal W_reg_22_9 : STD_LOGIC;
  signal W_reg_22_8 : STD_LOGIC;
  signal W_reg_22_7 : STD_LOGIC;
  signal W_reg_22_6 : STD_LOGIC;
  signal W_reg_22_5 : STD_LOGIC;
  signal W_reg_22_4 : STD_LOGIC;
  signal W_reg_22_3 : STD_LOGIC;
  signal W_reg_22_2 : STD_LOGIC;
  signal W_reg_22_1 : STD_LOGIC;
  signal W_reg_22_0 : STD_LOGIC;
  signal W_reg_22_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_22_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_22_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_22_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_22_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_22_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_22_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_22_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_22_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_22_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_22_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_22_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_22_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_22_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_22_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_22_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_22_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_22_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_22_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_22_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_22_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_22_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_22_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_22_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_22_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_22_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_22_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_22_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_22_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_22_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_22_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_23_31 : STD_LOGIC;
  signal W_reg_23_30 : STD_LOGIC;
  signal W_reg_23_29 : STD_LOGIC;
  signal W_reg_23_28 : STD_LOGIC;
  signal W_reg_23_27 : STD_LOGIC;
  signal W_reg_23_26 : STD_LOGIC;
  signal W_reg_23_25 : STD_LOGIC;
  signal W_reg_23_24 : STD_LOGIC;
  signal W_reg_23_23 : STD_LOGIC;
  signal W_reg_23_22 : STD_LOGIC;
  signal W_reg_23_21 : STD_LOGIC;
  signal W_reg_23_20 : STD_LOGIC;
  signal W_reg_23_19 : STD_LOGIC;
  signal W_reg_23_18 : STD_LOGIC;
  signal W_reg_23_17 : STD_LOGIC;
  signal W_reg_23_16 : STD_LOGIC;
  signal W_reg_23_15 : STD_LOGIC;
  signal W_reg_23_14 : STD_LOGIC;
  signal W_reg_23_13 : STD_LOGIC;
  signal W_reg_23_12 : STD_LOGIC;
  signal W_reg_23_11 : STD_LOGIC;
  signal W_reg_23_10 : STD_LOGIC;
  signal W_reg_23_9 : STD_LOGIC;
  signal W_reg_23_8 : STD_LOGIC;
  signal W_reg_23_7 : STD_LOGIC;
  signal W_reg_23_6 : STD_LOGIC;
  signal W_reg_23_5 : STD_LOGIC;
  signal W_reg_23_4 : STD_LOGIC;
  signal W_reg_23_3 : STD_LOGIC;
  signal W_reg_23_2 : STD_LOGIC;
  signal W_reg_23_1 : STD_LOGIC;
  signal W_reg_23_0 : STD_LOGIC;
  signal W_reg_23_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_23_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_23_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_23_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_23_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_23_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_23_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_23_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_23_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_23_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_23_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_23_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_23_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_23_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_23_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_23_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_23_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_23_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_23_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_23_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_23_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_23_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_23_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_23_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_23_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_23_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_23_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_23_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_23_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_23_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_23_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_24_31 : STD_LOGIC;
  signal W_reg_24_30 : STD_LOGIC;
  signal W_reg_24_29 : STD_LOGIC;
  signal W_reg_24_28 : STD_LOGIC;
  signal W_reg_24_27 : STD_LOGIC;
  signal W_reg_24_26 : STD_LOGIC;
  signal W_reg_24_25 : STD_LOGIC;
  signal W_reg_24_24 : STD_LOGIC;
  signal W_reg_24_23 : STD_LOGIC;
  signal W_reg_24_22 : STD_LOGIC;
  signal W_reg_24_21 : STD_LOGIC;
  signal W_reg_24_20 : STD_LOGIC;
  signal W_reg_24_19 : STD_LOGIC;
  signal W_reg_24_18 : STD_LOGIC;
  signal W_reg_24_17 : STD_LOGIC;
  signal W_reg_24_16 : STD_LOGIC;
  signal W_reg_24_15 : STD_LOGIC;
  signal W_reg_24_14 : STD_LOGIC;
  signal W_reg_24_13 : STD_LOGIC;
  signal W_reg_24_12 : STD_LOGIC;
  signal W_reg_24_11 : STD_LOGIC;
  signal W_reg_24_10 : STD_LOGIC;
  signal W_reg_24_9 : STD_LOGIC;
  signal W_reg_24_8 : STD_LOGIC;
  signal W_reg_24_7 : STD_LOGIC;
  signal W_reg_24_6 : STD_LOGIC;
  signal W_reg_24_5 : STD_LOGIC;
  signal W_reg_24_4 : STD_LOGIC;
  signal W_reg_24_3 : STD_LOGIC;
  signal W_reg_24_2 : STD_LOGIC;
  signal W_reg_24_1 : STD_LOGIC;
  signal W_reg_24_0 : STD_LOGIC;
  signal W_reg_24_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_24_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_24_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_24_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_24_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_24_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_24_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_24_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_24_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_24_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_24_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_24_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_24_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_24_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_24_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_24_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_24_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_24_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_24_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_24_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_24_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_24_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_24_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_24_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_24_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_24_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_24_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_24_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_24_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_24_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_24_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_25_31 : STD_LOGIC;
  signal W_reg_25_30 : STD_LOGIC;
  signal W_reg_25_29 : STD_LOGIC;
  signal W_reg_25_28 : STD_LOGIC;
  signal W_reg_25_27 : STD_LOGIC;
  signal W_reg_25_26 : STD_LOGIC;
  signal W_reg_25_25 : STD_LOGIC;
  signal W_reg_25_24 : STD_LOGIC;
  signal W_reg_25_23 : STD_LOGIC;
  signal W_reg_25_22 : STD_LOGIC;
  signal W_reg_25_21 : STD_LOGIC;
  signal W_reg_25_20 : STD_LOGIC;
  signal W_reg_25_19 : STD_LOGIC;
  signal W_reg_25_18 : STD_LOGIC;
  signal W_reg_25_17 : STD_LOGIC;
  signal W_reg_25_16 : STD_LOGIC;
  signal W_reg_25_15 : STD_LOGIC;
  signal W_reg_25_14 : STD_LOGIC;
  signal W_reg_25_13 : STD_LOGIC;
  signal W_reg_25_12 : STD_LOGIC;
  signal W_reg_25_11 : STD_LOGIC;
  signal W_reg_25_10 : STD_LOGIC;
  signal W_reg_25_9 : STD_LOGIC;
  signal W_reg_25_8 : STD_LOGIC;
  signal W_reg_25_7 : STD_LOGIC;
  signal W_reg_25_6 : STD_LOGIC;
  signal W_reg_25_5 : STD_LOGIC;
  signal W_reg_25_4 : STD_LOGIC;
  signal W_reg_25_3 : STD_LOGIC;
  signal W_reg_25_2 : STD_LOGIC;
  signal W_reg_25_1 : STD_LOGIC;
  signal W_reg_25_0 : STD_LOGIC;
  signal W_reg_25_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_25_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_25_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_25_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_25_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_25_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_25_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_25_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_25_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_25_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_25_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_25_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_25_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_25_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_25_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_25_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_25_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_25_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_25_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_25_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_25_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_25_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_25_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_25_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_25_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_25_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_25_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_25_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_25_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_25_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_25_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_26_31 : STD_LOGIC;
  signal W_reg_26_30 : STD_LOGIC;
  signal W_reg_26_29 : STD_LOGIC;
  signal W_reg_26_28 : STD_LOGIC;
  signal W_reg_26_27 : STD_LOGIC;
  signal W_reg_26_26 : STD_LOGIC;
  signal W_reg_26_25 : STD_LOGIC;
  signal W_reg_26_24 : STD_LOGIC;
  signal W_reg_26_23 : STD_LOGIC;
  signal W_reg_26_22 : STD_LOGIC;
  signal W_reg_26_21 : STD_LOGIC;
  signal W_reg_26_20 : STD_LOGIC;
  signal W_reg_26_19 : STD_LOGIC;
  signal W_reg_26_18 : STD_LOGIC;
  signal W_reg_26_17 : STD_LOGIC;
  signal W_reg_26_16 : STD_LOGIC;
  signal W_reg_26_15 : STD_LOGIC;
  signal W_reg_26_14 : STD_LOGIC;
  signal W_reg_26_13 : STD_LOGIC;
  signal W_reg_26_12 : STD_LOGIC;
  signal W_reg_26_11 : STD_LOGIC;
  signal W_reg_26_10 : STD_LOGIC;
  signal W_reg_26_9 : STD_LOGIC;
  signal W_reg_26_8 : STD_LOGIC;
  signal W_reg_26_7 : STD_LOGIC;
  signal W_reg_26_6 : STD_LOGIC;
  signal W_reg_26_5 : STD_LOGIC;
  signal W_reg_26_4 : STD_LOGIC;
  signal W_reg_26_3 : STD_LOGIC;
  signal W_reg_26_2 : STD_LOGIC;
  signal W_reg_26_1 : STD_LOGIC;
  signal W_reg_26_0 : STD_LOGIC;
  signal W_reg_26_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_26_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_26_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_26_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_26_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_26_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_26_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_26_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_26_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_26_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_26_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_26_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_26_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_26_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_26_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_26_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_26_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_26_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_26_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_26_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_26_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_26_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_26_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_26_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_26_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_26_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_26_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_26_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_26_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_26_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_26_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_27_31 : STD_LOGIC;
  signal W_reg_27_30 : STD_LOGIC;
  signal W_reg_27_29 : STD_LOGIC;
  signal W_reg_27_28 : STD_LOGIC;
  signal W_reg_27_27 : STD_LOGIC;
  signal W_reg_27_26 : STD_LOGIC;
  signal W_reg_27_25 : STD_LOGIC;
  signal W_reg_27_24 : STD_LOGIC;
  signal W_reg_27_23 : STD_LOGIC;
  signal W_reg_27_22 : STD_LOGIC;
  signal W_reg_27_21 : STD_LOGIC;
  signal W_reg_27_20 : STD_LOGIC;
  signal W_reg_27_19 : STD_LOGIC;
  signal W_reg_27_18 : STD_LOGIC;
  signal W_reg_27_17 : STD_LOGIC;
  signal W_reg_27_16 : STD_LOGIC;
  signal W_reg_27_15 : STD_LOGIC;
  signal W_reg_27_14 : STD_LOGIC;
  signal W_reg_27_13 : STD_LOGIC;
  signal W_reg_27_12 : STD_LOGIC;
  signal W_reg_27_11 : STD_LOGIC;
  signal W_reg_27_10 : STD_LOGIC;
  signal W_reg_27_9 : STD_LOGIC;
  signal W_reg_27_8 : STD_LOGIC;
  signal W_reg_27_7 : STD_LOGIC;
  signal W_reg_27_6 : STD_LOGIC;
  signal W_reg_27_5 : STD_LOGIC;
  signal W_reg_27_4 : STD_LOGIC;
  signal W_reg_27_3 : STD_LOGIC;
  signal W_reg_27_2 : STD_LOGIC;
  signal W_reg_27_1 : STD_LOGIC;
  signal W_reg_27_0 : STD_LOGIC;
  signal W_reg_27_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_27_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_27_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_27_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_27_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_27_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_27_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_27_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_27_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_27_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_27_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_27_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_27_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_27_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_27_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_27_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_27_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_27_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_27_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_27_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_27_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_27_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_27_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_27_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_27_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_27_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_27_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_27_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_27_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_27_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_27_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_28_31 : STD_LOGIC;
  signal W_reg_28_30 : STD_LOGIC;
  signal W_reg_28_29 : STD_LOGIC;
  signal W_reg_28_28 : STD_LOGIC;
  signal W_reg_28_27 : STD_LOGIC;
  signal W_reg_28_26 : STD_LOGIC;
  signal W_reg_28_25 : STD_LOGIC;
  signal W_reg_28_24 : STD_LOGIC;
  signal W_reg_28_23 : STD_LOGIC;
  signal W_reg_28_22 : STD_LOGIC;
  signal W_reg_28_21 : STD_LOGIC;
  signal W_reg_28_20 : STD_LOGIC;
  signal W_reg_28_19 : STD_LOGIC;
  signal W_reg_28_18 : STD_LOGIC;
  signal W_reg_28_17 : STD_LOGIC;
  signal W_reg_28_16 : STD_LOGIC;
  signal W_reg_28_15 : STD_LOGIC;
  signal W_reg_28_14 : STD_LOGIC;
  signal W_reg_28_13 : STD_LOGIC;
  signal W_reg_28_12 : STD_LOGIC;
  signal W_reg_28_11 : STD_LOGIC;
  signal W_reg_28_10 : STD_LOGIC;
  signal W_reg_28_9 : STD_LOGIC;
  signal W_reg_28_8 : STD_LOGIC;
  signal W_reg_28_7 : STD_LOGIC;
  signal W_reg_28_6 : STD_LOGIC;
  signal W_reg_28_5 : STD_LOGIC;
  signal W_reg_28_4 : STD_LOGIC;
  signal W_reg_28_3 : STD_LOGIC;
  signal W_reg_28_2 : STD_LOGIC;
  signal W_reg_28_1 : STD_LOGIC;
  signal W_reg_28_0 : STD_LOGIC;
  signal W_reg_28_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_28_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_28_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_28_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_28_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_28_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_28_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_28_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_28_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_28_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_28_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_28_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_28_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_28_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_28_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_28_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_28_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_28_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_28_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_28_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_28_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_28_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_28_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_28_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_28_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_28_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_28_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_28_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_28_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_28_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_28_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_29_31 : STD_LOGIC;
  signal W_reg_29_30 : STD_LOGIC;
  signal W_reg_29_29 : STD_LOGIC;
  signal W_reg_29_28 : STD_LOGIC;
  signal W_reg_29_27 : STD_LOGIC;
  signal W_reg_29_26 : STD_LOGIC;
  signal W_reg_29_25 : STD_LOGIC;
  signal W_reg_29_24 : STD_LOGIC;
  signal W_reg_29_23 : STD_LOGIC;
  signal W_reg_29_22 : STD_LOGIC;
  signal W_reg_29_21 : STD_LOGIC;
  signal W_reg_29_20 : STD_LOGIC;
  signal W_reg_29_19 : STD_LOGIC;
  signal W_reg_29_18 : STD_LOGIC;
  signal W_reg_29_17 : STD_LOGIC;
  signal W_reg_29_16 : STD_LOGIC;
  signal W_reg_29_15 : STD_LOGIC;
  signal W_reg_29_14 : STD_LOGIC;
  signal W_reg_29_13 : STD_LOGIC;
  signal W_reg_29_12 : STD_LOGIC;
  signal W_reg_29_11 : STD_LOGIC;
  signal W_reg_29_10 : STD_LOGIC;
  signal W_reg_29_9 : STD_LOGIC;
  signal W_reg_29_8 : STD_LOGIC;
  signal W_reg_29_7 : STD_LOGIC;
  signal W_reg_29_6 : STD_LOGIC;
  signal W_reg_29_5 : STD_LOGIC;
  signal W_reg_29_4 : STD_LOGIC;
  signal W_reg_29_3 : STD_LOGIC;
  signal W_reg_29_2 : STD_LOGIC;
  signal W_reg_29_1 : STD_LOGIC;
  signal W_reg_29_0 : STD_LOGIC;
  signal W_reg_29_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_29_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_29_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_29_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_29_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_29_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_29_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_29_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_29_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_29_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_29_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_29_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_29_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_29_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_29_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_29_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_29_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_29_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_29_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_29_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_29_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_29_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_29_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_29_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_29_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_29_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_29_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_29_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_29_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_29_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_29_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_2_31 : STD_LOGIC;
  signal W_reg_2_30 : STD_LOGIC;
  signal W_reg_2_29 : STD_LOGIC;
  signal W_reg_2_28 : STD_LOGIC;
  signal W_reg_2_27 : STD_LOGIC;
  signal W_reg_2_26 : STD_LOGIC;
  signal W_reg_2_25 : STD_LOGIC;
  signal W_reg_2_24 : STD_LOGIC;
  signal W_reg_2_23 : STD_LOGIC;
  signal W_reg_2_22 : STD_LOGIC;
  signal W_reg_2_21 : STD_LOGIC;
  signal W_reg_2_20 : STD_LOGIC;
  signal W_reg_2_19 : STD_LOGIC;
  signal W_reg_2_18 : STD_LOGIC;
  signal W_reg_2_17 : STD_LOGIC;
  signal W_reg_2_16 : STD_LOGIC;
  signal W_reg_2_15 : STD_LOGIC;
  signal W_reg_2_14 : STD_LOGIC;
  signal W_reg_2_13 : STD_LOGIC;
  signal W_reg_2_12 : STD_LOGIC;
  signal W_reg_2_11 : STD_LOGIC;
  signal W_reg_2_10 : STD_LOGIC;
  signal W_reg_2_9 : STD_LOGIC;
  signal W_reg_2_8 : STD_LOGIC;
  signal W_reg_2_7 : STD_LOGIC;
  signal W_reg_2_6 : STD_LOGIC;
  signal W_reg_2_5 : STD_LOGIC;
  signal W_reg_2_4 : STD_LOGIC;
  signal W_reg_2_3 : STD_LOGIC;
  signal W_reg_2_2 : STD_LOGIC;
  signal W_reg_2_1 : STD_LOGIC;
  signal W_reg_2_0 : STD_LOGIC;
  signal W_reg_30_31 : STD_LOGIC;
  signal W_reg_30_30 : STD_LOGIC;
  signal W_reg_30_29 : STD_LOGIC;
  signal W_reg_30_28 : STD_LOGIC;
  signal W_reg_30_27 : STD_LOGIC;
  signal W_reg_30_26 : STD_LOGIC;
  signal W_reg_30_25 : STD_LOGIC;
  signal W_reg_30_24 : STD_LOGIC;
  signal W_reg_30_23 : STD_LOGIC;
  signal W_reg_30_22 : STD_LOGIC;
  signal W_reg_30_21 : STD_LOGIC;
  signal W_reg_30_20 : STD_LOGIC;
  signal W_reg_30_19 : STD_LOGIC;
  signal W_reg_30_18 : STD_LOGIC;
  signal W_reg_30_17 : STD_LOGIC;
  signal W_reg_30_16 : STD_LOGIC;
  signal W_reg_30_15 : STD_LOGIC;
  signal W_reg_30_14 : STD_LOGIC;
  signal W_reg_30_13 : STD_LOGIC;
  signal W_reg_30_12 : STD_LOGIC;
  signal W_reg_30_11 : STD_LOGIC;
  signal W_reg_30_10 : STD_LOGIC;
  signal W_reg_30_9 : STD_LOGIC;
  signal W_reg_30_8 : STD_LOGIC;
  signal W_reg_30_7 : STD_LOGIC;
  signal W_reg_30_6 : STD_LOGIC;
  signal W_reg_30_5 : STD_LOGIC;
  signal W_reg_30_4 : STD_LOGIC;
  signal W_reg_30_3 : STD_LOGIC;
  signal W_reg_30_2 : STD_LOGIC;
  signal W_reg_30_1 : STD_LOGIC;
  signal W_reg_30_0 : STD_LOGIC;
  signal W_reg_30_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_30_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_30_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_30_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_30_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_30_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_30_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_30_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_30_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_30_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_30_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_30_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_30_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_30_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_30_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_30_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_30_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_30_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_30_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_30_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_30_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_30_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_30_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_30_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_30_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_30_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_30_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_30_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_30_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_30_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_30_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_31_31 : STD_LOGIC;
  signal W_reg_31_30 : STD_LOGIC;
  signal W_reg_31_29 : STD_LOGIC;
  signal W_reg_31_28 : STD_LOGIC;
  signal W_reg_31_27 : STD_LOGIC;
  signal W_reg_31_26 : STD_LOGIC;
  signal W_reg_31_25 : STD_LOGIC;
  signal W_reg_31_24 : STD_LOGIC;
  signal W_reg_31_23 : STD_LOGIC;
  signal W_reg_31_22 : STD_LOGIC;
  signal W_reg_31_21 : STD_LOGIC;
  signal W_reg_31_20 : STD_LOGIC;
  signal W_reg_31_19 : STD_LOGIC;
  signal W_reg_31_18 : STD_LOGIC;
  signal W_reg_31_17 : STD_LOGIC;
  signal W_reg_31_16 : STD_LOGIC;
  signal W_reg_31_15 : STD_LOGIC;
  signal W_reg_31_14 : STD_LOGIC;
  signal W_reg_31_13 : STD_LOGIC;
  signal W_reg_31_12 : STD_LOGIC;
  signal W_reg_31_11 : STD_LOGIC;
  signal W_reg_31_10 : STD_LOGIC;
  signal W_reg_31_9 : STD_LOGIC;
  signal W_reg_31_8 : STD_LOGIC;
  signal W_reg_31_7 : STD_LOGIC;
  signal W_reg_31_6 : STD_LOGIC;
  signal W_reg_31_5 : STD_LOGIC;
  signal W_reg_31_4 : STD_LOGIC;
  signal W_reg_31_3 : STD_LOGIC;
  signal W_reg_31_2 : STD_LOGIC;
  signal W_reg_31_1 : STD_LOGIC;
  signal W_reg_31_0 : STD_LOGIC;
  signal W_reg_31_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_31_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_31_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_31_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_31_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_31_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_31_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_31_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_31_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_31_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_31_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_31_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_31_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_31_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_31_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_31_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_31_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_31_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_31_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_31_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_31_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_31_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_31_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_31_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_31_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_31_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_31_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_31_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_31_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_31_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_31_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_32_31 : STD_LOGIC;
  signal W_reg_32_30 : STD_LOGIC;
  signal W_reg_32_29 : STD_LOGIC;
  signal W_reg_32_28 : STD_LOGIC;
  signal W_reg_32_27 : STD_LOGIC;
  signal W_reg_32_26 : STD_LOGIC;
  signal W_reg_32_25 : STD_LOGIC;
  signal W_reg_32_24 : STD_LOGIC;
  signal W_reg_32_23 : STD_LOGIC;
  signal W_reg_32_22 : STD_LOGIC;
  signal W_reg_32_21 : STD_LOGIC;
  signal W_reg_32_20 : STD_LOGIC;
  signal W_reg_32_19 : STD_LOGIC;
  signal W_reg_32_18 : STD_LOGIC;
  signal W_reg_32_17 : STD_LOGIC;
  signal W_reg_32_16 : STD_LOGIC;
  signal W_reg_32_15 : STD_LOGIC;
  signal W_reg_32_14 : STD_LOGIC;
  signal W_reg_32_13 : STD_LOGIC;
  signal W_reg_32_12 : STD_LOGIC;
  signal W_reg_32_11 : STD_LOGIC;
  signal W_reg_32_10 : STD_LOGIC;
  signal W_reg_32_9 : STD_LOGIC;
  signal W_reg_32_8 : STD_LOGIC;
  signal W_reg_32_7 : STD_LOGIC;
  signal W_reg_32_6 : STD_LOGIC;
  signal W_reg_32_5 : STD_LOGIC;
  signal W_reg_32_4 : STD_LOGIC;
  signal W_reg_32_3 : STD_LOGIC;
  signal W_reg_32_2 : STD_LOGIC;
  signal W_reg_32_1 : STD_LOGIC;
  signal W_reg_32_0 : STD_LOGIC;
  signal W_reg_32_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_32_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_32_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_32_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_32_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_32_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_32_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_32_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_32_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_32_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_32_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_32_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_32_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_32_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_32_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_32_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_32_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_32_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_32_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_32_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_32_31_i_2_n_1 : STD_LOGIC;
  signal W_reg_32_31_i_2_n_2 : STD_LOGIC;
  signal W_reg_32_31_i_2_n_3 : STD_LOGIC;
  signal W_reg_32_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_32_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_32_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_32_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_32_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_32_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_32_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_32_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_33_31 : STD_LOGIC;
  signal W_reg_33_30 : STD_LOGIC;
  signal W_reg_33_29 : STD_LOGIC;
  signal W_reg_33_28 : STD_LOGIC;
  signal W_reg_33_27 : STD_LOGIC;
  signal W_reg_33_26 : STD_LOGIC;
  signal W_reg_33_25 : STD_LOGIC;
  signal W_reg_33_24 : STD_LOGIC;
  signal W_reg_33_23 : STD_LOGIC;
  signal W_reg_33_22 : STD_LOGIC;
  signal W_reg_33_21 : STD_LOGIC;
  signal W_reg_33_20 : STD_LOGIC;
  signal W_reg_33_19 : STD_LOGIC;
  signal W_reg_33_18 : STD_LOGIC;
  signal W_reg_33_17 : STD_LOGIC;
  signal W_reg_33_16 : STD_LOGIC;
  signal W_reg_33_15 : STD_LOGIC;
  signal W_reg_33_14 : STD_LOGIC;
  signal W_reg_33_13 : STD_LOGIC;
  signal W_reg_33_12 : STD_LOGIC;
  signal W_reg_33_11 : STD_LOGIC;
  signal W_reg_33_10 : STD_LOGIC;
  signal W_reg_33_9 : STD_LOGIC;
  signal W_reg_33_8 : STD_LOGIC;
  signal W_reg_33_7 : STD_LOGIC;
  signal W_reg_33_6 : STD_LOGIC;
  signal W_reg_33_5 : STD_LOGIC;
  signal W_reg_33_4 : STD_LOGIC;
  signal W_reg_33_3 : STD_LOGIC;
  signal W_reg_33_2 : STD_LOGIC;
  signal W_reg_33_1 : STD_LOGIC;
  signal W_reg_33_0 : STD_LOGIC;
  signal W_reg_33_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_33_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_33_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_33_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_33_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_33_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_33_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_33_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_33_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_33_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_33_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_33_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_33_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_33_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_33_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_33_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_33_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_33_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_33_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_33_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_33_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_33_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_33_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_33_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_33_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_33_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_33_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_33_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_33_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_33_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_33_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_34_31 : STD_LOGIC;
  signal W_reg_34_30 : STD_LOGIC;
  signal W_reg_34_29 : STD_LOGIC;
  signal W_reg_34_28 : STD_LOGIC;
  signal W_reg_34_27 : STD_LOGIC;
  signal W_reg_34_26 : STD_LOGIC;
  signal W_reg_34_25 : STD_LOGIC;
  signal W_reg_34_24 : STD_LOGIC;
  signal W_reg_34_23 : STD_LOGIC;
  signal W_reg_34_22 : STD_LOGIC;
  signal W_reg_34_21 : STD_LOGIC;
  signal W_reg_34_20 : STD_LOGIC;
  signal W_reg_34_19 : STD_LOGIC;
  signal W_reg_34_18 : STD_LOGIC;
  signal W_reg_34_17 : STD_LOGIC;
  signal W_reg_34_16 : STD_LOGIC;
  signal W_reg_34_15 : STD_LOGIC;
  signal W_reg_34_14 : STD_LOGIC;
  signal W_reg_34_13 : STD_LOGIC;
  signal W_reg_34_12 : STD_LOGIC;
  signal W_reg_34_11 : STD_LOGIC;
  signal W_reg_34_10 : STD_LOGIC;
  signal W_reg_34_9 : STD_LOGIC;
  signal W_reg_34_8 : STD_LOGIC;
  signal W_reg_34_7 : STD_LOGIC;
  signal W_reg_34_6 : STD_LOGIC;
  signal W_reg_34_5 : STD_LOGIC;
  signal W_reg_34_4 : STD_LOGIC;
  signal W_reg_34_3 : STD_LOGIC;
  signal W_reg_34_2 : STD_LOGIC;
  signal W_reg_34_1 : STD_LOGIC;
  signal W_reg_34_0 : STD_LOGIC;
  signal W_reg_34_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_34_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_34_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_34_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_34_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_34_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_34_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_34_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_34_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_34_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_34_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_34_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_34_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_34_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_34_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_34_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_34_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_34_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_34_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_34_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_34_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_34_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_34_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_34_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_34_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_34_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_34_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_34_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_34_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_34_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_34_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_35_31 : STD_LOGIC;
  signal W_reg_35_30 : STD_LOGIC;
  signal W_reg_35_29 : STD_LOGIC;
  signal W_reg_35_28 : STD_LOGIC;
  signal W_reg_35_27 : STD_LOGIC;
  signal W_reg_35_26 : STD_LOGIC;
  signal W_reg_35_25 : STD_LOGIC;
  signal W_reg_35_24 : STD_LOGIC;
  signal W_reg_35_23 : STD_LOGIC;
  signal W_reg_35_22 : STD_LOGIC;
  signal W_reg_35_21 : STD_LOGIC;
  signal W_reg_35_20 : STD_LOGIC;
  signal W_reg_35_19 : STD_LOGIC;
  signal W_reg_35_18 : STD_LOGIC;
  signal W_reg_35_17 : STD_LOGIC;
  signal W_reg_35_16 : STD_LOGIC;
  signal W_reg_35_15 : STD_LOGIC;
  signal W_reg_35_14 : STD_LOGIC;
  signal W_reg_35_13 : STD_LOGIC;
  signal W_reg_35_12 : STD_LOGIC;
  signal W_reg_35_11 : STD_LOGIC;
  signal W_reg_35_10 : STD_LOGIC;
  signal W_reg_35_9 : STD_LOGIC;
  signal W_reg_35_8 : STD_LOGIC;
  signal W_reg_35_7 : STD_LOGIC;
  signal W_reg_35_6 : STD_LOGIC;
  signal W_reg_35_5 : STD_LOGIC;
  signal W_reg_35_4 : STD_LOGIC;
  signal W_reg_35_3 : STD_LOGIC;
  signal W_reg_35_2 : STD_LOGIC;
  signal W_reg_35_1 : STD_LOGIC;
  signal W_reg_35_0 : STD_LOGIC;
  signal W_reg_35_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_35_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_35_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_35_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_35_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_35_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_35_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_35_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_35_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_35_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_35_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_35_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_35_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_35_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_35_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_35_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_35_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_35_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_35_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_35_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_35_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_35_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_35_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_35_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_35_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_35_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_35_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_35_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_35_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_35_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_35_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_36_31 : STD_LOGIC;
  signal W_reg_36_30 : STD_LOGIC;
  signal W_reg_36_29 : STD_LOGIC;
  signal W_reg_36_28 : STD_LOGIC;
  signal W_reg_36_27 : STD_LOGIC;
  signal W_reg_36_26 : STD_LOGIC;
  signal W_reg_36_25 : STD_LOGIC;
  signal W_reg_36_24 : STD_LOGIC;
  signal W_reg_36_23 : STD_LOGIC;
  signal W_reg_36_22 : STD_LOGIC;
  signal W_reg_36_21 : STD_LOGIC;
  signal W_reg_36_20 : STD_LOGIC;
  signal W_reg_36_19 : STD_LOGIC;
  signal W_reg_36_18 : STD_LOGIC;
  signal W_reg_36_17 : STD_LOGIC;
  signal W_reg_36_16 : STD_LOGIC;
  signal W_reg_36_15 : STD_LOGIC;
  signal W_reg_36_14 : STD_LOGIC;
  signal W_reg_36_13 : STD_LOGIC;
  signal W_reg_36_12 : STD_LOGIC;
  signal W_reg_36_11 : STD_LOGIC;
  signal W_reg_36_10 : STD_LOGIC;
  signal W_reg_36_9 : STD_LOGIC;
  signal W_reg_36_8 : STD_LOGIC;
  signal W_reg_36_7 : STD_LOGIC;
  signal W_reg_36_6 : STD_LOGIC;
  signal W_reg_36_5 : STD_LOGIC;
  signal W_reg_36_4 : STD_LOGIC;
  signal W_reg_36_3 : STD_LOGIC;
  signal W_reg_36_2 : STD_LOGIC;
  signal W_reg_36_1 : STD_LOGIC;
  signal W_reg_36_0 : STD_LOGIC;
  signal W_reg_36_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_36_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_36_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_36_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_36_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_36_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_36_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_36_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_36_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_36_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_36_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_36_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_36_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_36_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_36_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_36_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_36_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_36_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_36_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_36_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_36_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_36_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_36_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_36_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_36_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_36_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_36_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_36_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_36_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_36_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_36_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_37_31 : STD_LOGIC;
  signal W_reg_37_30 : STD_LOGIC;
  signal W_reg_37_29 : STD_LOGIC;
  signal W_reg_37_28 : STD_LOGIC;
  signal W_reg_37_27 : STD_LOGIC;
  signal W_reg_37_26 : STD_LOGIC;
  signal W_reg_37_25 : STD_LOGIC;
  signal W_reg_37_24 : STD_LOGIC;
  signal W_reg_37_23 : STD_LOGIC;
  signal W_reg_37_22 : STD_LOGIC;
  signal W_reg_37_21 : STD_LOGIC;
  signal W_reg_37_20 : STD_LOGIC;
  signal W_reg_37_19 : STD_LOGIC;
  signal W_reg_37_18 : STD_LOGIC;
  signal W_reg_37_17 : STD_LOGIC;
  signal W_reg_37_16 : STD_LOGIC;
  signal W_reg_37_15 : STD_LOGIC;
  signal W_reg_37_14 : STD_LOGIC;
  signal W_reg_37_13 : STD_LOGIC;
  signal W_reg_37_12 : STD_LOGIC;
  signal W_reg_37_11 : STD_LOGIC;
  signal W_reg_37_10 : STD_LOGIC;
  signal W_reg_37_9 : STD_LOGIC;
  signal W_reg_37_8 : STD_LOGIC;
  signal W_reg_37_7 : STD_LOGIC;
  signal W_reg_37_6 : STD_LOGIC;
  signal W_reg_37_5 : STD_LOGIC;
  signal W_reg_37_4 : STD_LOGIC;
  signal W_reg_37_3 : STD_LOGIC;
  signal W_reg_37_2 : STD_LOGIC;
  signal W_reg_37_1 : STD_LOGIC;
  signal W_reg_37_0 : STD_LOGIC;
  signal W_reg_37_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_37_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_37_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_37_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_37_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_37_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_37_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_37_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_37_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_37_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_37_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_37_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_37_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_37_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_37_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_37_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_37_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_37_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_37_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_37_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_37_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_37_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_37_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_37_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_37_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_37_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_37_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_37_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_37_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_37_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_37_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_38_31 : STD_LOGIC;
  signal W_reg_38_30 : STD_LOGIC;
  signal W_reg_38_29 : STD_LOGIC;
  signal W_reg_38_28 : STD_LOGIC;
  signal W_reg_38_27 : STD_LOGIC;
  signal W_reg_38_26 : STD_LOGIC;
  signal W_reg_38_25 : STD_LOGIC;
  signal W_reg_38_24 : STD_LOGIC;
  signal W_reg_38_23 : STD_LOGIC;
  signal W_reg_38_22 : STD_LOGIC;
  signal W_reg_38_21 : STD_LOGIC;
  signal W_reg_38_20 : STD_LOGIC;
  signal W_reg_38_19 : STD_LOGIC;
  signal W_reg_38_18 : STD_LOGIC;
  signal W_reg_38_17 : STD_LOGIC;
  signal W_reg_38_16 : STD_LOGIC;
  signal W_reg_38_15 : STD_LOGIC;
  signal W_reg_38_14 : STD_LOGIC;
  signal W_reg_38_13 : STD_LOGIC;
  signal W_reg_38_12 : STD_LOGIC;
  signal W_reg_38_11 : STD_LOGIC;
  signal W_reg_38_10 : STD_LOGIC;
  signal W_reg_38_9 : STD_LOGIC;
  signal W_reg_38_8 : STD_LOGIC;
  signal W_reg_38_7 : STD_LOGIC;
  signal W_reg_38_6 : STD_LOGIC;
  signal W_reg_38_5 : STD_LOGIC;
  signal W_reg_38_4 : STD_LOGIC;
  signal W_reg_38_3 : STD_LOGIC;
  signal W_reg_38_2 : STD_LOGIC;
  signal W_reg_38_1 : STD_LOGIC;
  signal W_reg_38_0 : STD_LOGIC;
  signal W_reg_38_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_38_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_38_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_38_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_38_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_38_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_38_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_38_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_38_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_38_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_38_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_38_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_38_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_38_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_38_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_38_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_38_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_38_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_38_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_38_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_38_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_38_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_38_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_38_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_38_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_38_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_38_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_38_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_38_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_38_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_38_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_39_31 : STD_LOGIC;
  signal W_reg_39_30 : STD_LOGIC;
  signal W_reg_39_29 : STD_LOGIC;
  signal W_reg_39_28 : STD_LOGIC;
  signal W_reg_39_27 : STD_LOGIC;
  signal W_reg_39_26 : STD_LOGIC;
  signal W_reg_39_25 : STD_LOGIC;
  signal W_reg_39_24 : STD_LOGIC;
  signal W_reg_39_23 : STD_LOGIC;
  signal W_reg_39_22 : STD_LOGIC;
  signal W_reg_39_21 : STD_LOGIC;
  signal W_reg_39_20 : STD_LOGIC;
  signal W_reg_39_19 : STD_LOGIC;
  signal W_reg_39_18 : STD_LOGIC;
  signal W_reg_39_17 : STD_LOGIC;
  signal W_reg_39_16 : STD_LOGIC;
  signal W_reg_39_15 : STD_LOGIC;
  signal W_reg_39_14 : STD_LOGIC;
  signal W_reg_39_13 : STD_LOGIC;
  signal W_reg_39_12 : STD_LOGIC;
  signal W_reg_39_11 : STD_LOGIC;
  signal W_reg_39_10 : STD_LOGIC;
  signal W_reg_39_9 : STD_LOGIC;
  signal W_reg_39_8 : STD_LOGIC;
  signal W_reg_39_7 : STD_LOGIC;
  signal W_reg_39_6 : STD_LOGIC;
  signal W_reg_39_5 : STD_LOGIC;
  signal W_reg_39_4 : STD_LOGIC;
  signal W_reg_39_3 : STD_LOGIC;
  signal W_reg_39_2 : STD_LOGIC;
  signal W_reg_39_1 : STD_LOGIC;
  signal W_reg_39_0 : STD_LOGIC;
  signal W_reg_39_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_39_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_39_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_39_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_39_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_39_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_39_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_39_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_39_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_39_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_39_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_39_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_39_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_39_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_39_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_39_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_39_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_39_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_39_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_39_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_39_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_39_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_39_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_39_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_39_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_39_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_39_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_39_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_39_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_39_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_39_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_3_31 : STD_LOGIC;
  signal W_reg_3_30 : STD_LOGIC;
  signal W_reg_3_29 : STD_LOGIC;
  signal W_reg_3_28 : STD_LOGIC;
  signal W_reg_3_27 : STD_LOGIC;
  signal W_reg_3_26 : STD_LOGIC;
  signal W_reg_3_25 : STD_LOGIC;
  signal W_reg_3_24 : STD_LOGIC;
  signal W_reg_3_23 : STD_LOGIC;
  signal W_reg_3_22 : STD_LOGIC;
  signal W_reg_3_21 : STD_LOGIC;
  signal W_reg_3_20 : STD_LOGIC;
  signal W_reg_3_19 : STD_LOGIC;
  signal W_reg_3_18 : STD_LOGIC;
  signal W_reg_3_17 : STD_LOGIC;
  signal W_reg_3_16 : STD_LOGIC;
  signal W_reg_3_15 : STD_LOGIC;
  signal W_reg_3_14 : STD_LOGIC;
  signal W_reg_3_13 : STD_LOGIC;
  signal W_reg_3_12 : STD_LOGIC;
  signal W_reg_3_11 : STD_LOGIC;
  signal W_reg_3_10 : STD_LOGIC;
  signal W_reg_3_9 : STD_LOGIC;
  signal W_reg_3_8 : STD_LOGIC;
  signal W_reg_3_7 : STD_LOGIC;
  signal W_reg_3_6 : STD_LOGIC;
  signal W_reg_3_5 : STD_LOGIC;
  signal W_reg_3_4 : STD_LOGIC;
  signal W_reg_3_3 : STD_LOGIC;
  signal W_reg_3_2 : STD_LOGIC;
  signal W_reg_3_1 : STD_LOGIC;
  signal W_reg_3_0 : STD_LOGIC;
  signal W_reg_40_31 : STD_LOGIC;
  signal W_reg_40_30 : STD_LOGIC;
  signal W_reg_40_29 : STD_LOGIC;
  signal W_reg_40_28 : STD_LOGIC;
  signal W_reg_40_27 : STD_LOGIC;
  signal W_reg_40_26 : STD_LOGIC;
  signal W_reg_40_25 : STD_LOGIC;
  signal W_reg_40_24 : STD_LOGIC;
  signal W_reg_40_23 : STD_LOGIC;
  signal W_reg_40_22 : STD_LOGIC;
  signal W_reg_40_21 : STD_LOGIC;
  signal W_reg_40_20 : STD_LOGIC;
  signal W_reg_40_19 : STD_LOGIC;
  signal W_reg_40_18 : STD_LOGIC;
  signal W_reg_40_17 : STD_LOGIC;
  signal W_reg_40_16 : STD_LOGIC;
  signal W_reg_40_15 : STD_LOGIC;
  signal W_reg_40_14 : STD_LOGIC;
  signal W_reg_40_13 : STD_LOGIC;
  signal W_reg_40_12 : STD_LOGIC;
  signal W_reg_40_11 : STD_LOGIC;
  signal W_reg_40_10 : STD_LOGIC;
  signal W_reg_40_9 : STD_LOGIC;
  signal W_reg_40_8 : STD_LOGIC;
  signal W_reg_40_7 : STD_LOGIC;
  signal W_reg_40_6 : STD_LOGIC;
  signal W_reg_40_5 : STD_LOGIC;
  signal W_reg_40_4 : STD_LOGIC;
  signal W_reg_40_3 : STD_LOGIC;
  signal W_reg_40_2 : STD_LOGIC;
  signal W_reg_40_1 : STD_LOGIC;
  signal W_reg_40_0 : STD_LOGIC;
  signal W_reg_40_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_40_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_40_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_40_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_40_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_40_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_40_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_40_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_40_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_40_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_40_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_40_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_40_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_40_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_40_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_40_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_40_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_40_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_40_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_40_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_40_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_40_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_40_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_40_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_40_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_40_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_40_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_40_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_40_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_40_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_40_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_41_31 : STD_LOGIC;
  signal W_reg_41_30 : STD_LOGIC;
  signal W_reg_41_29 : STD_LOGIC;
  signal W_reg_41_28 : STD_LOGIC;
  signal W_reg_41_27 : STD_LOGIC;
  signal W_reg_41_26 : STD_LOGIC;
  signal W_reg_41_25 : STD_LOGIC;
  signal W_reg_41_24 : STD_LOGIC;
  signal W_reg_41_23 : STD_LOGIC;
  signal W_reg_41_22 : STD_LOGIC;
  signal W_reg_41_21 : STD_LOGIC;
  signal W_reg_41_20 : STD_LOGIC;
  signal W_reg_41_19 : STD_LOGIC;
  signal W_reg_41_18 : STD_LOGIC;
  signal W_reg_41_17 : STD_LOGIC;
  signal W_reg_41_16 : STD_LOGIC;
  signal W_reg_41_15 : STD_LOGIC;
  signal W_reg_41_14 : STD_LOGIC;
  signal W_reg_41_13 : STD_LOGIC;
  signal W_reg_41_12 : STD_LOGIC;
  signal W_reg_41_11 : STD_LOGIC;
  signal W_reg_41_10 : STD_LOGIC;
  signal W_reg_41_9 : STD_LOGIC;
  signal W_reg_41_8 : STD_LOGIC;
  signal W_reg_41_7 : STD_LOGIC;
  signal W_reg_41_6 : STD_LOGIC;
  signal W_reg_41_5 : STD_LOGIC;
  signal W_reg_41_4 : STD_LOGIC;
  signal W_reg_41_3 : STD_LOGIC;
  signal W_reg_41_2 : STD_LOGIC;
  signal W_reg_41_1 : STD_LOGIC;
  signal W_reg_41_0 : STD_LOGIC;
  signal W_reg_41_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_41_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_41_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_41_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_41_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_41_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_41_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_41_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_41_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_41_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_41_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_41_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_41_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_41_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_41_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_41_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_41_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_41_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_41_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_41_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_41_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_41_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_41_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_41_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_41_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_41_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_41_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_41_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_41_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_41_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_41_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_42_31 : STD_LOGIC;
  signal W_reg_42_30 : STD_LOGIC;
  signal W_reg_42_29 : STD_LOGIC;
  signal W_reg_42_28 : STD_LOGIC;
  signal W_reg_42_27 : STD_LOGIC;
  signal W_reg_42_26 : STD_LOGIC;
  signal W_reg_42_25 : STD_LOGIC;
  signal W_reg_42_24 : STD_LOGIC;
  signal W_reg_42_23 : STD_LOGIC;
  signal W_reg_42_22 : STD_LOGIC;
  signal W_reg_42_21 : STD_LOGIC;
  signal W_reg_42_20 : STD_LOGIC;
  signal W_reg_42_19 : STD_LOGIC;
  signal W_reg_42_18 : STD_LOGIC;
  signal W_reg_42_17 : STD_LOGIC;
  signal W_reg_42_16 : STD_LOGIC;
  signal W_reg_42_15 : STD_LOGIC;
  signal W_reg_42_14 : STD_LOGIC;
  signal W_reg_42_13 : STD_LOGIC;
  signal W_reg_42_12 : STD_LOGIC;
  signal W_reg_42_11 : STD_LOGIC;
  signal W_reg_42_10 : STD_LOGIC;
  signal W_reg_42_9 : STD_LOGIC;
  signal W_reg_42_8 : STD_LOGIC;
  signal W_reg_42_7 : STD_LOGIC;
  signal W_reg_42_6 : STD_LOGIC;
  signal W_reg_42_5 : STD_LOGIC;
  signal W_reg_42_4 : STD_LOGIC;
  signal W_reg_42_3 : STD_LOGIC;
  signal W_reg_42_2 : STD_LOGIC;
  signal W_reg_42_1 : STD_LOGIC;
  signal W_reg_42_0 : STD_LOGIC;
  signal W_reg_42_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_42_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_42_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_42_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_42_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_42_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_42_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_42_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_42_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_42_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_42_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_42_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_42_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_42_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_42_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_42_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_42_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_42_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_42_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_42_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_42_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_42_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_42_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_42_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_42_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_42_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_42_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_42_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_42_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_42_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_42_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_43_31 : STD_LOGIC;
  signal W_reg_43_30 : STD_LOGIC;
  signal W_reg_43_29 : STD_LOGIC;
  signal W_reg_43_28 : STD_LOGIC;
  signal W_reg_43_27 : STD_LOGIC;
  signal W_reg_43_26 : STD_LOGIC;
  signal W_reg_43_25 : STD_LOGIC;
  signal W_reg_43_24 : STD_LOGIC;
  signal W_reg_43_23 : STD_LOGIC;
  signal W_reg_43_22 : STD_LOGIC;
  signal W_reg_43_21 : STD_LOGIC;
  signal W_reg_43_20 : STD_LOGIC;
  signal W_reg_43_19 : STD_LOGIC;
  signal W_reg_43_18 : STD_LOGIC;
  signal W_reg_43_17 : STD_LOGIC;
  signal W_reg_43_16 : STD_LOGIC;
  signal W_reg_43_15 : STD_LOGIC;
  signal W_reg_43_14 : STD_LOGIC;
  signal W_reg_43_13 : STD_LOGIC;
  signal W_reg_43_12 : STD_LOGIC;
  signal W_reg_43_11 : STD_LOGIC;
  signal W_reg_43_10 : STD_LOGIC;
  signal W_reg_43_9 : STD_LOGIC;
  signal W_reg_43_8 : STD_LOGIC;
  signal W_reg_43_7 : STD_LOGIC;
  signal W_reg_43_6 : STD_LOGIC;
  signal W_reg_43_5 : STD_LOGIC;
  signal W_reg_43_4 : STD_LOGIC;
  signal W_reg_43_3 : STD_LOGIC;
  signal W_reg_43_2 : STD_LOGIC;
  signal W_reg_43_1 : STD_LOGIC;
  signal W_reg_43_0 : STD_LOGIC;
  signal W_reg_43_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_43_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_43_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_43_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_43_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_43_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_43_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_43_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_43_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_43_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_43_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_43_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_43_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_43_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_43_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_43_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_43_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_43_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_43_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_43_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_43_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_43_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_43_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_43_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_43_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_43_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_43_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_43_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_43_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_43_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_43_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_44_31 : STD_LOGIC;
  signal W_reg_44_30 : STD_LOGIC;
  signal W_reg_44_29 : STD_LOGIC;
  signal W_reg_44_28 : STD_LOGIC;
  signal W_reg_44_27 : STD_LOGIC;
  signal W_reg_44_26 : STD_LOGIC;
  signal W_reg_44_25 : STD_LOGIC;
  signal W_reg_44_24 : STD_LOGIC;
  signal W_reg_44_23 : STD_LOGIC;
  signal W_reg_44_22 : STD_LOGIC;
  signal W_reg_44_21 : STD_LOGIC;
  signal W_reg_44_20 : STD_LOGIC;
  signal W_reg_44_19 : STD_LOGIC;
  signal W_reg_44_18 : STD_LOGIC;
  signal W_reg_44_17 : STD_LOGIC;
  signal W_reg_44_16 : STD_LOGIC;
  signal W_reg_44_15 : STD_LOGIC;
  signal W_reg_44_14 : STD_LOGIC;
  signal W_reg_44_13 : STD_LOGIC;
  signal W_reg_44_12 : STD_LOGIC;
  signal W_reg_44_11 : STD_LOGIC;
  signal W_reg_44_10 : STD_LOGIC;
  signal W_reg_44_9 : STD_LOGIC;
  signal W_reg_44_8 : STD_LOGIC;
  signal W_reg_44_7 : STD_LOGIC;
  signal W_reg_44_6 : STD_LOGIC;
  signal W_reg_44_5 : STD_LOGIC;
  signal W_reg_44_4 : STD_LOGIC;
  signal W_reg_44_3 : STD_LOGIC;
  signal W_reg_44_2 : STD_LOGIC;
  signal W_reg_44_1 : STD_LOGIC;
  signal W_reg_44_0 : STD_LOGIC;
  signal W_reg_44_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_44_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_44_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_44_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_44_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_44_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_44_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_44_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_44_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_44_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_44_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_44_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_44_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_44_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_44_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_44_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_44_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_44_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_44_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_44_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_44_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_44_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_44_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_44_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_44_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_44_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_44_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_44_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_44_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_44_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_44_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_45_31 : STD_LOGIC;
  signal W_reg_45_30 : STD_LOGIC;
  signal W_reg_45_29 : STD_LOGIC;
  signal W_reg_45_28 : STD_LOGIC;
  signal W_reg_45_27 : STD_LOGIC;
  signal W_reg_45_26 : STD_LOGIC;
  signal W_reg_45_25 : STD_LOGIC;
  signal W_reg_45_24 : STD_LOGIC;
  signal W_reg_45_23 : STD_LOGIC;
  signal W_reg_45_22 : STD_LOGIC;
  signal W_reg_45_21 : STD_LOGIC;
  signal W_reg_45_20 : STD_LOGIC;
  signal W_reg_45_19 : STD_LOGIC;
  signal W_reg_45_18 : STD_LOGIC;
  signal W_reg_45_17 : STD_LOGIC;
  signal W_reg_45_16 : STD_LOGIC;
  signal W_reg_45_15 : STD_LOGIC;
  signal W_reg_45_14 : STD_LOGIC;
  signal W_reg_45_13 : STD_LOGIC;
  signal W_reg_45_12 : STD_LOGIC;
  signal W_reg_45_11 : STD_LOGIC;
  signal W_reg_45_10 : STD_LOGIC;
  signal W_reg_45_9 : STD_LOGIC;
  signal W_reg_45_8 : STD_LOGIC;
  signal W_reg_45_7 : STD_LOGIC;
  signal W_reg_45_6 : STD_LOGIC;
  signal W_reg_45_5 : STD_LOGIC;
  signal W_reg_45_4 : STD_LOGIC;
  signal W_reg_45_3 : STD_LOGIC;
  signal W_reg_45_2 : STD_LOGIC;
  signal W_reg_45_1 : STD_LOGIC;
  signal W_reg_45_0 : STD_LOGIC;
  signal W_reg_45_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_45_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_45_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_45_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_45_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_45_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_45_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_45_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_45_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_45_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_45_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_45_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_45_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_45_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_45_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_45_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_45_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_45_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_45_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_45_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_45_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_45_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_45_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_45_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_45_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_45_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_45_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_45_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_45_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_45_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_45_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_46_31 : STD_LOGIC;
  signal W_reg_46_30 : STD_LOGIC;
  signal W_reg_46_29 : STD_LOGIC;
  signal W_reg_46_28 : STD_LOGIC;
  signal W_reg_46_27 : STD_LOGIC;
  signal W_reg_46_26 : STD_LOGIC;
  signal W_reg_46_25 : STD_LOGIC;
  signal W_reg_46_24 : STD_LOGIC;
  signal W_reg_46_23 : STD_LOGIC;
  signal W_reg_46_22 : STD_LOGIC;
  signal W_reg_46_21 : STD_LOGIC;
  signal W_reg_46_20 : STD_LOGIC;
  signal W_reg_46_19 : STD_LOGIC;
  signal W_reg_46_18 : STD_LOGIC;
  signal W_reg_46_17 : STD_LOGIC;
  signal W_reg_46_16 : STD_LOGIC;
  signal W_reg_46_15 : STD_LOGIC;
  signal W_reg_46_14 : STD_LOGIC;
  signal W_reg_46_13 : STD_LOGIC;
  signal W_reg_46_12 : STD_LOGIC;
  signal W_reg_46_11 : STD_LOGIC;
  signal W_reg_46_10 : STD_LOGIC;
  signal W_reg_46_9 : STD_LOGIC;
  signal W_reg_46_8 : STD_LOGIC;
  signal W_reg_46_7 : STD_LOGIC;
  signal W_reg_46_6 : STD_LOGIC;
  signal W_reg_46_5 : STD_LOGIC;
  signal W_reg_46_4 : STD_LOGIC;
  signal W_reg_46_3 : STD_LOGIC;
  signal W_reg_46_2 : STD_LOGIC;
  signal W_reg_46_1 : STD_LOGIC;
  signal W_reg_46_0 : STD_LOGIC;
  signal W_reg_46_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_46_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_46_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_46_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_46_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_46_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_46_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_46_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_46_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_46_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_46_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_46_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_46_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_46_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_46_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_46_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_46_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_46_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_46_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_46_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_46_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_46_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_46_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_46_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_46_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_46_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_46_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_46_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_46_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_46_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_46_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_47_31 : STD_LOGIC;
  signal W_reg_47_30 : STD_LOGIC;
  signal W_reg_47_29 : STD_LOGIC;
  signal W_reg_47_28 : STD_LOGIC;
  signal W_reg_47_27 : STD_LOGIC;
  signal W_reg_47_26 : STD_LOGIC;
  signal W_reg_47_25 : STD_LOGIC;
  signal W_reg_47_24 : STD_LOGIC;
  signal W_reg_47_23 : STD_LOGIC;
  signal W_reg_47_22 : STD_LOGIC;
  signal W_reg_47_21 : STD_LOGIC;
  signal W_reg_47_20 : STD_LOGIC;
  signal W_reg_47_19 : STD_LOGIC;
  signal W_reg_47_18 : STD_LOGIC;
  signal W_reg_47_17 : STD_LOGIC;
  signal W_reg_47_16 : STD_LOGIC;
  signal W_reg_47_15 : STD_LOGIC;
  signal W_reg_47_14 : STD_LOGIC;
  signal W_reg_47_13 : STD_LOGIC;
  signal W_reg_47_12 : STD_LOGIC;
  signal W_reg_47_11 : STD_LOGIC;
  signal W_reg_47_10 : STD_LOGIC;
  signal W_reg_47_9 : STD_LOGIC;
  signal W_reg_47_8 : STD_LOGIC;
  signal W_reg_47_7 : STD_LOGIC;
  signal W_reg_47_6 : STD_LOGIC;
  signal W_reg_47_5 : STD_LOGIC;
  signal W_reg_47_4 : STD_LOGIC;
  signal W_reg_47_3 : STD_LOGIC;
  signal W_reg_47_2 : STD_LOGIC;
  signal W_reg_47_1 : STD_LOGIC;
  signal W_reg_47_0 : STD_LOGIC;
  signal W_reg_47_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_47_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_47_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_47_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_47_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_47_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_47_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_47_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_47_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_47_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_47_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_47_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_47_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_47_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_47_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_47_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_47_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_47_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_47_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_47_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_47_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_47_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_47_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_47_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_47_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_47_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_47_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_47_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_47_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_47_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_47_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_48_31 : STD_LOGIC;
  signal W_reg_48_30 : STD_LOGIC;
  signal W_reg_48_29 : STD_LOGIC;
  signal W_reg_48_28 : STD_LOGIC;
  signal W_reg_48_27 : STD_LOGIC;
  signal W_reg_48_26 : STD_LOGIC;
  signal W_reg_48_25 : STD_LOGIC;
  signal W_reg_48_24 : STD_LOGIC;
  signal W_reg_48_23 : STD_LOGIC;
  signal W_reg_48_22 : STD_LOGIC;
  signal W_reg_48_21 : STD_LOGIC;
  signal W_reg_48_20 : STD_LOGIC;
  signal W_reg_48_19 : STD_LOGIC;
  signal W_reg_48_18 : STD_LOGIC;
  signal W_reg_48_17 : STD_LOGIC;
  signal W_reg_48_16 : STD_LOGIC;
  signal W_reg_48_15 : STD_LOGIC;
  signal W_reg_48_14 : STD_LOGIC;
  signal W_reg_48_13 : STD_LOGIC;
  signal W_reg_48_12 : STD_LOGIC;
  signal W_reg_48_11 : STD_LOGIC;
  signal W_reg_48_10 : STD_LOGIC;
  signal W_reg_48_9 : STD_LOGIC;
  signal W_reg_48_8 : STD_LOGIC;
  signal W_reg_48_7 : STD_LOGIC;
  signal W_reg_48_6 : STD_LOGIC;
  signal W_reg_48_5 : STD_LOGIC;
  signal W_reg_48_4 : STD_LOGIC;
  signal W_reg_48_3 : STD_LOGIC;
  signal W_reg_48_2 : STD_LOGIC;
  signal W_reg_48_1 : STD_LOGIC;
  signal W_reg_48_0 : STD_LOGIC;
  signal W_reg_48_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_48_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_48_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_48_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_48_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_48_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_48_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_48_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_48_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_48_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_48_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_48_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_48_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_48_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_48_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_48_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_48_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_48_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_48_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_48_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_48_31_i_2_n_1 : STD_LOGIC;
  signal W_reg_48_31_i_2_n_2 : STD_LOGIC;
  signal W_reg_48_31_i_2_n_3 : STD_LOGIC;
  signal W_reg_48_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_48_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_48_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_48_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_48_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_48_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_48_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_48_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_49_31 : STD_LOGIC;
  signal W_reg_49_30 : STD_LOGIC;
  signal W_reg_49_29 : STD_LOGIC;
  signal W_reg_49_28 : STD_LOGIC;
  signal W_reg_49_27 : STD_LOGIC;
  signal W_reg_49_26 : STD_LOGIC;
  signal W_reg_49_25 : STD_LOGIC;
  signal W_reg_49_24 : STD_LOGIC;
  signal W_reg_49_23 : STD_LOGIC;
  signal W_reg_49_22 : STD_LOGIC;
  signal W_reg_49_21 : STD_LOGIC;
  signal W_reg_49_20 : STD_LOGIC;
  signal W_reg_49_19 : STD_LOGIC;
  signal W_reg_49_18 : STD_LOGIC;
  signal W_reg_49_17 : STD_LOGIC;
  signal W_reg_49_16 : STD_LOGIC;
  signal W_reg_49_15 : STD_LOGIC;
  signal W_reg_49_14 : STD_LOGIC;
  signal W_reg_49_13 : STD_LOGIC;
  signal W_reg_49_12 : STD_LOGIC;
  signal W_reg_49_11 : STD_LOGIC;
  signal W_reg_49_10 : STD_LOGIC;
  signal W_reg_49_9 : STD_LOGIC;
  signal W_reg_49_8 : STD_LOGIC;
  signal W_reg_49_7 : STD_LOGIC;
  signal W_reg_49_6 : STD_LOGIC;
  signal W_reg_49_5 : STD_LOGIC;
  signal W_reg_49_4 : STD_LOGIC;
  signal W_reg_49_3 : STD_LOGIC;
  signal W_reg_49_2 : STD_LOGIC;
  signal W_reg_49_1 : STD_LOGIC;
  signal W_reg_49_0 : STD_LOGIC;
  signal W_reg_49_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_49_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_49_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_49_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_49_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_49_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_49_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_49_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_49_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_49_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_49_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_49_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_49_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_49_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_49_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_49_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_49_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_49_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_49_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_49_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_49_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_49_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_49_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_49_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_49_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_49_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_49_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_49_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_49_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_49_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_49_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_4_31 : STD_LOGIC;
  signal W_reg_4_30 : STD_LOGIC;
  signal W_reg_4_29 : STD_LOGIC;
  signal W_reg_4_28 : STD_LOGIC;
  signal W_reg_4_27 : STD_LOGIC;
  signal W_reg_4_26 : STD_LOGIC;
  signal W_reg_4_25 : STD_LOGIC;
  signal W_reg_4_24 : STD_LOGIC;
  signal W_reg_4_23 : STD_LOGIC;
  signal W_reg_4_22 : STD_LOGIC;
  signal W_reg_4_21 : STD_LOGIC;
  signal W_reg_4_20 : STD_LOGIC;
  signal W_reg_4_19 : STD_LOGIC;
  signal W_reg_4_18 : STD_LOGIC;
  signal W_reg_4_17 : STD_LOGIC;
  signal W_reg_4_16 : STD_LOGIC;
  signal W_reg_4_15 : STD_LOGIC;
  signal W_reg_4_14 : STD_LOGIC;
  signal W_reg_4_13 : STD_LOGIC;
  signal W_reg_4_12 : STD_LOGIC;
  signal W_reg_4_11 : STD_LOGIC;
  signal W_reg_4_10 : STD_LOGIC;
  signal W_reg_4_9 : STD_LOGIC;
  signal W_reg_4_8 : STD_LOGIC;
  signal W_reg_4_7 : STD_LOGIC;
  signal W_reg_4_6 : STD_LOGIC;
  signal W_reg_4_5 : STD_LOGIC;
  signal W_reg_4_4 : STD_LOGIC;
  signal W_reg_4_3 : STD_LOGIC;
  signal W_reg_4_2 : STD_LOGIC;
  signal W_reg_4_1 : STD_LOGIC;
  signal W_reg_4_0 : STD_LOGIC;
  signal W_reg_50_31 : STD_LOGIC;
  signal W_reg_50_30 : STD_LOGIC;
  signal W_reg_50_29 : STD_LOGIC;
  signal W_reg_50_28 : STD_LOGIC;
  signal W_reg_50_27 : STD_LOGIC;
  signal W_reg_50_26 : STD_LOGIC;
  signal W_reg_50_25 : STD_LOGIC;
  signal W_reg_50_24 : STD_LOGIC;
  signal W_reg_50_23 : STD_LOGIC;
  signal W_reg_50_22 : STD_LOGIC;
  signal W_reg_50_21 : STD_LOGIC;
  signal W_reg_50_20 : STD_LOGIC;
  signal W_reg_50_19 : STD_LOGIC;
  signal W_reg_50_18 : STD_LOGIC;
  signal W_reg_50_17 : STD_LOGIC;
  signal W_reg_50_16 : STD_LOGIC;
  signal W_reg_50_15 : STD_LOGIC;
  signal W_reg_50_14 : STD_LOGIC;
  signal W_reg_50_13 : STD_LOGIC;
  signal W_reg_50_12 : STD_LOGIC;
  signal W_reg_50_11 : STD_LOGIC;
  signal W_reg_50_10 : STD_LOGIC;
  signal W_reg_50_9 : STD_LOGIC;
  signal W_reg_50_8 : STD_LOGIC;
  signal W_reg_50_7 : STD_LOGIC;
  signal W_reg_50_6 : STD_LOGIC;
  signal W_reg_50_5 : STD_LOGIC;
  signal W_reg_50_4 : STD_LOGIC;
  signal W_reg_50_3 : STD_LOGIC;
  signal W_reg_50_2 : STD_LOGIC;
  signal W_reg_50_1 : STD_LOGIC;
  signal W_reg_50_0 : STD_LOGIC;
  signal W_reg_50_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_50_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_50_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_50_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_50_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_50_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_50_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_50_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_50_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_50_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_50_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_50_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_50_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_50_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_50_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_50_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_50_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_50_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_50_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_50_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_50_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_50_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_50_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_50_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_50_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_50_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_50_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_50_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_50_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_50_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_50_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_51_31 : STD_LOGIC;
  signal W_reg_51_30 : STD_LOGIC;
  signal W_reg_51_29 : STD_LOGIC;
  signal W_reg_51_28 : STD_LOGIC;
  signal W_reg_51_27 : STD_LOGIC;
  signal W_reg_51_26 : STD_LOGIC;
  signal W_reg_51_25 : STD_LOGIC;
  signal W_reg_51_24 : STD_LOGIC;
  signal W_reg_51_23 : STD_LOGIC;
  signal W_reg_51_22 : STD_LOGIC;
  signal W_reg_51_21 : STD_LOGIC;
  signal W_reg_51_20 : STD_LOGIC;
  signal W_reg_51_19 : STD_LOGIC;
  signal W_reg_51_18 : STD_LOGIC;
  signal W_reg_51_17 : STD_LOGIC;
  signal W_reg_51_16 : STD_LOGIC;
  signal W_reg_51_15 : STD_LOGIC;
  signal W_reg_51_14 : STD_LOGIC;
  signal W_reg_51_13 : STD_LOGIC;
  signal W_reg_51_12 : STD_LOGIC;
  signal W_reg_51_11 : STD_LOGIC;
  signal W_reg_51_10 : STD_LOGIC;
  signal W_reg_51_9 : STD_LOGIC;
  signal W_reg_51_8 : STD_LOGIC;
  signal W_reg_51_7 : STD_LOGIC;
  signal W_reg_51_6 : STD_LOGIC;
  signal W_reg_51_5 : STD_LOGIC;
  signal W_reg_51_4 : STD_LOGIC;
  signal W_reg_51_3 : STD_LOGIC;
  signal W_reg_51_2 : STD_LOGIC;
  signal W_reg_51_1 : STD_LOGIC;
  signal W_reg_51_0 : STD_LOGIC;
  signal W_reg_51_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_51_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_51_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_51_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_51_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_51_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_51_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_51_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_51_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_51_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_51_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_51_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_51_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_51_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_51_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_51_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_51_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_51_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_51_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_51_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_51_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_51_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_51_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_51_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_51_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_51_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_51_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_51_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_51_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_51_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_51_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_52_31 : STD_LOGIC;
  signal W_reg_52_30 : STD_LOGIC;
  signal W_reg_52_29 : STD_LOGIC;
  signal W_reg_52_28 : STD_LOGIC;
  signal W_reg_52_27 : STD_LOGIC;
  signal W_reg_52_26 : STD_LOGIC;
  signal W_reg_52_25 : STD_LOGIC;
  signal W_reg_52_24 : STD_LOGIC;
  signal W_reg_52_23 : STD_LOGIC;
  signal W_reg_52_22 : STD_LOGIC;
  signal W_reg_52_21 : STD_LOGIC;
  signal W_reg_52_20 : STD_LOGIC;
  signal W_reg_52_19 : STD_LOGIC;
  signal W_reg_52_18 : STD_LOGIC;
  signal W_reg_52_17 : STD_LOGIC;
  signal W_reg_52_16 : STD_LOGIC;
  signal W_reg_52_15 : STD_LOGIC;
  signal W_reg_52_14 : STD_LOGIC;
  signal W_reg_52_13 : STD_LOGIC;
  signal W_reg_52_12 : STD_LOGIC;
  signal W_reg_52_11 : STD_LOGIC;
  signal W_reg_52_10 : STD_LOGIC;
  signal W_reg_52_9 : STD_LOGIC;
  signal W_reg_52_8 : STD_LOGIC;
  signal W_reg_52_7 : STD_LOGIC;
  signal W_reg_52_6 : STD_LOGIC;
  signal W_reg_52_5 : STD_LOGIC;
  signal W_reg_52_4 : STD_LOGIC;
  signal W_reg_52_3 : STD_LOGIC;
  signal W_reg_52_2 : STD_LOGIC;
  signal W_reg_52_1 : STD_LOGIC;
  signal W_reg_52_0 : STD_LOGIC;
  signal W_reg_52_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_52_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_52_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_52_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_52_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_52_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_52_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_52_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_52_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_52_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_52_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_52_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_52_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_52_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_52_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_52_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_52_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_52_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_52_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_52_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_52_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_52_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_52_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_52_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_52_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_52_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_52_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_52_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_52_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_52_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_52_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_53_31 : STD_LOGIC;
  signal W_reg_53_30 : STD_LOGIC;
  signal W_reg_53_29 : STD_LOGIC;
  signal W_reg_53_28 : STD_LOGIC;
  signal W_reg_53_27 : STD_LOGIC;
  signal W_reg_53_26 : STD_LOGIC;
  signal W_reg_53_25 : STD_LOGIC;
  signal W_reg_53_24 : STD_LOGIC;
  signal W_reg_53_23 : STD_LOGIC;
  signal W_reg_53_22 : STD_LOGIC;
  signal W_reg_53_21 : STD_LOGIC;
  signal W_reg_53_20 : STD_LOGIC;
  signal W_reg_53_19 : STD_LOGIC;
  signal W_reg_53_18 : STD_LOGIC;
  signal W_reg_53_17 : STD_LOGIC;
  signal W_reg_53_16 : STD_LOGIC;
  signal W_reg_53_15 : STD_LOGIC;
  signal W_reg_53_14 : STD_LOGIC;
  signal W_reg_53_13 : STD_LOGIC;
  signal W_reg_53_12 : STD_LOGIC;
  signal W_reg_53_11 : STD_LOGIC;
  signal W_reg_53_10 : STD_LOGIC;
  signal W_reg_53_9 : STD_LOGIC;
  signal W_reg_53_8 : STD_LOGIC;
  signal W_reg_53_7 : STD_LOGIC;
  signal W_reg_53_6 : STD_LOGIC;
  signal W_reg_53_5 : STD_LOGIC;
  signal W_reg_53_4 : STD_LOGIC;
  signal W_reg_53_3 : STD_LOGIC;
  signal W_reg_53_2 : STD_LOGIC;
  signal W_reg_53_1 : STD_LOGIC;
  signal W_reg_53_0 : STD_LOGIC;
  signal W_reg_53_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_53_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_53_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_53_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_53_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_53_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_53_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_53_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_53_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_53_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_53_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_53_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_53_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_53_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_53_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_53_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_53_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_53_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_53_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_53_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_53_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_53_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_53_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_53_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_53_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_53_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_53_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_53_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_53_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_53_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_53_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_54_31 : STD_LOGIC;
  signal W_reg_54_30 : STD_LOGIC;
  signal W_reg_54_29 : STD_LOGIC;
  signal W_reg_54_28 : STD_LOGIC;
  signal W_reg_54_27 : STD_LOGIC;
  signal W_reg_54_26 : STD_LOGIC;
  signal W_reg_54_25 : STD_LOGIC;
  signal W_reg_54_24 : STD_LOGIC;
  signal W_reg_54_23 : STD_LOGIC;
  signal W_reg_54_22 : STD_LOGIC;
  signal W_reg_54_21 : STD_LOGIC;
  signal W_reg_54_20 : STD_LOGIC;
  signal W_reg_54_19 : STD_LOGIC;
  signal W_reg_54_18 : STD_LOGIC;
  signal W_reg_54_17 : STD_LOGIC;
  signal W_reg_54_16 : STD_LOGIC;
  signal W_reg_54_15 : STD_LOGIC;
  signal W_reg_54_14 : STD_LOGIC;
  signal W_reg_54_13 : STD_LOGIC;
  signal W_reg_54_12 : STD_LOGIC;
  signal W_reg_54_11 : STD_LOGIC;
  signal W_reg_54_10 : STD_LOGIC;
  signal W_reg_54_9 : STD_LOGIC;
  signal W_reg_54_8 : STD_LOGIC;
  signal W_reg_54_7 : STD_LOGIC;
  signal W_reg_54_6 : STD_LOGIC;
  signal W_reg_54_5 : STD_LOGIC;
  signal W_reg_54_4 : STD_LOGIC;
  signal W_reg_54_3 : STD_LOGIC;
  signal W_reg_54_2 : STD_LOGIC;
  signal W_reg_54_1 : STD_LOGIC;
  signal W_reg_54_0 : STD_LOGIC;
  signal W_reg_54_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_54_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_54_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_54_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_54_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_54_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_54_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_54_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_54_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_54_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_54_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_54_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_54_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_54_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_54_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_54_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_54_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_54_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_54_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_54_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_54_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_54_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_54_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_54_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_54_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_54_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_54_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_54_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_54_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_54_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_54_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_55_31 : STD_LOGIC;
  signal W_reg_55_30 : STD_LOGIC;
  signal W_reg_55_29 : STD_LOGIC;
  signal W_reg_55_28 : STD_LOGIC;
  signal W_reg_55_27 : STD_LOGIC;
  signal W_reg_55_26 : STD_LOGIC;
  signal W_reg_55_25 : STD_LOGIC;
  signal W_reg_55_24 : STD_LOGIC;
  signal W_reg_55_23 : STD_LOGIC;
  signal W_reg_55_22 : STD_LOGIC;
  signal W_reg_55_21 : STD_LOGIC;
  signal W_reg_55_20 : STD_LOGIC;
  signal W_reg_55_19 : STD_LOGIC;
  signal W_reg_55_18 : STD_LOGIC;
  signal W_reg_55_17 : STD_LOGIC;
  signal W_reg_55_16 : STD_LOGIC;
  signal W_reg_55_15 : STD_LOGIC;
  signal W_reg_55_14 : STD_LOGIC;
  signal W_reg_55_13 : STD_LOGIC;
  signal W_reg_55_12 : STD_LOGIC;
  signal W_reg_55_11 : STD_LOGIC;
  signal W_reg_55_10 : STD_LOGIC;
  signal W_reg_55_9 : STD_LOGIC;
  signal W_reg_55_8 : STD_LOGIC;
  signal W_reg_55_7 : STD_LOGIC;
  signal W_reg_55_6 : STD_LOGIC;
  signal W_reg_55_5 : STD_LOGIC;
  signal W_reg_55_4 : STD_LOGIC;
  signal W_reg_55_3 : STD_LOGIC;
  signal W_reg_55_2 : STD_LOGIC;
  signal W_reg_55_1 : STD_LOGIC;
  signal W_reg_55_0 : STD_LOGIC;
  signal W_reg_55_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_55_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_55_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_55_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_55_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_55_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_55_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_55_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_55_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_55_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_55_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_55_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_55_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_55_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_55_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_55_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_55_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_55_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_55_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_55_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_55_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_55_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_55_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_55_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_55_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_55_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_55_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_55_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_55_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_55_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_55_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_56_31 : STD_LOGIC;
  signal W_reg_56_30 : STD_LOGIC;
  signal W_reg_56_29 : STD_LOGIC;
  signal W_reg_56_28 : STD_LOGIC;
  signal W_reg_56_27 : STD_LOGIC;
  signal W_reg_56_26 : STD_LOGIC;
  signal W_reg_56_25 : STD_LOGIC;
  signal W_reg_56_24 : STD_LOGIC;
  signal W_reg_56_23 : STD_LOGIC;
  signal W_reg_56_22 : STD_LOGIC;
  signal W_reg_56_21 : STD_LOGIC;
  signal W_reg_56_20 : STD_LOGIC;
  signal W_reg_56_19 : STD_LOGIC;
  signal W_reg_56_18 : STD_LOGIC;
  signal W_reg_56_17 : STD_LOGIC;
  signal W_reg_56_16 : STD_LOGIC;
  signal W_reg_56_15 : STD_LOGIC;
  signal W_reg_56_14 : STD_LOGIC;
  signal W_reg_56_13 : STD_LOGIC;
  signal W_reg_56_12 : STD_LOGIC;
  signal W_reg_56_11 : STD_LOGIC;
  signal W_reg_56_10 : STD_LOGIC;
  signal W_reg_56_9 : STD_LOGIC;
  signal W_reg_56_8 : STD_LOGIC;
  signal W_reg_56_7 : STD_LOGIC;
  signal W_reg_56_6 : STD_LOGIC;
  signal W_reg_56_5 : STD_LOGIC;
  signal W_reg_56_4 : STD_LOGIC;
  signal W_reg_56_3 : STD_LOGIC;
  signal W_reg_56_2 : STD_LOGIC;
  signal W_reg_56_1 : STD_LOGIC;
  signal W_reg_56_0 : STD_LOGIC;
  signal W_reg_56_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_56_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_56_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_56_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_56_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_56_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_56_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_56_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_56_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_56_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_56_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_56_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_56_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_56_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_56_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_56_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_56_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_56_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_56_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_56_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_56_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_56_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_56_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_56_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_56_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_56_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_56_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_56_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_56_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_56_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_56_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_57_31 : STD_LOGIC;
  signal W_reg_57_30 : STD_LOGIC;
  signal W_reg_57_29 : STD_LOGIC;
  signal W_reg_57_28 : STD_LOGIC;
  signal W_reg_57_27 : STD_LOGIC;
  signal W_reg_57_26 : STD_LOGIC;
  signal W_reg_57_25 : STD_LOGIC;
  signal W_reg_57_24 : STD_LOGIC;
  signal W_reg_57_23 : STD_LOGIC;
  signal W_reg_57_22 : STD_LOGIC;
  signal W_reg_57_21 : STD_LOGIC;
  signal W_reg_57_20 : STD_LOGIC;
  signal W_reg_57_19 : STD_LOGIC;
  signal W_reg_57_18 : STD_LOGIC;
  signal W_reg_57_17 : STD_LOGIC;
  signal W_reg_57_16 : STD_LOGIC;
  signal W_reg_57_15 : STD_LOGIC;
  signal W_reg_57_14 : STD_LOGIC;
  signal W_reg_57_13 : STD_LOGIC;
  signal W_reg_57_12 : STD_LOGIC;
  signal W_reg_57_11 : STD_LOGIC;
  signal W_reg_57_10 : STD_LOGIC;
  signal W_reg_57_9 : STD_LOGIC;
  signal W_reg_57_8 : STD_LOGIC;
  signal W_reg_57_7 : STD_LOGIC;
  signal W_reg_57_6 : STD_LOGIC;
  signal W_reg_57_5 : STD_LOGIC;
  signal W_reg_57_4 : STD_LOGIC;
  signal W_reg_57_3 : STD_LOGIC;
  signal W_reg_57_2 : STD_LOGIC;
  signal W_reg_57_1 : STD_LOGIC;
  signal W_reg_57_0 : STD_LOGIC;
  signal W_reg_57_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_57_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_57_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_57_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_57_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_57_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_57_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_57_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_57_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_57_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_57_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_57_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_57_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_57_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_57_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_57_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_57_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_57_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_57_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_57_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_57_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_57_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_57_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_57_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_57_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_57_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_57_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_57_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_57_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_57_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_57_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_58_31 : STD_LOGIC;
  signal W_reg_58_30 : STD_LOGIC;
  signal W_reg_58_29 : STD_LOGIC;
  signal W_reg_58_28 : STD_LOGIC;
  signal W_reg_58_27 : STD_LOGIC;
  signal W_reg_58_26 : STD_LOGIC;
  signal W_reg_58_25 : STD_LOGIC;
  signal W_reg_58_24 : STD_LOGIC;
  signal W_reg_58_23 : STD_LOGIC;
  signal W_reg_58_22 : STD_LOGIC;
  signal W_reg_58_21 : STD_LOGIC;
  signal W_reg_58_20 : STD_LOGIC;
  signal W_reg_58_19 : STD_LOGIC;
  signal W_reg_58_18 : STD_LOGIC;
  signal W_reg_58_17 : STD_LOGIC;
  signal W_reg_58_16 : STD_LOGIC;
  signal W_reg_58_15 : STD_LOGIC;
  signal W_reg_58_14 : STD_LOGIC;
  signal W_reg_58_13 : STD_LOGIC;
  signal W_reg_58_12 : STD_LOGIC;
  signal W_reg_58_11 : STD_LOGIC;
  signal W_reg_58_10 : STD_LOGIC;
  signal W_reg_58_9 : STD_LOGIC;
  signal W_reg_58_8 : STD_LOGIC;
  signal W_reg_58_7 : STD_LOGIC;
  signal W_reg_58_6 : STD_LOGIC;
  signal W_reg_58_5 : STD_LOGIC;
  signal W_reg_58_4 : STD_LOGIC;
  signal W_reg_58_3 : STD_LOGIC;
  signal W_reg_58_2 : STD_LOGIC;
  signal W_reg_58_1 : STD_LOGIC;
  signal W_reg_58_0 : STD_LOGIC;
  signal W_reg_58_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_58_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_58_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_58_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_58_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_58_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_58_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_58_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_58_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_58_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_58_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_58_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_58_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_58_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_58_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_58_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_58_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_58_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_58_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_58_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_58_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_58_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_58_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_58_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_58_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_58_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_58_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_58_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_58_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_58_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_58_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_59_31 : STD_LOGIC;
  signal W_reg_59_30 : STD_LOGIC;
  signal W_reg_59_29 : STD_LOGIC;
  signal W_reg_59_28 : STD_LOGIC;
  signal W_reg_59_27 : STD_LOGIC;
  signal W_reg_59_26 : STD_LOGIC;
  signal W_reg_59_25 : STD_LOGIC;
  signal W_reg_59_24 : STD_LOGIC;
  signal W_reg_59_23 : STD_LOGIC;
  signal W_reg_59_22 : STD_LOGIC;
  signal W_reg_59_21 : STD_LOGIC;
  signal W_reg_59_20 : STD_LOGIC;
  signal W_reg_59_19 : STD_LOGIC;
  signal W_reg_59_18 : STD_LOGIC;
  signal W_reg_59_17 : STD_LOGIC;
  signal W_reg_59_16 : STD_LOGIC;
  signal W_reg_59_15 : STD_LOGIC;
  signal W_reg_59_14 : STD_LOGIC;
  signal W_reg_59_13 : STD_LOGIC;
  signal W_reg_59_12 : STD_LOGIC;
  signal W_reg_59_11 : STD_LOGIC;
  signal W_reg_59_10 : STD_LOGIC;
  signal W_reg_59_9 : STD_LOGIC;
  signal W_reg_59_8 : STD_LOGIC;
  signal W_reg_59_7 : STD_LOGIC;
  signal W_reg_59_6 : STD_LOGIC;
  signal W_reg_59_5 : STD_LOGIC;
  signal W_reg_59_4 : STD_LOGIC;
  signal W_reg_59_3 : STD_LOGIC;
  signal W_reg_59_2 : STD_LOGIC;
  signal W_reg_59_1 : STD_LOGIC;
  signal W_reg_59_0 : STD_LOGIC;
  signal W_reg_59_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_59_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_59_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_59_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_59_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_59_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_59_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_59_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_59_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_59_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_59_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_59_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_59_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_59_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_59_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_59_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_59_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_59_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_59_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_59_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_59_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_59_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_59_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_59_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_59_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_59_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_59_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_59_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_59_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_59_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_59_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_5_31 : STD_LOGIC;
  signal W_reg_5_30 : STD_LOGIC;
  signal W_reg_5_29 : STD_LOGIC;
  signal W_reg_5_28 : STD_LOGIC;
  signal W_reg_5_27 : STD_LOGIC;
  signal W_reg_5_26 : STD_LOGIC;
  signal W_reg_5_25 : STD_LOGIC;
  signal W_reg_5_24 : STD_LOGIC;
  signal W_reg_5_23 : STD_LOGIC;
  signal W_reg_5_22 : STD_LOGIC;
  signal W_reg_5_21 : STD_LOGIC;
  signal W_reg_5_20 : STD_LOGIC;
  signal W_reg_5_19 : STD_LOGIC;
  signal W_reg_5_18 : STD_LOGIC;
  signal W_reg_5_17 : STD_LOGIC;
  signal W_reg_5_16 : STD_LOGIC;
  signal W_reg_5_15 : STD_LOGIC;
  signal W_reg_5_14 : STD_LOGIC;
  signal W_reg_5_13 : STD_LOGIC;
  signal W_reg_5_12 : STD_LOGIC;
  signal W_reg_5_11 : STD_LOGIC;
  signal W_reg_5_10 : STD_LOGIC;
  signal W_reg_5_9 : STD_LOGIC;
  signal W_reg_5_8 : STD_LOGIC;
  signal W_reg_5_7 : STD_LOGIC;
  signal W_reg_5_6 : STD_LOGIC;
  signal W_reg_5_5 : STD_LOGIC;
  signal W_reg_5_4 : STD_LOGIC;
  signal W_reg_5_3 : STD_LOGIC;
  signal W_reg_5_2 : STD_LOGIC;
  signal W_reg_5_1 : STD_LOGIC;
  signal W_reg_5_0 : STD_LOGIC;
  signal W_reg_60_31 : STD_LOGIC;
  signal W_reg_60_30 : STD_LOGIC;
  signal W_reg_60_29 : STD_LOGIC;
  signal W_reg_60_28 : STD_LOGIC;
  signal W_reg_60_27 : STD_LOGIC;
  signal W_reg_60_26 : STD_LOGIC;
  signal W_reg_60_25 : STD_LOGIC;
  signal W_reg_60_24 : STD_LOGIC;
  signal W_reg_60_23 : STD_LOGIC;
  signal W_reg_60_22 : STD_LOGIC;
  signal W_reg_60_21 : STD_LOGIC;
  signal W_reg_60_20 : STD_LOGIC;
  signal W_reg_60_19 : STD_LOGIC;
  signal W_reg_60_18 : STD_LOGIC;
  signal W_reg_60_17 : STD_LOGIC;
  signal W_reg_60_16 : STD_LOGIC;
  signal W_reg_60_15 : STD_LOGIC;
  signal W_reg_60_14 : STD_LOGIC;
  signal W_reg_60_13 : STD_LOGIC;
  signal W_reg_60_12 : STD_LOGIC;
  signal W_reg_60_11 : STD_LOGIC;
  signal W_reg_60_10 : STD_LOGIC;
  signal W_reg_60_9 : STD_LOGIC;
  signal W_reg_60_8 : STD_LOGIC;
  signal W_reg_60_7 : STD_LOGIC;
  signal W_reg_60_6 : STD_LOGIC;
  signal W_reg_60_5 : STD_LOGIC;
  signal W_reg_60_4 : STD_LOGIC;
  signal W_reg_60_3 : STD_LOGIC;
  signal W_reg_60_2 : STD_LOGIC;
  signal W_reg_60_1 : STD_LOGIC;
  signal W_reg_60_0 : STD_LOGIC;
  signal W_reg_60_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_60_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_60_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_60_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_60_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_60_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_60_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_60_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_60_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_60_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_60_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_60_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_60_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_60_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_60_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_60_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_60_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_60_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_60_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_60_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_60_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_60_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_60_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_60_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_60_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_60_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_60_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_60_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_60_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_60_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_60_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_61_31 : STD_LOGIC;
  signal W_reg_61_30 : STD_LOGIC;
  signal W_reg_61_29 : STD_LOGIC;
  signal W_reg_61_28 : STD_LOGIC;
  signal W_reg_61_27 : STD_LOGIC;
  signal W_reg_61_26 : STD_LOGIC;
  signal W_reg_61_25 : STD_LOGIC;
  signal W_reg_61_24 : STD_LOGIC;
  signal W_reg_61_23 : STD_LOGIC;
  signal W_reg_61_22 : STD_LOGIC;
  signal W_reg_61_21 : STD_LOGIC;
  signal W_reg_61_20 : STD_LOGIC;
  signal W_reg_61_19 : STD_LOGIC;
  signal W_reg_61_18 : STD_LOGIC;
  signal W_reg_61_17 : STD_LOGIC;
  signal W_reg_61_16 : STD_LOGIC;
  signal W_reg_61_15 : STD_LOGIC;
  signal W_reg_61_14 : STD_LOGIC;
  signal W_reg_61_13 : STD_LOGIC;
  signal W_reg_61_12 : STD_LOGIC;
  signal W_reg_61_11 : STD_LOGIC;
  signal W_reg_61_10 : STD_LOGIC;
  signal W_reg_61_9 : STD_LOGIC;
  signal W_reg_61_8 : STD_LOGIC;
  signal W_reg_61_7 : STD_LOGIC;
  signal W_reg_61_6 : STD_LOGIC;
  signal W_reg_61_5 : STD_LOGIC;
  signal W_reg_61_4 : STD_LOGIC;
  signal W_reg_61_3 : STD_LOGIC;
  signal W_reg_61_2 : STD_LOGIC;
  signal W_reg_61_1 : STD_LOGIC;
  signal W_reg_61_0 : STD_LOGIC;
  signal W_reg_61_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_61_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_61_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_61_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_61_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_61_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_61_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_61_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_61_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_61_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_61_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_61_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_61_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_61_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_61_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_61_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_61_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_61_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_61_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_61_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_61_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_61_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_61_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_61_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_61_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_61_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_61_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_61_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_61_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_61_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_61_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_62_31 : STD_LOGIC;
  signal W_reg_62_30 : STD_LOGIC;
  signal W_reg_62_29 : STD_LOGIC;
  signal W_reg_62_28 : STD_LOGIC;
  signal W_reg_62_27 : STD_LOGIC;
  signal W_reg_62_26 : STD_LOGIC;
  signal W_reg_62_25 : STD_LOGIC;
  signal W_reg_62_24 : STD_LOGIC;
  signal W_reg_62_23 : STD_LOGIC;
  signal W_reg_62_22 : STD_LOGIC;
  signal W_reg_62_21 : STD_LOGIC;
  signal W_reg_62_20 : STD_LOGIC;
  signal W_reg_62_19 : STD_LOGIC;
  signal W_reg_62_18 : STD_LOGIC;
  signal W_reg_62_17 : STD_LOGIC;
  signal W_reg_62_16 : STD_LOGIC;
  signal W_reg_62_15 : STD_LOGIC;
  signal W_reg_62_14 : STD_LOGIC;
  signal W_reg_62_13 : STD_LOGIC;
  signal W_reg_62_12 : STD_LOGIC;
  signal W_reg_62_11 : STD_LOGIC;
  signal W_reg_62_10 : STD_LOGIC;
  signal W_reg_62_9 : STD_LOGIC;
  signal W_reg_62_8 : STD_LOGIC;
  signal W_reg_62_7 : STD_LOGIC;
  signal W_reg_62_6 : STD_LOGIC;
  signal W_reg_62_5 : STD_LOGIC;
  signal W_reg_62_4 : STD_LOGIC;
  signal W_reg_62_3 : STD_LOGIC;
  signal W_reg_62_2 : STD_LOGIC;
  signal W_reg_62_1 : STD_LOGIC;
  signal W_reg_62_0 : STD_LOGIC;
  signal W_reg_62_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_62_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_62_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_62_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_62_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_62_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_62_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_62_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_62_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_62_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_62_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_62_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_62_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_62_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_62_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_62_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_62_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_62_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_62_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_62_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_62_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_62_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_62_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_62_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_62_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_62_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_62_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_62_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_62_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_62_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_62_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_63_31 : STD_LOGIC;
  signal W_reg_63_30 : STD_LOGIC;
  signal W_reg_63_29 : STD_LOGIC;
  signal W_reg_63_28 : STD_LOGIC;
  signal W_reg_63_27 : STD_LOGIC;
  signal W_reg_63_26 : STD_LOGIC;
  signal W_reg_63_25 : STD_LOGIC;
  signal W_reg_63_24 : STD_LOGIC;
  signal W_reg_63_23 : STD_LOGIC;
  signal W_reg_63_22 : STD_LOGIC;
  signal W_reg_63_21 : STD_LOGIC;
  signal W_reg_63_20 : STD_LOGIC;
  signal W_reg_63_19 : STD_LOGIC;
  signal W_reg_63_18 : STD_LOGIC;
  signal W_reg_63_17 : STD_LOGIC;
  signal W_reg_63_16 : STD_LOGIC;
  signal W_reg_63_15 : STD_LOGIC;
  signal W_reg_63_14 : STD_LOGIC;
  signal W_reg_63_13 : STD_LOGIC;
  signal W_reg_63_12 : STD_LOGIC;
  signal W_reg_63_11 : STD_LOGIC;
  signal W_reg_63_10 : STD_LOGIC;
  signal W_reg_63_9 : STD_LOGIC;
  signal W_reg_63_8 : STD_LOGIC;
  signal W_reg_63_7 : STD_LOGIC;
  signal W_reg_63_6 : STD_LOGIC;
  signal W_reg_63_5 : STD_LOGIC;
  signal W_reg_63_4 : STD_LOGIC;
  signal W_reg_63_3 : STD_LOGIC;
  signal W_reg_63_2 : STD_LOGIC;
  signal W_reg_63_1 : STD_LOGIC;
  signal W_reg_63_0 : STD_LOGIC;
  signal W_reg_63_11_i_1_n_0 : STD_LOGIC;
  signal W_reg_63_11_i_1_n_1 : STD_LOGIC;
  signal W_reg_63_11_i_1_n_2 : STD_LOGIC;
  signal W_reg_63_11_i_1_n_3 : STD_LOGIC;
  signal W_reg_63_15_i_1_n_0 : STD_LOGIC;
  signal W_reg_63_15_i_1_n_1 : STD_LOGIC;
  signal W_reg_63_15_i_1_n_2 : STD_LOGIC;
  signal W_reg_63_15_i_1_n_3 : STD_LOGIC;
  signal W_reg_63_19_i_1_n_0 : STD_LOGIC;
  signal W_reg_63_19_i_1_n_1 : STD_LOGIC;
  signal W_reg_63_19_i_1_n_2 : STD_LOGIC;
  signal W_reg_63_19_i_1_n_3 : STD_LOGIC;
  signal W_reg_63_23_i_1_n_0 : STD_LOGIC;
  signal W_reg_63_23_i_1_n_1 : STD_LOGIC;
  signal W_reg_63_23_i_1_n_2 : STD_LOGIC;
  signal W_reg_63_23_i_1_n_3 : STD_LOGIC;
  signal W_reg_63_27_i_1_n_0 : STD_LOGIC;
  signal W_reg_63_27_i_1_n_1 : STD_LOGIC;
  signal W_reg_63_27_i_1_n_2 : STD_LOGIC;
  signal W_reg_63_27_i_1_n_3 : STD_LOGIC;
  signal W_reg_63_31_i_1_n_1 : STD_LOGIC;
  signal W_reg_63_31_i_1_n_2 : STD_LOGIC;
  signal W_reg_63_31_i_1_n_3 : STD_LOGIC;
  signal W_reg_63_3_i_1_n_0 : STD_LOGIC;
  signal W_reg_63_3_i_1_n_1 : STD_LOGIC;
  signal W_reg_63_3_i_1_n_2 : STD_LOGIC;
  signal W_reg_63_3_i_1_n_3 : STD_LOGIC;
  signal W_reg_63_7_i_1_n_0 : STD_LOGIC;
  signal W_reg_63_7_i_1_n_1 : STD_LOGIC;
  signal W_reg_63_7_i_1_n_2 : STD_LOGIC;
  signal W_reg_63_7_i_1_n_3 : STD_LOGIC;
  signal W_reg_6_31 : STD_LOGIC;
  signal W_reg_6_30 : STD_LOGIC;
  signal W_reg_6_29 : STD_LOGIC;
  signal W_reg_6_28 : STD_LOGIC;
  signal W_reg_6_27 : STD_LOGIC;
  signal W_reg_6_26 : STD_LOGIC;
  signal W_reg_6_25 : STD_LOGIC;
  signal W_reg_6_24 : STD_LOGIC;
  signal W_reg_6_23 : STD_LOGIC;
  signal W_reg_6_22 : STD_LOGIC;
  signal W_reg_6_21 : STD_LOGIC;
  signal W_reg_6_20 : STD_LOGIC;
  signal W_reg_6_19 : STD_LOGIC;
  signal W_reg_6_18 : STD_LOGIC;
  signal W_reg_6_17 : STD_LOGIC;
  signal W_reg_6_16 : STD_LOGIC;
  signal W_reg_6_15 : STD_LOGIC;
  signal W_reg_6_14 : STD_LOGIC;
  signal W_reg_6_13 : STD_LOGIC;
  signal W_reg_6_12 : STD_LOGIC;
  signal W_reg_6_11 : STD_LOGIC;
  signal W_reg_6_10 : STD_LOGIC;
  signal W_reg_6_9 : STD_LOGIC;
  signal W_reg_6_8 : STD_LOGIC;
  signal W_reg_6_7 : STD_LOGIC;
  signal W_reg_6_6 : STD_LOGIC;
  signal W_reg_6_5 : STD_LOGIC;
  signal W_reg_6_4 : STD_LOGIC;
  signal W_reg_6_3 : STD_LOGIC;
  signal W_reg_6_2 : STD_LOGIC;
  signal W_reg_6_1 : STD_LOGIC;
  signal W_reg_6_0 : STD_LOGIC;
  signal W_reg_7_31 : STD_LOGIC;
  signal W_reg_7_30 : STD_LOGIC;
  signal W_reg_7_29 : STD_LOGIC;
  signal W_reg_7_28 : STD_LOGIC;
  signal W_reg_7_27 : STD_LOGIC;
  signal W_reg_7_26 : STD_LOGIC;
  signal W_reg_7_25 : STD_LOGIC;
  signal W_reg_7_24 : STD_LOGIC;
  signal W_reg_7_23 : STD_LOGIC;
  signal W_reg_7_22 : STD_LOGIC;
  signal W_reg_7_21 : STD_LOGIC;
  signal W_reg_7_20 : STD_LOGIC;
  signal W_reg_7_19 : STD_LOGIC;
  signal W_reg_7_18 : STD_LOGIC;
  signal W_reg_7_17 : STD_LOGIC;
  signal W_reg_7_16 : STD_LOGIC;
  signal W_reg_7_15 : STD_LOGIC;
  signal W_reg_7_14 : STD_LOGIC;
  signal W_reg_7_13 : STD_LOGIC;
  signal W_reg_7_12 : STD_LOGIC;
  signal W_reg_7_11 : STD_LOGIC;
  signal W_reg_7_10 : STD_LOGIC;
  signal W_reg_7_9 : STD_LOGIC;
  signal W_reg_7_8 : STD_LOGIC;
  signal W_reg_7_7 : STD_LOGIC;
  signal W_reg_7_6 : STD_LOGIC;
  signal W_reg_7_5 : STD_LOGIC;
  signal W_reg_7_4 : STD_LOGIC;
  signal W_reg_7_3 : STD_LOGIC;
  signal W_reg_7_2 : STD_LOGIC;
  signal W_reg_7_1 : STD_LOGIC;
  signal W_reg_7_0 : STD_LOGIC;
  signal W_reg_8_31 : STD_LOGIC;
  signal W_reg_8_30 : STD_LOGIC;
  signal W_reg_8_29 : STD_LOGIC;
  signal W_reg_8_28 : STD_LOGIC;
  signal W_reg_8_27 : STD_LOGIC;
  signal W_reg_8_26 : STD_LOGIC;
  signal W_reg_8_25 : STD_LOGIC;
  signal W_reg_8_24 : STD_LOGIC;
  signal W_reg_8_23 : STD_LOGIC;
  signal W_reg_8_22 : STD_LOGIC;
  signal W_reg_8_21 : STD_LOGIC;
  signal W_reg_8_20 : STD_LOGIC;
  signal W_reg_8_19 : STD_LOGIC;
  signal W_reg_8_18 : STD_LOGIC;
  signal W_reg_8_17 : STD_LOGIC;
  signal W_reg_8_16 : STD_LOGIC;
  signal W_reg_8_15 : STD_LOGIC;
  signal W_reg_8_14 : STD_LOGIC;
  signal W_reg_8_13 : STD_LOGIC;
  signal W_reg_8_12 : STD_LOGIC;
  signal W_reg_8_11 : STD_LOGIC;
  signal W_reg_8_10 : STD_LOGIC;
  signal W_reg_8_9 : STD_LOGIC;
  signal W_reg_8_8 : STD_LOGIC;
  signal W_reg_8_7 : STD_LOGIC;
  signal W_reg_8_6 : STD_LOGIC;
  signal W_reg_8_5 : STD_LOGIC;
  signal W_reg_8_4 : STD_LOGIC;
  signal W_reg_8_3 : STD_LOGIC;
  signal W_reg_8_2 : STD_LOGIC;
  signal W_reg_8_1 : STD_LOGIC;
  signal W_reg_8_0 : STD_LOGIC;
  signal W_reg_9_31 : STD_LOGIC;
  signal W_reg_9_30 : STD_LOGIC;
  signal W_reg_9_29 : STD_LOGIC;
  signal W_reg_9_28 : STD_LOGIC;
  signal W_reg_9_27 : STD_LOGIC;
  signal W_reg_9_26 : STD_LOGIC;
  signal W_reg_9_25 : STD_LOGIC;
  signal W_reg_9_24 : STD_LOGIC;
  signal W_reg_9_23 : STD_LOGIC;
  signal W_reg_9_22 : STD_LOGIC;
  signal W_reg_9_21 : STD_LOGIC;
  signal W_reg_9_20 : STD_LOGIC;
  signal W_reg_9_19 : STD_LOGIC;
  signal W_reg_9_18 : STD_LOGIC;
  signal W_reg_9_17 : STD_LOGIC;
  signal W_reg_9_16 : STD_LOGIC;
  signal W_reg_9_15 : STD_LOGIC;
  signal W_reg_9_14 : STD_LOGIC;
  signal W_reg_9_13 : STD_LOGIC;
  signal W_reg_9_12 : STD_LOGIC;
  signal W_reg_9_11 : STD_LOGIC;
  signal W_reg_9_10 : STD_LOGIC;
  signal W_reg_9_9 : STD_LOGIC;
  signal W_reg_9_8 : STD_LOGIC;
  signal W_reg_9_7 : STD_LOGIC;
  signal W_reg_9_6 : STD_LOGIC;
  signal W_reg_9_5 : STD_LOGIC;
  signal W_reg_9_4 : STD_LOGIC;
  signal W_reg_9_3 : STD_LOGIC;
  signal W_reg_9_2 : STD_LOGIC;
  signal W_reg_9_1 : STD_LOGIC;
  signal W_reg_9_0 : STD_LOGIC;
  signal x_31 : STD_LOGIC;
  signal x_30 : STD_LOGIC;
  signal x_29 : STD_LOGIC;
  signal x_28 : STD_LOGIC;
  signal x_27 : STD_LOGIC;
  signal x_26 : STD_LOGIC;
  signal x_25 : STD_LOGIC;
  signal x_24 : STD_LOGIC;
  signal x_23 : STD_LOGIC;
  signal x_22 : STD_LOGIC;
  signal x_21 : STD_LOGIC;
  signal x_20 : STD_LOGIC;
  signal x_19 : STD_LOGIC;
  signal x_18 : STD_LOGIC;
  signal x_17 : STD_LOGIC;
  signal x_16 : STD_LOGIC;
  signal x_15 : STD_LOGIC;
  signal x_14 : STD_LOGIC;
  signal x_13 : STD_LOGIC;
  signal x_12 : STD_LOGIC;
  signal x_11 : STD_LOGIC;
  signal x_10 : STD_LOGIC;
  signal x_9 : STD_LOGIC;
  signal x_8 : STD_LOGIC;
  signal x_7 : STD_LOGIC;
  signal x_6 : STD_LOGIC;
  signal x_5 : STD_LOGIC;
  signal x_4 : STD_LOGIC;
  signal x_3 : STD_LOGIC;
  signal x_2 : STD_LOGIC;
  signal x_1 : STD_LOGIC;
  signal x_0 : STD_LOGIC;
  signal x100_out_31 : STD_LOGIC;
  signal x100_out_30 : STD_LOGIC;
  signal x100_out_29 : STD_LOGIC;
  signal x100_out_28 : STD_LOGIC;
  signal x100_out_27 : STD_LOGIC;
  signal x100_out_26 : STD_LOGIC;
  signal x100_out_25 : STD_LOGIC;
  signal x100_out_24 : STD_LOGIC;
  signal x100_out_23 : STD_LOGIC;
  signal x100_out_22 : STD_LOGIC;
  signal x100_out_21 : STD_LOGIC;
  signal x100_out_20 : STD_LOGIC;
  signal x100_out_19 : STD_LOGIC;
  signal x100_out_18 : STD_LOGIC;
  signal x100_out_17 : STD_LOGIC;
  signal x100_out_16 : STD_LOGIC;
  signal x100_out_15 : STD_LOGIC;
  signal x100_out_14 : STD_LOGIC;
  signal x100_out_13 : STD_LOGIC;
  signal x100_out_12 : STD_LOGIC;
  signal x100_out_11 : STD_LOGIC;
  signal x100_out_10 : STD_LOGIC;
  signal x100_out_9 : STD_LOGIC;
  signal x100_out_8 : STD_LOGIC;
  signal x100_out_7 : STD_LOGIC;
  signal x100_out_6 : STD_LOGIC;
  signal x100_out_5 : STD_LOGIC;
  signal x100_out_4 : STD_LOGIC;
  signal x100_out_3 : STD_LOGIC;
  signal x100_out_2 : STD_LOGIC;
  signal x100_out_1 : STD_LOGIC;
  signal x100_out_0 : STD_LOGIC;
  signal x102_out_31 : STD_LOGIC;
  signal x102_out_30 : STD_LOGIC;
  signal x102_out_29 : STD_LOGIC;
  signal x102_out_28 : STD_LOGIC;
  signal x102_out_27 : STD_LOGIC;
  signal x102_out_26 : STD_LOGIC;
  signal x102_out_25 : STD_LOGIC;
  signal x102_out_24 : STD_LOGIC;
  signal x102_out_23 : STD_LOGIC;
  signal x102_out_22 : STD_LOGIC;
  signal x102_out_21 : STD_LOGIC;
  signal x102_out_20 : STD_LOGIC;
  signal x102_out_19 : STD_LOGIC;
  signal x102_out_18 : STD_LOGIC;
  signal x102_out_17 : STD_LOGIC;
  signal x102_out_16 : STD_LOGIC;
  signal x102_out_15 : STD_LOGIC;
  signal x102_out_14 : STD_LOGIC;
  signal x102_out_13 : STD_LOGIC;
  signal x102_out_12 : STD_LOGIC;
  signal x102_out_11 : STD_LOGIC;
  signal x102_out_10 : STD_LOGIC;
  signal x102_out_9 : STD_LOGIC;
  signal x102_out_8 : STD_LOGIC;
  signal x102_out_7 : STD_LOGIC;
  signal x102_out_6 : STD_LOGIC;
  signal x102_out_5 : STD_LOGIC;
  signal x102_out_4 : STD_LOGIC;
  signal x102_out_3 : STD_LOGIC;
  signal x102_out_2 : STD_LOGIC;
  signal x102_out_1 : STD_LOGIC;
  signal x102_out_0 : STD_LOGIC;
  signal x104_out_31 : STD_LOGIC;
  signal x104_out_30 : STD_LOGIC;
  signal x104_out_29 : STD_LOGIC;
  signal x104_out_28 : STD_LOGIC;
  signal x104_out_27 : STD_LOGIC;
  signal x104_out_26 : STD_LOGIC;
  signal x104_out_25 : STD_LOGIC;
  signal x104_out_24 : STD_LOGIC;
  signal x104_out_23 : STD_LOGIC;
  signal x104_out_22 : STD_LOGIC;
  signal x104_out_21 : STD_LOGIC;
  signal x104_out_20 : STD_LOGIC;
  signal x104_out_19 : STD_LOGIC;
  signal x104_out_18 : STD_LOGIC;
  signal x104_out_17 : STD_LOGIC;
  signal x104_out_16 : STD_LOGIC;
  signal x104_out_15 : STD_LOGIC;
  signal x104_out_14 : STD_LOGIC;
  signal x104_out_13 : STD_LOGIC;
  signal x104_out_12 : STD_LOGIC;
  signal x104_out_11 : STD_LOGIC;
  signal x104_out_10 : STD_LOGIC;
  signal x104_out_9 : STD_LOGIC;
  signal x104_out_8 : STD_LOGIC;
  signal x104_out_7 : STD_LOGIC;
  signal x104_out_6 : STD_LOGIC;
  signal x104_out_5 : STD_LOGIC;
  signal x104_out_4 : STD_LOGIC;
  signal x104_out_3 : STD_LOGIC;
  signal x104_out_2 : STD_LOGIC;
  signal x104_out_1 : STD_LOGIC;
  signal x104_out_0 : STD_LOGIC;
  signal x106_out_31 : STD_LOGIC;
  signal x106_out_30 : STD_LOGIC;
  signal x106_out_29 : STD_LOGIC;
  signal x106_out_28 : STD_LOGIC;
  signal x106_out_27 : STD_LOGIC;
  signal x106_out_26 : STD_LOGIC;
  signal x106_out_25 : STD_LOGIC;
  signal x106_out_24 : STD_LOGIC;
  signal x106_out_23 : STD_LOGIC;
  signal x106_out_22 : STD_LOGIC;
  signal x106_out_21 : STD_LOGIC;
  signal x106_out_20 : STD_LOGIC;
  signal x106_out_19 : STD_LOGIC;
  signal x106_out_18 : STD_LOGIC;
  signal x106_out_17 : STD_LOGIC;
  signal x106_out_16 : STD_LOGIC;
  signal x106_out_15 : STD_LOGIC;
  signal x106_out_14 : STD_LOGIC;
  signal x106_out_13 : STD_LOGIC;
  signal x106_out_12 : STD_LOGIC;
  signal x106_out_11 : STD_LOGIC;
  signal x106_out_10 : STD_LOGIC;
  signal x106_out_9 : STD_LOGIC;
  signal x106_out_8 : STD_LOGIC;
  signal x106_out_7 : STD_LOGIC;
  signal x106_out_6 : STD_LOGIC;
  signal x106_out_5 : STD_LOGIC;
  signal x106_out_4 : STD_LOGIC;
  signal x106_out_3 : STD_LOGIC;
  signal x106_out_2 : STD_LOGIC;
  signal x106_out_1 : STD_LOGIC;
  signal x106_out_0 : STD_LOGIC;
  signal x108_out_31 : STD_LOGIC;
  signal x108_out_30 : STD_LOGIC;
  signal x108_out_29 : STD_LOGIC;
  signal x108_out_28 : STD_LOGIC;
  signal x108_out_27 : STD_LOGIC;
  signal x108_out_26 : STD_LOGIC;
  signal x108_out_25 : STD_LOGIC;
  signal x108_out_24 : STD_LOGIC;
  signal x108_out_23 : STD_LOGIC;
  signal x108_out_22 : STD_LOGIC;
  signal x108_out_21 : STD_LOGIC;
  signal x108_out_20 : STD_LOGIC;
  signal x108_out_19 : STD_LOGIC;
  signal x108_out_18 : STD_LOGIC;
  signal x108_out_17 : STD_LOGIC;
  signal x108_out_16 : STD_LOGIC;
  signal x108_out_15 : STD_LOGIC;
  signal x108_out_14 : STD_LOGIC;
  signal x108_out_13 : STD_LOGIC;
  signal x108_out_12 : STD_LOGIC;
  signal x108_out_11 : STD_LOGIC;
  signal x108_out_10 : STD_LOGIC;
  signal x108_out_9 : STD_LOGIC;
  signal x108_out_8 : STD_LOGIC;
  signal x108_out_7 : STD_LOGIC;
  signal x108_out_6 : STD_LOGIC;
  signal x108_out_5 : STD_LOGIC;
  signal x108_out_4 : STD_LOGIC;
  signal x108_out_3 : STD_LOGIC;
  signal x108_out_2 : STD_LOGIC;
  signal x108_out_1 : STD_LOGIC;
  signal x108_out_0 : STD_LOGIC;
  signal x110_out_31 : STD_LOGIC;
  signal x110_out_30 : STD_LOGIC;
  signal x110_out_29 : STD_LOGIC;
  signal x110_out_28 : STD_LOGIC;
  signal x110_out_27 : STD_LOGIC;
  signal x110_out_26 : STD_LOGIC;
  signal x110_out_25 : STD_LOGIC;
  signal x110_out_24 : STD_LOGIC;
  signal x110_out_23 : STD_LOGIC;
  signal x110_out_22 : STD_LOGIC;
  signal x110_out_21 : STD_LOGIC;
  signal x110_out_20 : STD_LOGIC;
  signal x110_out_19 : STD_LOGIC;
  signal x110_out_18 : STD_LOGIC;
  signal x110_out_17 : STD_LOGIC;
  signal x110_out_16 : STD_LOGIC;
  signal x110_out_15 : STD_LOGIC;
  signal x110_out_14 : STD_LOGIC;
  signal x110_out_13 : STD_LOGIC;
  signal x110_out_12 : STD_LOGIC;
  signal x110_out_11 : STD_LOGIC;
  signal x110_out_10 : STD_LOGIC;
  signal x110_out_9 : STD_LOGIC;
  signal x110_out_8 : STD_LOGIC;
  signal x110_out_7 : STD_LOGIC;
  signal x110_out_6 : STD_LOGIC;
  signal x110_out_5 : STD_LOGIC;
  signal x110_out_4 : STD_LOGIC;
  signal x110_out_3 : STD_LOGIC;
  signal x110_out_2 : STD_LOGIC;
  signal x110_out_1 : STD_LOGIC;
  signal x110_out_0 : STD_LOGIC;
  signal x111_out_31 : STD_LOGIC;
  signal x111_out_30 : STD_LOGIC;
  signal x111_out_29 : STD_LOGIC;
  signal x111_out_28 : STD_LOGIC;
  signal x111_out_27 : STD_LOGIC;
  signal x111_out_26 : STD_LOGIC;
  signal x111_out_25 : STD_LOGIC;
  signal x111_out_24 : STD_LOGIC;
  signal x111_out_23 : STD_LOGIC;
  signal x111_out_22 : STD_LOGIC;
  signal x111_out_21 : STD_LOGIC;
  signal x111_out_20 : STD_LOGIC;
  signal x111_out_19 : STD_LOGIC;
  signal x111_out_18 : STD_LOGIC;
  signal x111_out_17 : STD_LOGIC;
  signal x111_out_16 : STD_LOGIC;
  signal x111_out_15 : STD_LOGIC;
  signal x111_out_14 : STD_LOGIC;
  signal x111_out_13 : STD_LOGIC;
  signal x111_out_12 : STD_LOGIC;
  signal x111_out_11 : STD_LOGIC;
  signal x111_out_10 : STD_LOGIC;
  signal x111_out_9 : STD_LOGIC;
  signal x111_out_8 : STD_LOGIC;
  signal x111_out_7 : STD_LOGIC;
  signal x111_out_6 : STD_LOGIC;
  signal x111_out_5 : STD_LOGIC;
  signal x111_out_4 : STD_LOGIC;
  signal x111_out_3 : STD_LOGIC;
  signal x111_out_2 : STD_LOGIC;
  signal x111_out_1 : STD_LOGIC;
  signal x111_out_0 : STD_LOGIC;
  signal x112_out_31 : STD_LOGIC;
  signal x112_out_30 : STD_LOGIC;
  signal x112_out_29 : STD_LOGIC;
  signal x112_out_28 : STD_LOGIC;
  signal x112_out_27 : STD_LOGIC;
  signal x112_out_26 : STD_LOGIC;
  signal x112_out_25 : STD_LOGIC;
  signal x112_out_24 : STD_LOGIC;
  signal x112_out_23 : STD_LOGIC;
  signal x112_out_22 : STD_LOGIC;
  signal x112_out_21 : STD_LOGIC;
  signal x112_out_20 : STD_LOGIC;
  signal x112_out_19 : STD_LOGIC;
  signal x112_out_18 : STD_LOGIC;
  signal x112_out_17 : STD_LOGIC;
  signal x112_out_16 : STD_LOGIC;
  signal x112_out_15 : STD_LOGIC;
  signal x112_out_14 : STD_LOGIC;
  signal x112_out_13 : STD_LOGIC;
  signal x112_out_12 : STD_LOGIC;
  signal x112_out_11 : STD_LOGIC;
  signal x112_out_10 : STD_LOGIC;
  signal x112_out_9 : STD_LOGIC;
  signal x112_out_8 : STD_LOGIC;
  signal x112_out_7 : STD_LOGIC;
  signal x112_out_6 : STD_LOGIC;
  signal x112_out_5 : STD_LOGIC;
  signal x112_out_4 : STD_LOGIC;
  signal x112_out_3 : STD_LOGIC;
  signal x112_out_2 : STD_LOGIC;
  signal x112_out_1 : STD_LOGIC;
  signal x112_out_0 : STD_LOGIC;
  signal x113_out_31 : STD_LOGIC;
  signal x113_out_30 : STD_LOGIC;
  signal x113_out_29 : STD_LOGIC;
  signal x113_out_28 : STD_LOGIC;
  signal x113_out_27 : STD_LOGIC;
  signal x113_out_26 : STD_LOGIC;
  signal x113_out_25 : STD_LOGIC;
  signal x113_out_24 : STD_LOGIC;
  signal x113_out_23 : STD_LOGIC;
  signal x113_out_22 : STD_LOGIC;
  signal x113_out_21 : STD_LOGIC;
  signal x113_out_20 : STD_LOGIC;
  signal x113_out_19 : STD_LOGIC;
  signal x113_out_18 : STD_LOGIC;
  signal x113_out_17 : STD_LOGIC;
  signal x113_out_16 : STD_LOGIC;
  signal x113_out_15 : STD_LOGIC;
  signal x113_out_14 : STD_LOGIC;
  signal x113_out_13 : STD_LOGIC;
  signal x113_out_12 : STD_LOGIC;
  signal x113_out_11 : STD_LOGIC;
  signal x113_out_10 : STD_LOGIC;
  signal x113_out_9 : STD_LOGIC;
  signal x113_out_8 : STD_LOGIC;
  signal x113_out_7 : STD_LOGIC;
  signal x113_out_6 : STD_LOGIC;
  signal x113_out_5 : STD_LOGIC;
  signal x113_out_4 : STD_LOGIC;
  signal x113_out_3 : STD_LOGIC;
  signal x113_out_2 : STD_LOGIC;
  signal x113_out_1 : STD_LOGIC;
  signal x113_out_0 : STD_LOGIC;
  signal x114_out_31 : STD_LOGIC;
  signal x114_out_30 : STD_LOGIC;
  signal x114_out_29 : STD_LOGIC;
  signal x114_out_28 : STD_LOGIC;
  signal x114_out_27 : STD_LOGIC;
  signal x114_out_26 : STD_LOGIC;
  signal x114_out_25 : STD_LOGIC;
  signal x114_out_24 : STD_LOGIC;
  signal x114_out_23 : STD_LOGIC;
  signal x114_out_22 : STD_LOGIC;
  signal x114_out_21 : STD_LOGIC;
  signal x114_out_20 : STD_LOGIC;
  signal x114_out_19 : STD_LOGIC;
  signal x114_out_18 : STD_LOGIC;
  signal x114_out_17 : STD_LOGIC;
  signal x114_out_16 : STD_LOGIC;
  signal x114_out_15 : STD_LOGIC;
  signal x114_out_14 : STD_LOGIC;
  signal x114_out_13 : STD_LOGIC;
  signal x114_out_12 : STD_LOGIC;
  signal x114_out_11 : STD_LOGIC;
  signal x114_out_10 : STD_LOGIC;
  signal x114_out_9 : STD_LOGIC;
  signal x114_out_8 : STD_LOGIC;
  signal x114_out_7 : STD_LOGIC;
  signal x114_out_6 : STD_LOGIC;
  signal x114_out_5 : STD_LOGIC;
  signal x114_out_4 : STD_LOGIC;
  signal x114_out_3 : STD_LOGIC;
  signal x114_out_2 : STD_LOGIC;
  signal x114_out_1 : STD_LOGIC;
  signal x114_out_0 : STD_LOGIC;
  signal x115_out_31 : STD_LOGIC;
  signal x115_out_30 : STD_LOGIC;
  signal x115_out_29 : STD_LOGIC;
  signal x115_out_28 : STD_LOGIC;
  signal x115_out_27 : STD_LOGIC;
  signal x115_out_26 : STD_LOGIC;
  signal x115_out_25 : STD_LOGIC;
  signal x115_out_24 : STD_LOGIC;
  signal x115_out_23 : STD_LOGIC;
  signal x115_out_22 : STD_LOGIC;
  signal x115_out_21 : STD_LOGIC;
  signal x115_out_20 : STD_LOGIC;
  signal x115_out_19 : STD_LOGIC;
  signal x115_out_18 : STD_LOGIC;
  signal x115_out_17 : STD_LOGIC;
  signal x115_out_16 : STD_LOGIC;
  signal x115_out_15 : STD_LOGIC;
  signal x115_out_14 : STD_LOGIC;
  signal x115_out_13 : STD_LOGIC;
  signal x115_out_12 : STD_LOGIC;
  signal x115_out_11 : STD_LOGIC;
  signal x115_out_10 : STD_LOGIC;
  signal x115_out_9 : STD_LOGIC;
  signal x115_out_8 : STD_LOGIC;
  signal x115_out_7 : STD_LOGIC;
  signal x115_out_6 : STD_LOGIC;
  signal x115_out_5 : STD_LOGIC;
  signal x115_out_4 : STD_LOGIC;
  signal x115_out_3 : STD_LOGIC;
  signal x115_out_2 : STD_LOGIC;
  signal x115_out_1 : STD_LOGIC;
  signal x115_out_0 : STD_LOGIC;
  signal x116_out_31 : STD_LOGIC;
  signal x116_out_30 : STD_LOGIC;
  signal x116_out_29 : STD_LOGIC;
  signal x116_out_28 : STD_LOGIC;
  signal x116_out_27 : STD_LOGIC;
  signal x116_out_26 : STD_LOGIC;
  signal x116_out_25 : STD_LOGIC;
  signal x116_out_24 : STD_LOGIC;
  signal x116_out_23 : STD_LOGIC;
  signal x116_out_22 : STD_LOGIC;
  signal x116_out_21 : STD_LOGIC;
  signal x116_out_20 : STD_LOGIC;
  signal x116_out_19 : STD_LOGIC;
  signal x116_out_18 : STD_LOGIC;
  signal x116_out_17 : STD_LOGIC;
  signal x116_out_16 : STD_LOGIC;
  signal x116_out_15 : STD_LOGIC;
  signal x116_out_14 : STD_LOGIC;
  signal x116_out_13 : STD_LOGIC;
  signal x116_out_12 : STD_LOGIC;
  signal x116_out_11 : STD_LOGIC;
  signal x116_out_10 : STD_LOGIC;
  signal x116_out_9 : STD_LOGIC;
  signal x116_out_8 : STD_LOGIC;
  signal x116_out_7 : STD_LOGIC;
  signal x116_out_6 : STD_LOGIC;
  signal x116_out_5 : STD_LOGIC;
  signal x116_out_4 : STD_LOGIC;
  signal x116_out_3 : STD_LOGIC;
  signal x116_out_2 : STD_LOGIC;
  signal x116_out_1 : STD_LOGIC;
  signal x116_out_0 : STD_LOGIC;
  signal x117_out_31 : STD_LOGIC;
  signal x117_out_30 : STD_LOGIC;
  signal x117_out_29 : STD_LOGIC;
  signal x117_out_28 : STD_LOGIC;
  signal x117_out_27 : STD_LOGIC;
  signal x117_out_26 : STD_LOGIC;
  signal x117_out_25 : STD_LOGIC;
  signal x117_out_24 : STD_LOGIC;
  signal x117_out_23 : STD_LOGIC;
  signal x117_out_22 : STD_LOGIC;
  signal x117_out_21 : STD_LOGIC;
  signal x117_out_20 : STD_LOGIC;
  signal x117_out_19 : STD_LOGIC;
  signal x117_out_18 : STD_LOGIC;
  signal x117_out_17 : STD_LOGIC;
  signal x117_out_16 : STD_LOGIC;
  signal x117_out_15 : STD_LOGIC;
  signal x117_out_14 : STD_LOGIC;
  signal x117_out_13 : STD_LOGIC;
  signal x117_out_12 : STD_LOGIC;
  signal x117_out_11 : STD_LOGIC;
  signal x117_out_10 : STD_LOGIC;
  signal x117_out_9 : STD_LOGIC;
  signal x117_out_8 : STD_LOGIC;
  signal x117_out_7 : STD_LOGIC;
  signal x117_out_6 : STD_LOGIC;
  signal x117_out_5 : STD_LOGIC;
  signal x117_out_4 : STD_LOGIC;
  signal x117_out_3 : STD_LOGIC;
  signal x117_out_2 : STD_LOGIC;
  signal x117_out_1 : STD_LOGIC;
  signal x117_out_0 : STD_LOGIC;
  signal x11_out_31 : STD_LOGIC;
  signal x11_out_30 : STD_LOGIC;
  signal x11_out_29 : STD_LOGIC;
  signal x11_out_28 : STD_LOGIC;
  signal x11_out_27 : STD_LOGIC;
  signal x11_out_26 : STD_LOGIC;
  signal x11_out_25 : STD_LOGIC;
  signal x11_out_24 : STD_LOGIC;
  signal x11_out_23 : STD_LOGIC;
  signal x11_out_22 : STD_LOGIC;
  signal x11_out_21 : STD_LOGIC;
  signal x11_out_20 : STD_LOGIC;
  signal x11_out_19 : STD_LOGIC;
  signal x11_out_18 : STD_LOGIC;
  signal x11_out_17 : STD_LOGIC;
  signal x11_out_16 : STD_LOGIC;
  signal x11_out_15 : STD_LOGIC;
  signal x11_out_14 : STD_LOGIC;
  signal x11_out_13 : STD_LOGIC;
  signal x11_out_12 : STD_LOGIC;
  signal x11_out_11 : STD_LOGIC;
  signal x11_out_10 : STD_LOGIC;
  signal x11_out_9 : STD_LOGIC;
  signal x11_out_8 : STD_LOGIC;
  signal x11_out_7 : STD_LOGIC;
  signal x11_out_6 : STD_LOGIC;
  signal x11_out_5 : STD_LOGIC;
  signal x11_out_4 : STD_LOGIC;
  signal x11_out_3 : STD_LOGIC;
  signal x11_out_2 : STD_LOGIC;
  signal x11_out_1 : STD_LOGIC;
  signal x11_out_0 : STD_LOGIC;
  signal x14_out_31 : STD_LOGIC;
  signal x14_out_30 : STD_LOGIC;
  signal x14_out_29 : STD_LOGIC;
  signal x14_out_28 : STD_LOGIC;
  signal x14_out_27 : STD_LOGIC;
  signal x14_out_26 : STD_LOGIC;
  signal x14_out_25 : STD_LOGIC;
  signal x14_out_24 : STD_LOGIC;
  signal x14_out_23 : STD_LOGIC;
  signal x14_out_22 : STD_LOGIC;
  signal x14_out_21 : STD_LOGIC;
  signal x14_out_20 : STD_LOGIC;
  signal x14_out_19 : STD_LOGIC;
  signal x14_out_18 : STD_LOGIC;
  signal x14_out_17 : STD_LOGIC;
  signal x14_out_16 : STD_LOGIC;
  signal x14_out_15 : STD_LOGIC;
  signal x14_out_14 : STD_LOGIC;
  signal x14_out_13 : STD_LOGIC;
  signal x14_out_12 : STD_LOGIC;
  signal x14_out_11 : STD_LOGIC;
  signal x14_out_10 : STD_LOGIC;
  signal x14_out_9 : STD_LOGIC;
  signal x14_out_8 : STD_LOGIC;
  signal x14_out_7 : STD_LOGIC;
  signal x14_out_6 : STD_LOGIC;
  signal x14_out_5 : STD_LOGIC;
  signal x14_out_4 : STD_LOGIC;
  signal x14_out_3 : STD_LOGIC;
  signal x14_out_2 : STD_LOGIC;
  signal x14_out_1 : STD_LOGIC;
  signal x14_out_0 : STD_LOGIC;
  signal x17_out_31 : STD_LOGIC;
  signal x17_out_30 : STD_LOGIC;
  signal x17_out_29 : STD_LOGIC;
  signal x17_out_28 : STD_LOGIC;
  signal x17_out_27 : STD_LOGIC;
  signal x17_out_26 : STD_LOGIC;
  signal x17_out_25 : STD_LOGIC;
  signal x17_out_24 : STD_LOGIC;
  signal x17_out_23 : STD_LOGIC;
  signal x17_out_22 : STD_LOGIC;
  signal x17_out_21 : STD_LOGIC;
  signal x17_out_20 : STD_LOGIC;
  signal x17_out_19 : STD_LOGIC;
  signal x17_out_18 : STD_LOGIC;
  signal x17_out_17 : STD_LOGIC;
  signal x17_out_16 : STD_LOGIC;
  signal x17_out_15 : STD_LOGIC;
  signal x17_out_14 : STD_LOGIC;
  signal x17_out_13 : STD_LOGIC;
  signal x17_out_12 : STD_LOGIC;
  signal x17_out_11 : STD_LOGIC;
  signal x17_out_10 : STD_LOGIC;
  signal x17_out_9 : STD_LOGIC;
  signal x17_out_8 : STD_LOGIC;
  signal x17_out_7 : STD_LOGIC;
  signal x17_out_6 : STD_LOGIC;
  signal x17_out_5 : STD_LOGIC;
  signal x17_out_4 : STD_LOGIC;
  signal x17_out_3 : STD_LOGIC;
  signal x17_out_2 : STD_LOGIC;
  signal x17_out_1 : STD_LOGIC;
  signal x17_out_0 : STD_LOGIC;
  signal x20_out_31 : STD_LOGIC;
  signal x20_out_30 : STD_LOGIC;
  signal x20_out_29 : STD_LOGIC;
  signal x20_out_28 : STD_LOGIC;
  signal x20_out_27 : STD_LOGIC;
  signal x20_out_26 : STD_LOGIC;
  signal x20_out_25 : STD_LOGIC;
  signal x20_out_24 : STD_LOGIC;
  signal x20_out_23 : STD_LOGIC;
  signal x20_out_22 : STD_LOGIC;
  signal x20_out_21 : STD_LOGIC;
  signal x20_out_20 : STD_LOGIC;
  signal x20_out_19 : STD_LOGIC;
  signal x20_out_18 : STD_LOGIC;
  signal x20_out_17 : STD_LOGIC;
  signal x20_out_16 : STD_LOGIC;
  signal x20_out_15 : STD_LOGIC;
  signal x20_out_14 : STD_LOGIC;
  signal x20_out_13 : STD_LOGIC;
  signal x20_out_12 : STD_LOGIC;
  signal x20_out_11 : STD_LOGIC;
  signal x20_out_10 : STD_LOGIC;
  signal x20_out_9 : STD_LOGIC;
  signal x20_out_8 : STD_LOGIC;
  signal x20_out_7 : STD_LOGIC;
  signal x20_out_6 : STD_LOGIC;
  signal x20_out_5 : STD_LOGIC;
  signal x20_out_4 : STD_LOGIC;
  signal x20_out_3 : STD_LOGIC;
  signal x20_out_2 : STD_LOGIC;
  signal x20_out_1 : STD_LOGIC;
  signal x20_out_0 : STD_LOGIC;
  signal x23_out_31 : STD_LOGIC;
  signal x23_out_30 : STD_LOGIC;
  signal x23_out_29 : STD_LOGIC;
  signal x23_out_28 : STD_LOGIC;
  signal x23_out_27 : STD_LOGIC;
  signal x23_out_26 : STD_LOGIC;
  signal x23_out_25 : STD_LOGIC;
  signal x23_out_24 : STD_LOGIC;
  signal x23_out_23 : STD_LOGIC;
  signal x23_out_22 : STD_LOGIC;
  signal x23_out_21 : STD_LOGIC;
  signal x23_out_20 : STD_LOGIC;
  signal x23_out_19 : STD_LOGIC;
  signal x23_out_18 : STD_LOGIC;
  signal x23_out_17 : STD_LOGIC;
  signal x23_out_16 : STD_LOGIC;
  signal x23_out_15 : STD_LOGIC;
  signal x23_out_14 : STD_LOGIC;
  signal x23_out_13 : STD_LOGIC;
  signal x23_out_12 : STD_LOGIC;
  signal x23_out_11 : STD_LOGIC;
  signal x23_out_10 : STD_LOGIC;
  signal x23_out_9 : STD_LOGIC;
  signal x23_out_8 : STD_LOGIC;
  signal x23_out_7 : STD_LOGIC;
  signal x23_out_6 : STD_LOGIC;
  signal x23_out_5 : STD_LOGIC;
  signal x23_out_4 : STD_LOGIC;
  signal x23_out_3 : STD_LOGIC;
  signal x23_out_2 : STD_LOGIC;
  signal x23_out_1 : STD_LOGIC;
  signal x23_out_0 : STD_LOGIC;
  signal x26_out_31 : STD_LOGIC;
  signal x26_out_30 : STD_LOGIC;
  signal x26_out_29 : STD_LOGIC;
  signal x26_out_28 : STD_LOGIC;
  signal x26_out_27 : STD_LOGIC;
  signal x26_out_26 : STD_LOGIC;
  signal x26_out_25 : STD_LOGIC;
  signal x26_out_24 : STD_LOGIC;
  signal x26_out_23 : STD_LOGIC;
  signal x26_out_22 : STD_LOGIC;
  signal x26_out_21 : STD_LOGIC;
  signal x26_out_20 : STD_LOGIC;
  signal x26_out_19 : STD_LOGIC;
  signal x26_out_18 : STD_LOGIC;
  signal x26_out_17 : STD_LOGIC;
  signal x26_out_16 : STD_LOGIC;
  signal x26_out_15 : STD_LOGIC;
  signal x26_out_14 : STD_LOGIC;
  signal x26_out_13 : STD_LOGIC;
  signal x26_out_12 : STD_LOGIC;
  signal x26_out_11 : STD_LOGIC;
  signal x26_out_10 : STD_LOGIC;
  signal x26_out_9 : STD_LOGIC;
  signal x26_out_8 : STD_LOGIC;
  signal x26_out_7 : STD_LOGIC;
  signal x26_out_6 : STD_LOGIC;
  signal x26_out_5 : STD_LOGIC;
  signal x26_out_4 : STD_LOGIC;
  signal x26_out_3 : STD_LOGIC;
  signal x26_out_2 : STD_LOGIC;
  signal x26_out_1 : STD_LOGIC;
  signal x26_out_0 : STD_LOGIC;
  signal x29_out_31 : STD_LOGIC;
  signal x29_out_30 : STD_LOGIC;
  signal x29_out_29 : STD_LOGIC;
  signal x29_out_28 : STD_LOGIC;
  signal x29_out_27 : STD_LOGIC;
  signal x29_out_26 : STD_LOGIC;
  signal x29_out_25 : STD_LOGIC;
  signal x29_out_24 : STD_LOGIC;
  signal x29_out_23 : STD_LOGIC;
  signal x29_out_22 : STD_LOGIC;
  signal x29_out_21 : STD_LOGIC;
  signal x29_out_20 : STD_LOGIC;
  signal x29_out_19 : STD_LOGIC;
  signal x29_out_18 : STD_LOGIC;
  signal x29_out_17 : STD_LOGIC;
  signal x29_out_16 : STD_LOGIC;
  signal x29_out_15 : STD_LOGIC;
  signal x29_out_14 : STD_LOGIC;
  signal x29_out_13 : STD_LOGIC;
  signal x29_out_12 : STD_LOGIC;
  signal x29_out_11 : STD_LOGIC;
  signal x29_out_10 : STD_LOGIC;
  signal x29_out_9 : STD_LOGIC;
  signal x29_out_8 : STD_LOGIC;
  signal x29_out_7 : STD_LOGIC;
  signal x29_out_6 : STD_LOGIC;
  signal x29_out_5 : STD_LOGIC;
  signal x29_out_4 : STD_LOGIC;
  signal x29_out_3 : STD_LOGIC;
  signal x29_out_2 : STD_LOGIC;
  signal x29_out_1 : STD_LOGIC;
  signal x29_out_0 : STD_LOGIC;
  signal x32_out_31 : STD_LOGIC;
  signal x32_out_30 : STD_LOGIC;
  signal x32_out_29 : STD_LOGIC;
  signal x32_out_28 : STD_LOGIC;
  signal x32_out_27 : STD_LOGIC;
  signal x32_out_26 : STD_LOGIC;
  signal x32_out_25 : STD_LOGIC;
  signal x32_out_24 : STD_LOGIC;
  signal x32_out_23 : STD_LOGIC;
  signal x32_out_22 : STD_LOGIC;
  signal x32_out_21 : STD_LOGIC;
  signal x32_out_20 : STD_LOGIC;
  signal x32_out_19 : STD_LOGIC;
  signal x32_out_18 : STD_LOGIC;
  signal x32_out_17 : STD_LOGIC;
  signal x32_out_16 : STD_LOGIC;
  signal x32_out_15 : STD_LOGIC;
  signal x32_out_14 : STD_LOGIC;
  signal x32_out_13 : STD_LOGIC;
  signal x32_out_12 : STD_LOGIC;
  signal x32_out_11 : STD_LOGIC;
  signal x32_out_10 : STD_LOGIC;
  signal x32_out_9 : STD_LOGIC;
  signal x32_out_8 : STD_LOGIC;
  signal x32_out_7 : STD_LOGIC;
  signal x32_out_6 : STD_LOGIC;
  signal x32_out_5 : STD_LOGIC;
  signal x32_out_4 : STD_LOGIC;
  signal x32_out_3 : STD_LOGIC;
  signal x32_out_2 : STD_LOGIC;
  signal x32_out_1 : STD_LOGIC;
  signal x32_out_0 : STD_LOGIC;
  signal x35_out_31 : STD_LOGIC;
  signal x35_out_30 : STD_LOGIC;
  signal x35_out_29 : STD_LOGIC;
  signal x35_out_28 : STD_LOGIC;
  signal x35_out_27 : STD_LOGIC;
  signal x35_out_26 : STD_LOGIC;
  signal x35_out_25 : STD_LOGIC;
  signal x35_out_24 : STD_LOGIC;
  signal x35_out_23 : STD_LOGIC;
  signal x35_out_22 : STD_LOGIC;
  signal x35_out_21 : STD_LOGIC;
  signal x35_out_20 : STD_LOGIC;
  signal x35_out_19 : STD_LOGIC;
  signal x35_out_18 : STD_LOGIC;
  signal x35_out_17 : STD_LOGIC;
  signal x35_out_16 : STD_LOGIC;
  signal x35_out_15 : STD_LOGIC;
  signal x35_out_14 : STD_LOGIC;
  signal x35_out_13 : STD_LOGIC;
  signal x35_out_12 : STD_LOGIC;
  signal x35_out_11 : STD_LOGIC;
  signal x35_out_10 : STD_LOGIC;
  signal x35_out_9 : STD_LOGIC;
  signal x35_out_8 : STD_LOGIC;
  signal x35_out_7 : STD_LOGIC;
  signal x35_out_6 : STD_LOGIC;
  signal x35_out_5 : STD_LOGIC;
  signal x35_out_4 : STD_LOGIC;
  signal x35_out_3 : STD_LOGIC;
  signal x35_out_2 : STD_LOGIC;
  signal x35_out_1 : STD_LOGIC;
  signal x35_out_0 : STD_LOGIC;
  signal x38_out_31 : STD_LOGIC;
  signal x38_out_30 : STD_LOGIC;
  signal x38_out_29 : STD_LOGIC;
  signal x38_out_28 : STD_LOGIC;
  signal x38_out_27 : STD_LOGIC;
  signal x38_out_26 : STD_LOGIC;
  signal x38_out_25 : STD_LOGIC;
  signal x38_out_24 : STD_LOGIC;
  signal x38_out_23 : STD_LOGIC;
  signal x38_out_22 : STD_LOGIC;
  signal x38_out_21 : STD_LOGIC;
  signal x38_out_20 : STD_LOGIC;
  signal x38_out_19 : STD_LOGIC;
  signal x38_out_18 : STD_LOGIC;
  signal x38_out_17 : STD_LOGIC;
  signal x38_out_16 : STD_LOGIC;
  signal x38_out_15 : STD_LOGIC;
  signal x38_out_14 : STD_LOGIC;
  signal x38_out_13 : STD_LOGIC;
  signal x38_out_12 : STD_LOGIC;
  signal x38_out_11 : STD_LOGIC;
  signal x38_out_10 : STD_LOGIC;
  signal x38_out_9 : STD_LOGIC;
  signal x38_out_8 : STD_LOGIC;
  signal x38_out_7 : STD_LOGIC;
  signal x38_out_6 : STD_LOGIC;
  signal x38_out_5 : STD_LOGIC;
  signal x38_out_4 : STD_LOGIC;
  signal x38_out_3 : STD_LOGIC;
  signal x38_out_2 : STD_LOGIC;
  signal x38_out_1 : STD_LOGIC;
  signal x38_out_0 : STD_LOGIC;
  signal x41_out_31 : STD_LOGIC;
  signal x41_out_30 : STD_LOGIC;
  signal x41_out_29 : STD_LOGIC;
  signal x41_out_28 : STD_LOGIC;
  signal x41_out_27 : STD_LOGIC;
  signal x41_out_26 : STD_LOGIC;
  signal x41_out_25 : STD_LOGIC;
  signal x41_out_24 : STD_LOGIC;
  signal x41_out_23 : STD_LOGIC;
  signal x41_out_22 : STD_LOGIC;
  signal x41_out_21 : STD_LOGIC;
  signal x41_out_20 : STD_LOGIC;
  signal x41_out_19 : STD_LOGIC;
  signal x41_out_18 : STD_LOGIC;
  signal x41_out_17 : STD_LOGIC;
  signal x41_out_16 : STD_LOGIC;
  signal x41_out_15 : STD_LOGIC;
  signal x41_out_14 : STD_LOGIC;
  signal x41_out_13 : STD_LOGIC;
  signal x41_out_12 : STD_LOGIC;
  signal x41_out_11 : STD_LOGIC;
  signal x41_out_10 : STD_LOGIC;
  signal x41_out_9 : STD_LOGIC;
  signal x41_out_8 : STD_LOGIC;
  signal x41_out_7 : STD_LOGIC;
  signal x41_out_6 : STD_LOGIC;
  signal x41_out_5 : STD_LOGIC;
  signal x41_out_4 : STD_LOGIC;
  signal x41_out_3 : STD_LOGIC;
  signal x41_out_2 : STD_LOGIC;
  signal x41_out_1 : STD_LOGIC;
  signal x41_out_0 : STD_LOGIC;
  signal x44_out_31 : STD_LOGIC;
  signal x44_out_30 : STD_LOGIC;
  signal x44_out_29 : STD_LOGIC;
  signal x44_out_28 : STD_LOGIC;
  signal x44_out_27 : STD_LOGIC;
  signal x44_out_26 : STD_LOGIC;
  signal x44_out_25 : STD_LOGIC;
  signal x44_out_24 : STD_LOGIC;
  signal x44_out_23 : STD_LOGIC;
  signal x44_out_22 : STD_LOGIC;
  signal x44_out_21 : STD_LOGIC;
  signal x44_out_20 : STD_LOGIC;
  signal x44_out_19 : STD_LOGIC;
  signal x44_out_18 : STD_LOGIC;
  signal x44_out_17 : STD_LOGIC;
  signal x44_out_16 : STD_LOGIC;
  signal x44_out_15 : STD_LOGIC;
  signal x44_out_14 : STD_LOGIC;
  signal x44_out_13 : STD_LOGIC;
  signal x44_out_12 : STD_LOGIC;
  signal x44_out_11 : STD_LOGIC;
  signal x44_out_10 : STD_LOGIC;
  signal x44_out_9 : STD_LOGIC;
  signal x44_out_8 : STD_LOGIC;
  signal x44_out_7 : STD_LOGIC;
  signal x44_out_6 : STD_LOGIC;
  signal x44_out_5 : STD_LOGIC;
  signal x44_out_4 : STD_LOGIC;
  signal x44_out_3 : STD_LOGIC;
  signal x44_out_2 : STD_LOGIC;
  signal x44_out_1 : STD_LOGIC;
  signal x44_out_0 : STD_LOGIC;
  signal x47_out_31 : STD_LOGIC;
  signal x47_out_30 : STD_LOGIC;
  signal x47_out_29 : STD_LOGIC;
  signal x47_out_28 : STD_LOGIC;
  signal x47_out_27 : STD_LOGIC;
  signal x47_out_26 : STD_LOGIC;
  signal x47_out_25 : STD_LOGIC;
  signal x47_out_24 : STD_LOGIC;
  signal x47_out_23 : STD_LOGIC;
  signal x47_out_22 : STD_LOGIC;
  signal x47_out_21 : STD_LOGIC;
  signal x47_out_20 : STD_LOGIC;
  signal x47_out_19 : STD_LOGIC;
  signal x47_out_18 : STD_LOGIC;
  signal x47_out_17 : STD_LOGIC;
  signal x47_out_16 : STD_LOGIC;
  signal x47_out_15 : STD_LOGIC;
  signal x47_out_14 : STD_LOGIC;
  signal x47_out_13 : STD_LOGIC;
  signal x47_out_12 : STD_LOGIC;
  signal x47_out_11 : STD_LOGIC;
  signal x47_out_10 : STD_LOGIC;
  signal x47_out_9 : STD_LOGIC;
  signal x47_out_8 : STD_LOGIC;
  signal x47_out_7 : STD_LOGIC;
  signal x47_out_6 : STD_LOGIC;
  signal x47_out_5 : STD_LOGIC;
  signal x47_out_4 : STD_LOGIC;
  signal x47_out_3 : STD_LOGIC;
  signal x47_out_2 : STD_LOGIC;
  signal x47_out_1 : STD_LOGIC;
  signal x47_out_0 : STD_LOGIC;
  signal x50_out_31 : STD_LOGIC;
  signal x50_out_30 : STD_LOGIC;
  signal x50_out_29 : STD_LOGIC;
  signal x50_out_28 : STD_LOGIC;
  signal x50_out_27 : STD_LOGIC;
  signal x50_out_26 : STD_LOGIC;
  signal x50_out_25 : STD_LOGIC;
  signal x50_out_24 : STD_LOGIC;
  signal x50_out_23 : STD_LOGIC;
  signal x50_out_22 : STD_LOGIC;
  signal x50_out_21 : STD_LOGIC;
  signal x50_out_20 : STD_LOGIC;
  signal x50_out_19 : STD_LOGIC;
  signal x50_out_18 : STD_LOGIC;
  signal x50_out_17 : STD_LOGIC;
  signal x50_out_16 : STD_LOGIC;
  signal x50_out_15 : STD_LOGIC;
  signal x50_out_14 : STD_LOGIC;
  signal x50_out_13 : STD_LOGIC;
  signal x50_out_12 : STD_LOGIC;
  signal x50_out_11 : STD_LOGIC;
  signal x50_out_10 : STD_LOGIC;
  signal x50_out_9 : STD_LOGIC;
  signal x50_out_8 : STD_LOGIC;
  signal x50_out_7 : STD_LOGIC;
  signal x50_out_6 : STD_LOGIC;
  signal x50_out_5 : STD_LOGIC;
  signal x50_out_4 : STD_LOGIC;
  signal x50_out_3 : STD_LOGIC;
  signal x50_out_2 : STD_LOGIC;
  signal x50_out_1 : STD_LOGIC;
  signal x50_out_0 : STD_LOGIC;
  signal x53_out_31 : STD_LOGIC;
  signal x53_out_30 : STD_LOGIC;
  signal x53_out_29 : STD_LOGIC;
  signal x53_out_28 : STD_LOGIC;
  signal x53_out_27 : STD_LOGIC;
  signal x53_out_26 : STD_LOGIC;
  signal x53_out_25 : STD_LOGIC;
  signal x53_out_24 : STD_LOGIC;
  signal x53_out_23 : STD_LOGIC;
  signal x53_out_22 : STD_LOGIC;
  signal x53_out_21 : STD_LOGIC;
  signal x53_out_20 : STD_LOGIC;
  signal x53_out_19 : STD_LOGIC;
  signal x53_out_18 : STD_LOGIC;
  signal x53_out_17 : STD_LOGIC;
  signal x53_out_16 : STD_LOGIC;
  signal x53_out_15 : STD_LOGIC;
  signal x53_out_14 : STD_LOGIC;
  signal x53_out_13 : STD_LOGIC;
  signal x53_out_12 : STD_LOGIC;
  signal x53_out_11 : STD_LOGIC;
  signal x53_out_10 : STD_LOGIC;
  signal x53_out_9 : STD_LOGIC;
  signal x53_out_8 : STD_LOGIC;
  signal x53_out_7 : STD_LOGIC;
  signal x53_out_6 : STD_LOGIC;
  signal x53_out_5 : STD_LOGIC;
  signal x53_out_4 : STD_LOGIC;
  signal x53_out_3 : STD_LOGIC;
  signal x53_out_2 : STD_LOGIC;
  signal x53_out_1 : STD_LOGIC;
  signal x53_out_0 : STD_LOGIC;
  signal x56_out_31 : STD_LOGIC;
  signal x56_out_30 : STD_LOGIC;
  signal x56_out_29 : STD_LOGIC;
  signal x56_out_28 : STD_LOGIC;
  signal x56_out_27 : STD_LOGIC;
  signal x56_out_26 : STD_LOGIC;
  signal x56_out_25 : STD_LOGIC;
  signal x56_out_24 : STD_LOGIC;
  signal x56_out_23 : STD_LOGIC;
  signal x56_out_22 : STD_LOGIC;
  signal x56_out_21 : STD_LOGIC;
  signal x56_out_20 : STD_LOGIC;
  signal x56_out_19 : STD_LOGIC;
  signal x56_out_18 : STD_LOGIC;
  signal x56_out_17 : STD_LOGIC;
  signal x56_out_16 : STD_LOGIC;
  signal x56_out_15 : STD_LOGIC;
  signal x56_out_14 : STD_LOGIC;
  signal x56_out_13 : STD_LOGIC;
  signal x56_out_12 : STD_LOGIC;
  signal x56_out_11 : STD_LOGIC;
  signal x56_out_10 : STD_LOGIC;
  signal x56_out_9 : STD_LOGIC;
  signal x56_out_8 : STD_LOGIC;
  signal x56_out_7 : STD_LOGIC;
  signal x56_out_6 : STD_LOGIC;
  signal x56_out_5 : STD_LOGIC;
  signal x56_out_4 : STD_LOGIC;
  signal x56_out_3 : STD_LOGIC;
  signal x56_out_2 : STD_LOGIC;
  signal x56_out_1 : STD_LOGIC;
  signal x56_out_0 : STD_LOGIC;
  signal x59_out_31 : STD_LOGIC;
  signal x59_out_30 : STD_LOGIC;
  signal x59_out_29 : STD_LOGIC;
  signal x59_out_28 : STD_LOGIC;
  signal x59_out_27 : STD_LOGIC;
  signal x59_out_26 : STD_LOGIC;
  signal x59_out_25 : STD_LOGIC;
  signal x59_out_24 : STD_LOGIC;
  signal x59_out_23 : STD_LOGIC;
  signal x59_out_22 : STD_LOGIC;
  signal x59_out_21 : STD_LOGIC;
  signal x59_out_20 : STD_LOGIC;
  signal x59_out_19 : STD_LOGIC;
  signal x59_out_18 : STD_LOGIC;
  signal x59_out_17 : STD_LOGIC;
  signal x59_out_16 : STD_LOGIC;
  signal x59_out_15 : STD_LOGIC;
  signal x59_out_14 : STD_LOGIC;
  signal x59_out_13 : STD_LOGIC;
  signal x59_out_12 : STD_LOGIC;
  signal x59_out_11 : STD_LOGIC;
  signal x59_out_10 : STD_LOGIC;
  signal x59_out_9 : STD_LOGIC;
  signal x59_out_8 : STD_LOGIC;
  signal x59_out_7 : STD_LOGIC;
  signal x59_out_6 : STD_LOGIC;
  signal x59_out_5 : STD_LOGIC;
  signal x59_out_4 : STD_LOGIC;
  signal x59_out_3 : STD_LOGIC;
  signal x59_out_2 : STD_LOGIC;
  signal x59_out_1 : STD_LOGIC;
  signal x59_out_0 : STD_LOGIC;
  signal x62_out_31 : STD_LOGIC;
  signal x62_out_30 : STD_LOGIC;
  signal x62_out_29 : STD_LOGIC;
  signal x62_out_28 : STD_LOGIC;
  signal x62_out_27 : STD_LOGIC;
  signal x62_out_26 : STD_LOGIC;
  signal x62_out_25 : STD_LOGIC;
  signal x62_out_24 : STD_LOGIC;
  signal x62_out_23 : STD_LOGIC;
  signal x62_out_22 : STD_LOGIC;
  signal x62_out_21 : STD_LOGIC;
  signal x62_out_20 : STD_LOGIC;
  signal x62_out_19 : STD_LOGIC;
  signal x62_out_18 : STD_LOGIC;
  signal x62_out_17 : STD_LOGIC;
  signal x62_out_16 : STD_LOGIC;
  signal x62_out_15 : STD_LOGIC;
  signal x62_out_14 : STD_LOGIC;
  signal x62_out_13 : STD_LOGIC;
  signal x62_out_12 : STD_LOGIC;
  signal x62_out_11 : STD_LOGIC;
  signal x62_out_10 : STD_LOGIC;
  signal x62_out_9 : STD_LOGIC;
  signal x62_out_8 : STD_LOGIC;
  signal x62_out_7 : STD_LOGIC;
  signal x62_out_6 : STD_LOGIC;
  signal x62_out_5 : STD_LOGIC;
  signal x62_out_4 : STD_LOGIC;
  signal x62_out_3 : STD_LOGIC;
  signal x62_out_2 : STD_LOGIC;
  signal x62_out_1 : STD_LOGIC;
  signal x62_out_0 : STD_LOGIC;
  signal x65_out_31 : STD_LOGIC;
  signal x65_out_30 : STD_LOGIC;
  signal x65_out_29 : STD_LOGIC;
  signal x65_out_28 : STD_LOGIC;
  signal x65_out_27 : STD_LOGIC;
  signal x65_out_26 : STD_LOGIC;
  signal x65_out_25 : STD_LOGIC;
  signal x65_out_24 : STD_LOGIC;
  signal x65_out_23 : STD_LOGIC;
  signal x65_out_22 : STD_LOGIC;
  signal x65_out_21 : STD_LOGIC;
  signal x65_out_20 : STD_LOGIC;
  signal x65_out_19 : STD_LOGIC;
  signal x65_out_18 : STD_LOGIC;
  signal x65_out_17 : STD_LOGIC;
  signal x65_out_16 : STD_LOGIC;
  signal x65_out_15 : STD_LOGIC;
  signal x65_out_14 : STD_LOGIC;
  signal x65_out_13 : STD_LOGIC;
  signal x65_out_12 : STD_LOGIC;
  signal x65_out_11 : STD_LOGIC;
  signal x65_out_10 : STD_LOGIC;
  signal x65_out_9 : STD_LOGIC;
  signal x65_out_8 : STD_LOGIC;
  signal x65_out_7 : STD_LOGIC;
  signal x65_out_6 : STD_LOGIC;
  signal x65_out_5 : STD_LOGIC;
  signal x65_out_4 : STD_LOGIC;
  signal x65_out_3 : STD_LOGIC;
  signal x65_out_2 : STD_LOGIC;
  signal x65_out_1 : STD_LOGIC;
  signal x65_out_0 : STD_LOGIC;
  signal x68_out_31 : STD_LOGIC;
  signal x68_out_30 : STD_LOGIC;
  signal x68_out_29 : STD_LOGIC;
  signal x68_out_28 : STD_LOGIC;
  signal x68_out_27 : STD_LOGIC;
  signal x68_out_26 : STD_LOGIC;
  signal x68_out_25 : STD_LOGIC;
  signal x68_out_24 : STD_LOGIC;
  signal x68_out_23 : STD_LOGIC;
  signal x68_out_22 : STD_LOGIC;
  signal x68_out_21 : STD_LOGIC;
  signal x68_out_20 : STD_LOGIC;
  signal x68_out_19 : STD_LOGIC;
  signal x68_out_18 : STD_LOGIC;
  signal x68_out_17 : STD_LOGIC;
  signal x68_out_16 : STD_LOGIC;
  signal x68_out_15 : STD_LOGIC;
  signal x68_out_14 : STD_LOGIC;
  signal x68_out_13 : STD_LOGIC;
  signal x68_out_12 : STD_LOGIC;
  signal x68_out_11 : STD_LOGIC;
  signal x68_out_10 : STD_LOGIC;
  signal x68_out_9 : STD_LOGIC;
  signal x68_out_8 : STD_LOGIC;
  signal x68_out_7 : STD_LOGIC;
  signal x68_out_6 : STD_LOGIC;
  signal x68_out_5 : STD_LOGIC;
  signal x68_out_4 : STD_LOGIC;
  signal x68_out_3 : STD_LOGIC;
  signal x68_out_2 : STD_LOGIC;
  signal x68_out_1 : STD_LOGIC;
  signal x68_out_0 : STD_LOGIC;
  signal x71_out_31 : STD_LOGIC;
  signal x71_out_30 : STD_LOGIC;
  signal x71_out_29 : STD_LOGIC;
  signal x71_out_28 : STD_LOGIC;
  signal x71_out_27 : STD_LOGIC;
  signal x71_out_26 : STD_LOGIC;
  signal x71_out_25 : STD_LOGIC;
  signal x71_out_24 : STD_LOGIC;
  signal x71_out_23 : STD_LOGIC;
  signal x71_out_22 : STD_LOGIC;
  signal x71_out_21 : STD_LOGIC;
  signal x71_out_20 : STD_LOGIC;
  signal x71_out_19 : STD_LOGIC;
  signal x71_out_18 : STD_LOGIC;
  signal x71_out_17 : STD_LOGIC;
  signal x71_out_16 : STD_LOGIC;
  signal x71_out_15 : STD_LOGIC;
  signal x71_out_14 : STD_LOGIC;
  signal x71_out_13 : STD_LOGIC;
  signal x71_out_12 : STD_LOGIC;
  signal x71_out_11 : STD_LOGIC;
  signal x71_out_10 : STD_LOGIC;
  signal x71_out_9 : STD_LOGIC;
  signal x71_out_8 : STD_LOGIC;
  signal x71_out_7 : STD_LOGIC;
  signal x71_out_6 : STD_LOGIC;
  signal x71_out_5 : STD_LOGIC;
  signal x71_out_4 : STD_LOGIC;
  signal x71_out_3 : STD_LOGIC;
  signal x71_out_2 : STD_LOGIC;
  signal x71_out_1 : STD_LOGIC;
  signal x71_out_0 : STD_LOGIC;
  signal x74_out_31 : STD_LOGIC;
  signal x74_out_30 : STD_LOGIC;
  signal x74_out_29 : STD_LOGIC;
  signal x74_out_28 : STD_LOGIC;
  signal x74_out_27 : STD_LOGIC;
  signal x74_out_26 : STD_LOGIC;
  signal x74_out_25 : STD_LOGIC;
  signal x74_out_24 : STD_LOGIC;
  signal x74_out_23 : STD_LOGIC;
  signal x74_out_22 : STD_LOGIC;
  signal x74_out_21 : STD_LOGIC;
  signal x74_out_20 : STD_LOGIC;
  signal x74_out_19 : STD_LOGIC;
  signal x74_out_18 : STD_LOGIC;
  signal x74_out_17 : STD_LOGIC;
  signal x74_out_16 : STD_LOGIC;
  signal x74_out_15 : STD_LOGIC;
  signal x74_out_14 : STD_LOGIC;
  signal x74_out_13 : STD_LOGIC;
  signal x74_out_12 : STD_LOGIC;
  signal x74_out_11 : STD_LOGIC;
  signal x74_out_10 : STD_LOGIC;
  signal x74_out_9 : STD_LOGIC;
  signal x74_out_8 : STD_LOGIC;
  signal x74_out_7 : STD_LOGIC;
  signal x74_out_6 : STD_LOGIC;
  signal x74_out_5 : STD_LOGIC;
  signal x74_out_4 : STD_LOGIC;
  signal x74_out_3 : STD_LOGIC;
  signal x74_out_2 : STD_LOGIC;
  signal x74_out_1 : STD_LOGIC;
  signal x74_out_0 : STD_LOGIC;
  signal x77_out_31 : STD_LOGIC;
  signal x77_out_30 : STD_LOGIC;
  signal x77_out_29 : STD_LOGIC;
  signal x77_out_28 : STD_LOGIC;
  signal x77_out_27 : STD_LOGIC;
  signal x77_out_26 : STD_LOGIC;
  signal x77_out_25 : STD_LOGIC;
  signal x77_out_24 : STD_LOGIC;
  signal x77_out_23 : STD_LOGIC;
  signal x77_out_22 : STD_LOGIC;
  signal x77_out_21 : STD_LOGIC;
  signal x77_out_20 : STD_LOGIC;
  signal x77_out_19 : STD_LOGIC;
  signal x77_out_18 : STD_LOGIC;
  signal x77_out_17 : STD_LOGIC;
  signal x77_out_16 : STD_LOGIC;
  signal x77_out_15 : STD_LOGIC;
  signal x77_out_14 : STD_LOGIC;
  signal x77_out_13 : STD_LOGIC;
  signal x77_out_12 : STD_LOGIC;
  signal x77_out_11 : STD_LOGIC;
  signal x77_out_10 : STD_LOGIC;
  signal x77_out_9 : STD_LOGIC;
  signal x77_out_8 : STD_LOGIC;
  signal x77_out_7 : STD_LOGIC;
  signal x77_out_6 : STD_LOGIC;
  signal x77_out_5 : STD_LOGIC;
  signal x77_out_4 : STD_LOGIC;
  signal x77_out_3 : STD_LOGIC;
  signal x77_out_2 : STD_LOGIC;
  signal x77_out_1 : STD_LOGIC;
  signal x77_out_0 : STD_LOGIC;
  signal x80_out_31 : STD_LOGIC;
  signal x80_out_30 : STD_LOGIC;
  signal x80_out_29 : STD_LOGIC;
  signal x80_out_28 : STD_LOGIC;
  signal x80_out_27 : STD_LOGIC;
  signal x80_out_26 : STD_LOGIC;
  signal x80_out_25 : STD_LOGIC;
  signal x80_out_24 : STD_LOGIC;
  signal x80_out_23 : STD_LOGIC;
  signal x80_out_22 : STD_LOGIC;
  signal x80_out_21 : STD_LOGIC;
  signal x80_out_20 : STD_LOGIC;
  signal x80_out_19 : STD_LOGIC;
  signal x80_out_18 : STD_LOGIC;
  signal x80_out_17 : STD_LOGIC;
  signal x80_out_16 : STD_LOGIC;
  signal x80_out_15 : STD_LOGIC;
  signal x80_out_14 : STD_LOGIC;
  signal x80_out_13 : STD_LOGIC;
  signal x80_out_12 : STD_LOGIC;
  signal x80_out_11 : STD_LOGIC;
  signal x80_out_10 : STD_LOGIC;
  signal x80_out_9 : STD_LOGIC;
  signal x80_out_8 : STD_LOGIC;
  signal x80_out_7 : STD_LOGIC;
  signal x80_out_6 : STD_LOGIC;
  signal x80_out_5 : STD_LOGIC;
  signal x80_out_4 : STD_LOGIC;
  signal x80_out_3 : STD_LOGIC;
  signal x80_out_2 : STD_LOGIC;
  signal x80_out_1 : STD_LOGIC;
  signal x80_out_0 : STD_LOGIC;
  signal x83_out_31 : STD_LOGIC;
  signal x83_out_30 : STD_LOGIC;
  signal x83_out_29 : STD_LOGIC;
  signal x83_out_28 : STD_LOGIC;
  signal x83_out_27 : STD_LOGIC;
  signal x83_out_26 : STD_LOGIC;
  signal x83_out_25 : STD_LOGIC;
  signal x83_out_24 : STD_LOGIC;
  signal x83_out_23 : STD_LOGIC;
  signal x83_out_22 : STD_LOGIC;
  signal x83_out_21 : STD_LOGIC;
  signal x83_out_20 : STD_LOGIC;
  signal x83_out_19 : STD_LOGIC;
  signal x83_out_18 : STD_LOGIC;
  signal x83_out_17 : STD_LOGIC;
  signal x83_out_16 : STD_LOGIC;
  signal x83_out_15 : STD_LOGIC;
  signal x83_out_14 : STD_LOGIC;
  signal x83_out_13 : STD_LOGIC;
  signal x83_out_12 : STD_LOGIC;
  signal x83_out_11 : STD_LOGIC;
  signal x83_out_10 : STD_LOGIC;
  signal x83_out_9 : STD_LOGIC;
  signal x83_out_8 : STD_LOGIC;
  signal x83_out_7 : STD_LOGIC;
  signal x83_out_6 : STD_LOGIC;
  signal x83_out_5 : STD_LOGIC;
  signal x83_out_4 : STD_LOGIC;
  signal x83_out_3 : STD_LOGIC;
  signal x83_out_2 : STD_LOGIC;
  signal x83_out_1 : STD_LOGIC;
  signal x83_out_0 : STD_LOGIC;
  signal x86_out_31 : STD_LOGIC;
  signal x86_out_30 : STD_LOGIC;
  signal x86_out_29 : STD_LOGIC;
  signal x86_out_28 : STD_LOGIC;
  signal x86_out_27 : STD_LOGIC;
  signal x86_out_26 : STD_LOGIC;
  signal x86_out_25 : STD_LOGIC;
  signal x86_out_24 : STD_LOGIC;
  signal x86_out_23 : STD_LOGIC;
  signal x86_out_22 : STD_LOGIC;
  signal x86_out_21 : STD_LOGIC;
  signal x86_out_20 : STD_LOGIC;
  signal x86_out_19 : STD_LOGIC;
  signal x86_out_18 : STD_LOGIC;
  signal x86_out_17 : STD_LOGIC;
  signal x86_out_16 : STD_LOGIC;
  signal x86_out_15 : STD_LOGIC;
  signal x86_out_14 : STD_LOGIC;
  signal x86_out_13 : STD_LOGIC;
  signal x86_out_12 : STD_LOGIC;
  signal x86_out_11 : STD_LOGIC;
  signal x86_out_10 : STD_LOGIC;
  signal x86_out_9 : STD_LOGIC;
  signal x86_out_8 : STD_LOGIC;
  signal x86_out_7 : STD_LOGIC;
  signal x86_out_6 : STD_LOGIC;
  signal x86_out_5 : STD_LOGIC;
  signal x86_out_4 : STD_LOGIC;
  signal x86_out_3 : STD_LOGIC;
  signal x86_out_2 : STD_LOGIC;
  signal x86_out_1 : STD_LOGIC;
  signal x86_out_0 : STD_LOGIC;
  signal x89_out_31 : STD_LOGIC;
  signal x89_out_30 : STD_LOGIC;
  signal x89_out_29 : STD_LOGIC;
  signal x89_out_28 : STD_LOGIC;
  signal x89_out_27 : STD_LOGIC;
  signal x89_out_26 : STD_LOGIC;
  signal x89_out_25 : STD_LOGIC;
  signal x89_out_24 : STD_LOGIC;
  signal x89_out_23 : STD_LOGIC;
  signal x89_out_22 : STD_LOGIC;
  signal x89_out_21 : STD_LOGIC;
  signal x89_out_20 : STD_LOGIC;
  signal x89_out_19 : STD_LOGIC;
  signal x89_out_18 : STD_LOGIC;
  signal x89_out_17 : STD_LOGIC;
  signal x89_out_16 : STD_LOGIC;
  signal x89_out_15 : STD_LOGIC;
  signal x89_out_14 : STD_LOGIC;
  signal x89_out_13 : STD_LOGIC;
  signal x89_out_12 : STD_LOGIC;
  signal x89_out_11 : STD_LOGIC;
  signal x89_out_10 : STD_LOGIC;
  signal x89_out_9 : STD_LOGIC;
  signal x89_out_8 : STD_LOGIC;
  signal x89_out_7 : STD_LOGIC;
  signal x89_out_6 : STD_LOGIC;
  signal x89_out_5 : STD_LOGIC;
  signal x89_out_4 : STD_LOGIC;
  signal x89_out_3 : STD_LOGIC;
  signal x89_out_2 : STD_LOGIC;
  signal x89_out_1 : STD_LOGIC;
  signal x89_out_0 : STD_LOGIC;
  signal x8_out_31 : STD_LOGIC;
  signal x8_out_30 : STD_LOGIC;
  signal x8_out_29 : STD_LOGIC;
  signal x8_out_28 : STD_LOGIC;
  signal x8_out_27 : STD_LOGIC;
  signal x8_out_26 : STD_LOGIC;
  signal x8_out_25 : STD_LOGIC;
  signal x8_out_24 : STD_LOGIC;
  signal x8_out_23 : STD_LOGIC;
  signal x8_out_22 : STD_LOGIC;
  signal x8_out_21 : STD_LOGIC;
  signal x8_out_20 : STD_LOGIC;
  signal x8_out_19 : STD_LOGIC;
  signal x8_out_18 : STD_LOGIC;
  signal x8_out_17 : STD_LOGIC;
  signal x8_out_16 : STD_LOGIC;
  signal x8_out_15 : STD_LOGIC;
  signal x8_out_14 : STD_LOGIC;
  signal x8_out_13 : STD_LOGIC;
  signal x8_out_12 : STD_LOGIC;
  signal x8_out_11 : STD_LOGIC;
  signal x8_out_10 : STD_LOGIC;
  signal x8_out_9 : STD_LOGIC;
  signal x8_out_8 : STD_LOGIC;
  signal x8_out_7 : STD_LOGIC;
  signal x8_out_6 : STD_LOGIC;
  signal x8_out_5 : STD_LOGIC;
  signal x8_out_4 : STD_LOGIC;
  signal x8_out_3 : STD_LOGIC;
  signal x8_out_2 : STD_LOGIC;
  signal x8_out_1 : STD_LOGIC;
  signal x8_out_0 : STD_LOGIC;
  signal x92_out_31 : STD_LOGIC;
  signal x92_out_30 : STD_LOGIC;
  signal x92_out_29 : STD_LOGIC;
  signal x92_out_28 : STD_LOGIC;
  signal x92_out_27 : STD_LOGIC;
  signal x92_out_26 : STD_LOGIC;
  signal x92_out_25 : STD_LOGIC;
  signal x92_out_24 : STD_LOGIC;
  signal x92_out_23 : STD_LOGIC;
  signal x92_out_22 : STD_LOGIC;
  signal x92_out_21 : STD_LOGIC;
  signal x92_out_20 : STD_LOGIC;
  signal x92_out_19 : STD_LOGIC;
  signal x92_out_18 : STD_LOGIC;
  signal x92_out_17 : STD_LOGIC;
  signal x92_out_16 : STD_LOGIC;
  signal x92_out_15 : STD_LOGIC;
  signal x92_out_14 : STD_LOGIC;
  signal x92_out_13 : STD_LOGIC;
  signal x92_out_12 : STD_LOGIC;
  signal x92_out_11 : STD_LOGIC;
  signal x92_out_10 : STD_LOGIC;
  signal x92_out_9 : STD_LOGIC;
  signal x92_out_8 : STD_LOGIC;
  signal x92_out_7 : STD_LOGIC;
  signal x92_out_6 : STD_LOGIC;
  signal x92_out_5 : STD_LOGIC;
  signal x92_out_4 : STD_LOGIC;
  signal x92_out_3 : STD_LOGIC;
  signal x92_out_2 : STD_LOGIC;
  signal x92_out_1 : STD_LOGIC;
  signal x92_out_0 : STD_LOGIC;
  signal x94_out_31 : STD_LOGIC;
  signal x94_out_30 : STD_LOGIC;
  signal x94_out_29 : STD_LOGIC;
  signal x94_out_28 : STD_LOGIC;
  signal x94_out_27 : STD_LOGIC;
  signal x94_out_26 : STD_LOGIC;
  signal x94_out_25 : STD_LOGIC;
  signal x94_out_24 : STD_LOGIC;
  signal x94_out_23 : STD_LOGIC;
  signal x94_out_22 : STD_LOGIC;
  signal x94_out_21 : STD_LOGIC;
  signal x94_out_20 : STD_LOGIC;
  signal x94_out_19 : STD_LOGIC;
  signal x94_out_18 : STD_LOGIC;
  signal x94_out_17 : STD_LOGIC;
  signal x94_out_16 : STD_LOGIC;
  signal x94_out_15 : STD_LOGIC;
  signal x94_out_14 : STD_LOGIC;
  signal x94_out_13 : STD_LOGIC;
  signal x94_out_12 : STD_LOGIC;
  signal x94_out_11 : STD_LOGIC;
  signal x94_out_10 : STD_LOGIC;
  signal x94_out_9 : STD_LOGIC;
  signal x94_out_8 : STD_LOGIC;
  signal x94_out_7 : STD_LOGIC;
  signal x94_out_6 : STD_LOGIC;
  signal x94_out_5 : STD_LOGIC;
  signal x94_out_4 : STD_LOGIC;
  signal x94_out_3 : STD_LOGIC;
  signal x94_out_2 : STD_LOGIC;
  signal x94_out_1 : STD_LOGIC;
  signal x94_out_0 : STD_LOGIC;
  signal x96_out_31 : STD_LOGIC;
  signal x96_out_30 : STD_LOGIC;
  signal x96_out_29 : STD_LOGIC;
  signal x96_out_28 : STD_LOGIC;
  signal x96_out_27 : STD_LOGIC;
  signal x96_out_26 : STD_LOGIC;
  signal x96_out_25 : STD_LOGIC;
  signal x96_out_24 : STD_LOGIC;
  signal x96_out_23 : STD_LOGIC;
  signal x96_out_22 : STD_LOGIC;
  signal x96_out_21 : STD_LOGIC;
  signal x96_out_20 : STD_LOGIC;
  signal x96_out_19 : STD_LOGIC;
  signal x96_out_18 : STD_LOGIC;
  signal x96_out_17 : STD_LOGIC;
  signal x96_out_16 : STD_LOGIC;
  signal x96_out_15 : STD_LOGIC;
  signal x96_out_14 : STD_LOGIC;
  signal x96_out_13 : STD_LOGIC;
  signal x96_out_12 : STD_LOGIC;
  signal x96_out_11 : STD_LOGIC;
  signal x96_out_10 : STD_LOGIC;
  signal x96_out_9 : STD_LOGIC;
  signal x96_out_8 : STD_LOGIC;
  signal x96_out_7 : STD_LOGIC;
  signal x96_out_6 : STD_LOGIC;
  signal x96_out_5 : STD_LOGIC;
  signal x96_out_4 : STD_LOGIC;
  signal x96_out_3 : STD_LOGIC;
  signal x96_out_2 : STD_LOGIC;
  signal x96_out_1 : STD_LOGIC;
  signal x96_out_0 : STD_LOGIC;
  signal x98_out_31 : STD_LOGIC;
  signal x98_out_30 : STD_LOGIC;
  signal x98_out_29 : STD_LOGIC;
  signal x98_out_28 : STD_LOGIC;
  signal x98_out_27 : STD_LOGIC;
  signal x98_out_26 : STD_LOGIC;
  signal x98_out_25 : STD_LOGIC;
  signal x98_out_24 : STD_LOGIC;
  signal x98_out_23 : STD_LOGIC;
  signal x98_out_22 : STD_LOGIC;
  signal x98_out_21 : STD_LOGIC;
  signal x98_out_20 : STD_LOGIC;
  signal x98_out_19 : STD_LOGIC;
  signal x98_out_18 : STD_LOGIC;
  signal x98_out_17 : STD_LOGIC;
  signal x98_out_16 : STD_LOGIC;
  signal x98_out_15 : STD_LOGIC;
  signal x98_out_14 : STD_LOGIC;
  signal x98_out_13 : STD_LOGIC;
  signal x98_out_12 : STD_LOGIC;
  signal x98_out_11 : STD_LOGIC;
  signal x98_out_10 : STD_LOGIC;
  signal x98_out_9 : STD_LOGIC;
  signal x98_out_8 : STD_LOGIC;
  signal x98_out_7 : STD_LOGIC;
  signal x98_out_6 : STD_LOGIC;
  signal x98_out_5 : STD_LOGIC;
  signal x98_out_4 : STD_LOGIC;
  signal x98_out_3 : STD_LOGIC;
  signal x98_out_2 : STD_LOGIC;
  signal x98_out_1 : STD_LOGIC;
  signal x98_out_0 : STD_LOGIC;
begin
a_0_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in7_0,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_224,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => a_0_i_1_n_0
);
a_10_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in7_10,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_234,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => a_10_i_1_n_0
);
a_11_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in7_11,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_235,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => a_11_i_1_n_0
);
a_11_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => T1_0_11,
   I1 => T2_11,
   O => a_11_i_3_n_0
);
a_11_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => T1_0_10,
   I1 => T2_10,
   O => a_11_i_4_n_0
);
a_11_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => T1_0_9,
   I1 => T2_9,
   O => a_11_i_5_n_0
);
a_11_i_6 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => T1_0_8,
   I1 => T2_8,
   O => a_11_i_6_n_0
);
a_12_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in7_12,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_236,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => a_12_i_1_n_0
);
a_13_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in7_13,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_237,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => a_13_i_1_n_0
);
a_14_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in7_14,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_238,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => a_14_i_1_n_0
);
a_15_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in7_15,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_239,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => a_15_i_1_n_0
);
a_15_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => T1_0_15,
   I1 => T2_15,
   O => a_15_i_3_n_0
);
a_15_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => T1_0_14,
   I1 => T2_14,
   O => a_15_i_4_n_0
);
a_15_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => T1_0_13,
   I1 => T2_13,
   O => a_15_i_5_n_0
);
a_15_i_6 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => T1_0_12,
   I1 => T2_12,
   O => a_15_i_6_n_0
);
a_16_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in7_16,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_240,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => a_16_i_1_n_0
);
a_17_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in7_17,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_241,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => a_17_i_1_n_0
);
a_18_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in7_18,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_242,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => a_18_i_1_n_0
);
a_19_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in7_19,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_243,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => a_19_i_1_n_0
);
a_19_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => T1_0_19,
   I1 => T2_19,
   O => a_19_i_3_n_0
);
a_19_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => T1_0_18,
   I1 => T2_18,
   O => a_19_i_4_n_0
);
a_19_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => T1_0_17,
   I1 => T2_17,
   O => a_19_i_5_n_0
);
a_19_i_6 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => T1_0_16,
   I1 => T2_16,
   O => a_19_i_6_n_0
);
a_1_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in7_1,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_225,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => a_1_i_1_n_0
);
a_20_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in7_20,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_244,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => a_20_i_1_n_0
);
a_21_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in7_21,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_245,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => a_21_i_1_n_0
);
a_22_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in7_22,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_246,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => a_22_i_1_n_0
);
a_23_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in7_23,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_247,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => a_23_i_1_n_0
);
a_23_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => T1_0_23,
   I1 => T2_23,
   O => a_23_i_3_n_0
);
a_23_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => T1_0_22,
   I1 => T2_22,
   O => a_23_i_4_n_0
);
a_23_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => T1_0_21,
   I1 => T2_21,
   O => a_23_i_5_n_0
);
a_23_i_6 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => T1_0_20,
   I1 => T2_20,
   O => a_23_i_6_n_0
);
a_24_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in7_24,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_248,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => a_24_i_1_n_0
);
a_25_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in7_25,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_249,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => a_25_i_1_n_0
);
a_26_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in7_26,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_250,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => a_26_i_1_n_0
);
a_27_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in7_27,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_251,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => a_27_i_1_n_0
);
a_27_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => T1_0_27,
   I1 => T2_27,
   O => a_27_i_3_n_0
);
a_27_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => T1_0_26,
   I1 => T2_26,
   O => a_27_i_4_n_0
);
a_27_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => T1_0_25,
   I1 => T2_25,
   O => a_27_i_5_n_0
);
a_27_i_6 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => T1_0_24,
   I1 => T2_24,
   O => a_27_i_6_n_0
);
a_28_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in7_28,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_252,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => a_28_i_1_n_0
);
a_29_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in7_29,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_253,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => a_29_i_1_n_0
);
a_2_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in7_2,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_226,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => a_2_i_1_n_0
);
a_30_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in7_30,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_254,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => a_30_i_1_n_0
);
a_31_i_1 : LUT3
  generic map(
   INIT => X"54"
  )
 port map (
   I0 => rst_IBUF,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   I2 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   O => a_31_i_1_n_0
);
a_31_i_2 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in7_31,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_255,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => a_31_i_2_n_0
);
a_31_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => T2_31,
   I1 => T1_0_31,
   O => a_31_i_4_n_0
);
a_31_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => T1_0_30,
   I1 => T2_30,
   O => a_31_i_5_n_0
);
a_31_i_6 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => T1_0_29,
   I1 => T2_29,
   O => a_31_i_6_n_0
);
a_31_i_7 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => T1_0_28,
   I1 => T2_28,
   O => a_31_i_7_n_0
);
a_3_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in7_3,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_227,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => a_3_i_1_n_0
);
a_3_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => T1_0_3,
   I1 => T2_3,
   O => a_3_i_3_n_0
);
a_3_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => T1_0_2,
   I1 => T2_2,
   O => a_3_i_4_n_0
);
a_3_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => T1_0_1,
   I1 => T2_1,
   O => a_3_i_5_n_0
);
a_3_i_6 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => T1_0_0,
   I1 => T2_0,
   O => a_3_i_6_n_0
);
a_4_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in7_4,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_228,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => a_4_i_1_n_0
);
a_5_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in7_5,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_229,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => a_5_i_1_n_0
);
a_6_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in7_6,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_230,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => a_6_i_1_n_0
);
a_7_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in7_7,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_231,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => a_7_i_1_n_0
);
a_7_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => T1_0_7,
   I1 => T2_7,
   O => a_7_i_3_n_0
);
a_7_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => T1_0_6,
   I1 => T2_6,
   O => a_7_i_4_n_0
);
a_7_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => T1_0_5,
   I1 => T2_5,
   O => a_7_i_5_n_0
);
a_7_i_6 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => T1_0_4,
   I1 => T2_4,
   O => a_7_i_6_n_0
);
a_8_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in7_8,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_232,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => a_8_i_1_n_0
);
a_9_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in7_9,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_233,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => a_9_i_1_n_0
);
a_reg_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => a_0_i_1_n_0,
   R => '0',
   Q => ROTR2_out_13
);
a_reg_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => a_10_i_1_n_0,
   R => '0',
   Q => ROTR2_out_3
);
a_reg_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => a_11_i_1_n_0,
   R => '0',
   Q => ROTR2_out_2
);
a_reg_11_i_2 : CARRY4
 port map (
   CI => a_reg_7_i_2_n_0,
   CYINIT => '0',
   DI(0) => T1_0_8,
   DI(1) => T1_0_9,
   DI(2) => T1_0_10,
   DI(3) => T1_0_11,
   S(0) => a_11_i_6_n_0,
   S(1) => a_11_i_5_n_0,
   S(2) => a_11_i_4_n_0,
   S(3) => a_11_i_3_n_0,
   CO(0) => a_reg_11_i_2_n_3,
   CO(1) => a_reg_11_i_2_n_2,
   CO(2) => a_reg_11_i_2_n_1,
   CO(3) => a_reg_11_i_2_n_0,
   O(0) => in7_8,
   O(1) => in7_9,
   O(2) => in7_10,
   O(3) => in7_11
);
a_reg_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => a_12_i_1_n_0,
   R => '0',
   Q => ROTR2_out_1
);
a_reg_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => a_13_i_1_n_0,
   R => '0',
   Q => ROTR2_out_32
);
a_reg_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => a_14_i_1_n_0,
   R => '0',
   Q => ROTR2_out_31
);
a_reg_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => a_15_i_1_n_0,
   R => '0',
   Q => ROTR2_out_30
);
a_reg_15_i_2 : CARRY4
 port map (
   CI => a_reg_11_i_2_n_0,
   CYINIT => '0',
   DI(0) => T1_0_12,
   DI(1) => T1_0_13,
   DI(2) => T1_0_14,
   DI(3) => T1_0_15,
   S(0) => a_15_i_6_n_0,
   S(1) => a_15_i_5_n_0,
   S(2) => a_15_i_4_n_0,
   S(3) => a_15_i_3_n_0,
   CO(0) => a_reg_15_i_2_n_3,
   CO(1) => a_reg_15_i_2_n_2,
   CO(2) => a_reg_15_i_2_n_1,
   CO(3) => a_reg_15_i_2_n_0,
   O(0) => in7_12,
   O(1) => in7_13,
   O(2) => in7_14,
   O(3) => in7_15
);
a_reg_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => a_16_i_1_n_0,
   R => '0',
   Q => ROTR2_out_29
);
a_reg_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => a_17_i_1_n_0,
   R => '0',
   Q => ROTR2_out_28
);
a_reg_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => a_18_i_1_n_0,
   R => '0',
   Q => ROTR2_out_27
);
a_reg_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => a_19_i_1_n_0,
   R => '0',
   Q => ROTR2_out_26
);
a_reg_19_i_2 : CARRY4
 port map (
   CI => a_reg_15_i_2_n_0,
   CYINIT => '0',
   DI(0) => T1_0_16,
   DI(1) => T1_0_17,
   DI(2) => T1_0_18,
   DI(3) => T1_0_19,
   S(0) => a_19_i_6_n_0,
   S(1) => a_19_i_5_n_0,
   S(2) => a_19_i_4_n_0,
   S(3) => a_19_i_3_n_0,
   CO(0) => a_reg_19_i_2_n_3,
   CO(1) => a_reg_19_i_2_n_2,
   CO(2) => a_reg_19_i_2_n_1,
   CO(3) => a_reg_19_i_2_n_0,
   O(0) => in7_16,
   O(1) => in7_17,
   O(2) => in7_18,
   O(3) => in7_19
);
a_reg_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => a_1_i_1_n_0,
   R => '0',
   Q => ROTR2_out_12
);
a_reg_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => a_20_i_1_n_0,
   R => '0',
   Q => ROTR2_out_25
);
a_reg_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => a_21_i_1_n_0,
   R => '0',
   Q => ROTR2_out_24
);
a_reg_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => a_22_i_1_n_0,
   R => '0',
   Q => ROTR2_out_23
);
a_reg_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => a_23_i_1_n_0,
   R => '0',
   Q => ROTR2_out_22
);
a_reg_23_i_2 : CARRY4
 port map (
   CI => a_reg_19_i_2_n_0,
   CYINIT => '0',
   DI(0) => T1_0_20,
   DI(1) => T1_0_21,
   DI(2) => T1_0_22,
   DI(3) => T1_0_23,
   S(0) => a_23_i_6_n_0,
   S(1) => a_23_i_5_n_0,
   S(2) => a_23_i_4_n_0,
   S(3) => a_23_i_3_n_0,
   CO(0) => a_reg_23_i_2_n_3,
   CO(1) => a_reg_23_i_2_n_2,
   CO(2) => a_reg_23_i_2_n_1,
   CO(3) => a_reg_23_i_2_n_0,
   O(0) => in7_20,
   O(1) => in7_21,
   O(2) => in7_22,
   O(3) => in7_23
);
a_reg_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => a_24_i_1_n_0,
   R => '0',
   Q => ROTR2_out_21
);
a_reg_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => a_25_i_1_n_0,
   R => '0',
   Q => ROTR2_out_20
);
a_reg_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => a_26_i_1_n_0,
   R => '0',
   Q => ROTR2_out_19
);
a_reg_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => a_27_i_1_n_0,
   R => '0',
   Q => ROTR2_out_18
);
a_reg_27_i_2 : CARRY4
 port map (
   CI => a_reg_23_i_2_n_0,
   CYINIT => '0',
   DI(0) => T1_0_24,
   DI(1) => T1_0_25,
   DI(2) => T1_0_26,
   DI(3) => T1_0_27,
   S(0) => a_27_i_6_n_0,
   S(1) => a_27_i_5_n_0,
   S(2) => a_27_i_4_n_0,
   S(3) => a_27_i_3_n_0,
   CO(0) => a_reg_27_i_2_n_3,
   CO(1) => a_reg_27_i_2_n_2,
   CO(2) => a_reg_27_i_2_n_1,
   CO(3) => a_reg_27_i_2_n_0,
   O(0) => in7_24,
   O(1) => in7_25,
   O(2) => in7_26,
   O(3) => in7_27
);
a_reg_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => a_28_i_1_n_0,
   R => '0',
   Q => ROTR2_out_17
);
a_reg_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => a_29_i_1_n_0,
   R => '0',
   Q => ROTR2_out_16
);
a_reg_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => a_2_i_1_n_0,
   R => '0',
   Q => ROTR2_out_11
);
a_reg_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => a_30_i_1_n_0,
   R => '0',
   Q => ROTR2_out_15
);
a_reg_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => a_31_i_2_n_0,
   R => '0',
   Q => ROTR2_out_14
);
a_reg_31_i_3 : CARRY4
 port map (
   CI => a_reg_27_i_2_n_0,
   CYINIT => '0',
   DI(0) => T1_0_28,
   DI(1) => T1_0_29,
   DI(2) => T1_0_30,
   DI(3) => '0',
   S(0) => a_31_i_7_n_0,
   S(1) => a_31_i_6_n_0,
   S(2) => a_31_i_5_n_0,
   S(3) => a_31_i_4_n_0,
   CO(0) => a_reg_31_i_3_n_3,
   CO(1) => a_reg_31_i_3_n_2,
   CO(2) => a_reg_31_i_3_n_1,
   CO(3) => NLW_a_reg_31_i_3_CO_UNCONNECTED_3,
   O(0) => in7_28,
   O(1) => in7_29,
   O(2) => in7_30,
   O(3) => in7_31
);
a_reg_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => a_3_i_1_n_0,
   R => '0',
   Q => ROTR2_out_10
);
a_reg_3_i_2 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => T1_0_0,
   DI(1) => T1_0_1,
   DI(2) => T1_0_2,
   DI(3) => T1_0_3,
   S(0) => a_3_i_6_n_0,
   S(1) => a_3_i_5_n_0,
   S(2) => a_3_i_4_n_0,
   S(3) => a_3_i_3_n_0,
   CO(0) => a_reg_3_i_2_n_3,
   CO(1) => a_reg_3_i_2_n_2,
   CO(2) => a_reg_3_i_2_n_1,
   CO(3) => a_reg_3_i_2_n_0,
   O(0) => in7_0,
   O(1) => in7_1,
   O(2) => in7_2,
   O(3) => in7_3
);
a_reg_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => a_4_i_1_n_0,
   R => '0',
   Q => ROTR2_out_9
);
a_reg_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => a_5_i_1_n_0,
   R => '0',
   Q => ROTR2_out_8
);
a_reg_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => a_6_i_1_n_0,
   R => '0',
   Q => ROTR2_out_7
);
a_reg_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => a_7_i_1_n_0,
   R => '0',
   Q => ROTR2_out_6
);
a_reg_7_i_2 : CARRY4
 port map (
   CI => a_reg_3_i_2_n_0,
   CYINIT => '0',
   DI(0) => T1_0_4,
   DI(1) => T1_0_5,
   DI(2) => T1_0_6,
   DI(3) => T1_0_7,
   S(0) => a_7_i_6_n_0,
   S(1) => a_7_i_5_n_0,
   S(2) => a_7_i_4_n_0,
   S(3) => a_7_i_3_n_0,
   CO(0) => a_reg_7_i_2_n_3,
   CO(1) => a_reg_7_i_2_n_2,
   CO(2) => a_reg_7_i_2_n_1,
   CO(3) => a_reg_7_i_2_n_0,
   O(0) => in7_4,
   O(1) => in7_5,
   O(2) => in7_6,
   O(3) => in7_7
);
a_reg_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => a_8_i_1_n_0,
   R => '0',
   Q => ROTR2_out_5
);
a_reg_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => a_9_i_1_n_0,
   R => '0',
   Q => ROTR2_out_4
);
b_0_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I1 => ROTR2_out_13,
   I2 => data_out_OBUF_192,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => b_0_i_1_n_0
);
b_10_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I1 => ROTR2_out_3,
   I2 => data_out_OBUF_202,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => b_10_i_1_n_0
);
b_11_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I1 => ROTR2_out_2,
   I2 => data_out_OBUF_203,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => b_11_i_1_n_0
);
b_12_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I1 => ROTR2_out_1,
   I2 => data_out_OBUF_204,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => b_12_i_1_n_0
);
b_13_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I1 => ROTR2_out_32,
   I2 => data_out_OBUF_205,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => b_13_i_1_n_0
);
b_14_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I1 => ROTR2_out_31,
   I2 => data_out_OBUF_206,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => b_14_i_1_n_0
);
b_15_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I1 => ROTR2_out_30,
   I2 => data_out_OBUF_207,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => b_15_i_1_n_0
);
b_16_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I1 => ROTR2_out_29,
   I2 => data_out_OBUF_208,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => b_16_i_1_n_0
);
b_17_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I1 => ROTR2_out_28,
   I2 => data_out_OBUF_209,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => b_17_i_1_n_0
);
b_18_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I1 => ROTR2_out_27,
   I2 => data_out_OBUF_210,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => b_18_i_1_n_0
);
b_19_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I1 => ROTR2_out_26,
   I2 => data_out_OBUF_211,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => b_19_i_1_n_0
);
b_1_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I1 => ROTR2_out_12,
   I2 => data_out_OBUF_193,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => b_1_i_1_n_0
);
b_20_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I1 => ROTR2_out_25,
   I2 => data_out_OBUF_212,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => b_20_i_1_n_0
);
b_21_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I1 => ROTR2_out_24,
   I2 => data_out_OBUF_213,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => b_21_i_1_n_0
);
b_22_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I1 => ROTR2_out_23,
   I2 => data_out_OBUF_214,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => b_22_i_1_n_0
);
b_23_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I1 => ROTR2_out_22,
   I2 => data_out_OBUF_215,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => b_23_i_1_n_0
);
b_24_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I1 => ROTR2_out_21,
   I2 => data_out_OBUF_216,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => b_24_i_1_n_0
);
b_25_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I1 => ROTR2_out_20,
   I2 => data_out_OBUF_217,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => b_25_i_1_n_0
);
b_26_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I1 => ROTR2_out_19,
   I2 => data_out_OBUF_218,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => b_26_i_1_n_0
);
b_27_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I1 => ROTR2_out_18,
   I2 => data_out_OBUF_219,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => b_27_i_1_n_0
);
b_28_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I1 => ROTR2_out_17,
   I2 => data_out_OBUF_220,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => b_28_i_1_n_0
);
b_29_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I1 => ROTR2_out_16,
   I2 => data_out_OBUF_221,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => b_29_i_1_n_0
);
b_2_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I1 => ROTR2_out_11,
   I2 => data_out_OBUF_194,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => b_2_i_1_n_0
);
b_30_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I1 => ROTR2_out_15,
   I2 => data_out_OBUF_222,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => b_30_i_1_n_0
);
b_31_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I1 => ROTR2_out_14,
   I2 => data_out_OBUF_223,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => b_31_i_1_n_0
);
b_3_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I1 => ROTR2_out_10,
   I2 => data_out_OBUF_195,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => b_3_i_1_n_0
);
b_4_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I1 => ROTR2_out_9,
   I2 => data_out_OBUF_196,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => b_4_i_1_n_0
);
b_5_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I1 => ROTR2_out_8,
   I2 => data_out_OBUF_197,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => b_5_i_1_n_0
);
b_6_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I1 => ROTR2_out_7,
   I2 => data_out_OBUF_198,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => b_6_i_1_n_0
);
b_7_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I1 => ROTR2_out_6,
   I2 => data_out_OBUF_199,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => b_7_i_1_n_0
);
b_8_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I1 => ROTR2_out_5,
   I2 => data_out_OBUF_200,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => b_8_i_1_n_0
);
b_9_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I1 => ROTR2_out_4,
   I2 => data_out_OBUF_201,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => b_9_i_1_n_0
);
b_reg_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => b_0_i_1_n_0,
   R => '0',
   Q => b_reg_n_0_0
);
b_reg_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => b_10_i_1_n_0,
   R => '0',
   Q => b_reg_n_0_10
);
b_reg_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => b_11_i_1_n_0,
   R => '0',
   Q => b_reg_n_0_11
);
b_reg_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => b_12_i_1_n_0,
   R => '0',
   Q => b_reg_n_0_12
);
b_reg_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => b_13_i_1_n_0,
   R => '0',
   Q => b_reg_n_0_13
);
b_reg_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => b_14_i_1_n_0,
   R => '0',
   Q => b_reg_n_0_14
);
b_reg_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => b_15_i_1_n_0,
   R => '0',
   Q => b_reg_n_0_15
);
b_reg_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => b_16_i_1_n_0,
   R => '0',
   Q => b_reg_n_0_16
);
b_reg_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => b_17_i_1_n_0,
   R => '0',
   Q => b_reg_n_0_17
);
b_reg_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => b_18_i_1_n_0,
   R => '0',
   Q => b_reg_n_0_18
);
b_reg_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => b_19_i_1_n_0,
   R => '0',
   Q => b_reg_n_0_19
);
b_reg_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => b_1_i_1_n_0,
   R => '0',
   Q => b_reg_n_0_1
);
b_reg_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => b_20_i_1_n_0,
   R => '0',
   Q => b_reg_n_0_20
);
b_reg_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => b_21_i_1_n_0,
   R => '0',
   Q => b_reg_n_0_21
);
b_reg_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => b_22_i_1_n_0,
   R => '0',
   Q => b_reg_n_0_22
);
b_reg_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => b_23_i_1_n_0,
   R => '0',
   Q => b_reg_n_0_23
);
b_reg_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => b_24_i_1_n_0,
   R => '0',
   Q => b_reg_n_0_24
);
b_reg_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => b_25_i_1_n_0,
   R => '0',
   Q => b_reg_n_0_25
);
b_reg_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => b_26_i_1_n_0,
   R => '0',
   Q => b_reg_n_0_26
);
b_reg_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => b_27_i_1_n_0,
   R => '0',
   Q => b_reg_n_0_27
);
b_reg_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => b_28_i_1_n_0,
   R => '0',
   Q => b_reg_n_0_28
);
b_reg_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => b_29_i_1_n_0,
   R => '0',
   Q => b_reg_n_0_29
);
b_reg_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => b_2_i_1_n_0,
   R => '0',
   Q => b_reg_n_0_2
);
b_reg_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => b_30_i_1_n_0,
   R => '0',
   Q => b_reg_n_0_30
);
b_reg_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => b_31_i_1_n_0,
   R => '0',
   Q => b_reg_n_0_31
);
b_reg_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => b_3_i_1_n_0,
   R => '0',
   Q => b_reg_n_0_3
);
b_reg_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => b_4_i_1_n_0,
   R => '0',
   Q => b_reg_n_0_4
);
b_reg_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => b_5_i_1_n_0,
   R => '0',
   Q => b_reg_n_0_5
);
b_reg_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => b_6_i_1_n_0,
   R => '0',
   Q => b_reg_n_0_6
);
b_reg_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => b_7_i_1_n_0,
   R => '0',
   Q => b_reg_n_0_7
);
b_reg_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => b_8_i_1_n_0,
   R => '0',
   Q => b_reg_n_0_8
);
b_reg_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => b_9_i_1_n_0,
   R => '0',
   Q => b_reg_n_0_9
);
clk_IBUF_BUFG_inst : BUFG
 port map (
   I => clk_IBUF,
   O => clk_IBUF_BUFG
);
clk_IBUF_inst : IBUF
 port map (
   I => clk,
   O => clk_IBUF
);
c_0_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => b_reg_n_0_0,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_160,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => c_0_i_1_n_0
);
c_10_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => b_reg_n_0_10,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_170,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => c_10_i_1_n_0
);
c_11_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => b_reg_n_0_11,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_171,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => c_11_i_1_n_0
);
c_12_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => b_reg_n_0_12,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_172,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => c_12_i_1_n_0
);
c_13_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => b_reg_n_0_13,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_173,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => c_13_i_1_n_0
);
c_14_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => b_reg_n_0_14,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_174,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => c_14_i_1_n_0
);
c_15_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => b_reg_n_0_15,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_175,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => c_15_i_1_n_0
);
c_16_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => b_reg_n_0_16,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_176,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => c_16_i_1_n_0
);
c_17_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => b_reg_n_0_17,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_177,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => c_17_i_1_n_0
);
c_18_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => b_reg_n_0_18,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_178,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => c_18_i_1_n_0
);
c_19_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => b_reg_n_0_19,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_179,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => c_19_i_1_n_0
);
c_1_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => b_reg_n_0_1,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_161,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => c_1_i_1_n_0
);
c_20_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => b_reg_n_0_20,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_180,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => c_20_i_1_n_0
);
c_21_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => b_reg_n_0_21,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_181,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => c_21_i_1_n_0
);
c_22_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => b_reg_n_0_22,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_182,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => c_22_i_1_n_0
);
c_23_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => b_reg_n_0_23,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_183,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => c_23_i_1_n_0
);
c_24_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => b_reg_n_0_24,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_184,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => c_24_i_1_n_0
);
c_25_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => b_reg_n_0_25,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_185,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => c_25_i_1_n_0
);
c_26_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => b_reg_n_0_26,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_186,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => c_26_i_1_n_0
);
c_27_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => b_reg_n_0_27,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_187,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => c_27_i_1_n_0
);
c_28_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => b_reg_n_0_28,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_188,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => c_28_i_1_n_0
);
c_29_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => b_reg_n_0_29,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_189,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => c_29_i_1_n_0
);
c_2_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => b_reg_n_0_2,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_162,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => c_2_i_1_n_0
);
c_30_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => b_reg_n_0_30,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_190,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => c_30_i_1_n_0
);
c_31_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => b_reg_n_0_31,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_191,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => c_31_i_1_n_0
);
c_3_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => b_reg_n_0_3,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_163,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => c_3_i_1_n_0
);
c_4_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => b_reg_n_0_4,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_164,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => c_4_i_1_n_0
);
c_5_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => b_reg_n_0_5,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_165,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => c_5_i_1_n_0
);
c_6_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => b_reg_n_0_6,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_166,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => c_6_i_1_n_0
);
c_7_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => b_reg_n_0_7,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_167,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => c_7_i_1_n_0
);
c_8_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => b_reg_n_0_8,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_168,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => c_8_i_1_n_0
);
c_9_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => b_reg_n_0_9,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_169,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => c_9_i_1_n_0
);
c_reg_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => c_0_i_1_n_0,
   R => '0',
   Q => c_reg_n_0_0
);
c_reg_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => c_10_i_1_n_0,
   R => '0',
   Q => c_reg_n_0_10
);
c_reg_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => c_11_i_1_n_0,
   R => '0',
   Q => c_reg_n_0_11
);
c_reg_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => c_12_i_1_n_0,
   R => '0',
   Q => c_reg_n_0_12
);
c_reg_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => c_13_i_1_n_0,
   R => '0',
   Q => c_reg_n_0_13
);
c_reg_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => c_14_i_1_n_0,
   R => '0',
   Q => c_reg_n_0_14
);
c_reg_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => c_15_i_1_n_0,
   R => '0',
   Q => c_reg_n_0_15
);
c_reg_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => c_16_i_1_n_0,
   R => '0',
   Q => c_reg_n_0_16
);
c_reg_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => c_17_i_1_n_0,
   R => '0',
   Q => c_reg_n_0_17
);
c_reg_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => c_18_i_1_n_0,
   R => '0',
   Q => c_reg_n_0_18
);
c_reg_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => c_19_i_1_n_0,
   R => '0',
   Q => c_reg_n_0_19
);
c_reg_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => c_1_i_1_n_0,
   R => '0',
   Q => c_reg_n_0_1
);
c_reg_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => c_20_i_1_n_0,
   R => '0',
   Q => c_reg_n_0_20
);
c_reg_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => c_21_i_1_n_0,
   R => '0',
   Q => c_reg_n_0_21
);
c_reg_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => c_22_i_1_n_0,
   R => '0',
   Q => c_reg_n_0_22
);
c_reg_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => c_23_i_1_n_0,
   R => '0',
   Q => c_reg_n_0_23
);
c_reg_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => c_24_i_1_n_0,
   R => '0',
   Q => c_reg_n_0_24
);
c_reg_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => c_25_i_1_n_0,
   R => '0',
   Q => c_reg_n_0_25
);
c_reg_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => c_26_i_1_n_0,
   R => '0',
   Q => c_reg_n_0_26
);
c_reg_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => c_27_i_1_n_0,
   R => '0',
   Q => c_reg_n_0_27
);
c_reg_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => c_28_i_1_n_0,
   R => '0',
   Q => c_reg_n_0_28
);
c_reg_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => c_29_i_1_n_0,
   R => '0',
   Q => c_reg_n_0_29
);
c_reg_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => c_2_i_1_n_0,
   R => '0',
   Q => c_reg_n_0_2
);
c_reg_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => c_30_i_1_n_0,
   R => '0',
   Q => c_reg_n_0_30
);
c_reg_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => c_31_i_1_n_0,
   R => '0',
   Q => c_reg_n_0_31
);
c_reg_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => c_3_i_1_n_0,
   R => '0',
   Q => c_reg_n_0_3
);
c_reg_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => c_4_i_1_n_0,
   R => '0',
   Q => c_reg_n_0_4
);
c_reg_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => c_5_i_1_n_0,
   R => '0',
   Q => c_reg_n_0_5
);
c_reg_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => c_6_i_1_n_0,
   R => '0',
   Q => c_reg_n_0_6
);
c_reg_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => c_7_i_1_n_0,
   R => '0',
   Q => c_reg_n_0_7
);
c_reg_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => c_8_i_1_n_0,
   R => '0',
   Q => c_reg_n_0_8
);
c_reg_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => c_9_i_1_n_0,
   R => '0',
   Q => c_reg_n_0_9
);
data_out_OBUF_0_inst : OBUF
 port map (
   I => data_out_OBUF_0,
   O => data_out_0
);
data_out_OBUF_100_inst : OBUF
 port map (
   I => data_out_OBUF_100,
   O => data_out_100
);
data_out_OBUF_101_inst : OBUF
 port map (
   I => data_out_OBUF_101,
   O => data_out_101
);
data_out_OBUF_102_inst : OBUF
 port map (
   I => data_out_OBUF_102,
   O => data_out_102
);
data_out_OBUF_103_inst : OBUF
 port map (
   I => data_out_OBUF_103,
   O => data_out_103
);
data_out_OBUF_104_inst : OBUF
 port map (
   I => data_out_OBUF_104,
   O => data_out_104
);
data_out_OBUF_105_inst : OBUF
 port map (
   I => data_out_OBUF_105,
   O => data_out_105
);
data_out_OBUF_106_inst : OBUF
 port map (
   I => data_out_OBUF_106,
   O => data_out_106
);
data_out_OBUF_107_inst : OBUF
 port map (
   I => data_out_OBUF_107,
   O => data_out_107
);
data_out_OBUF_108_inst : OBUF
 port map (
   I => data_out_OBUF_108,
   O => data_out_108
);
data_out_OBUF_109_inst : OBUF
 port map (
   I => data_out_OBUF_109,
   O => data_out_109
);
data_out_OBUF_10_inst : OBUF
 port map (
   I => data_out_OBUF_10,
   O => data_out_10
);
data_out_OBUF_110_inst : OBUF
 port map (
   I => data_out_OBUF_110,
   O => data_out_110
);
data_out_OBUF_111_inst : OBUF
 port map (
   I => data_out_OBUF_111,
   O => data_out_111
);
data_out_OBUF_112_inst : OBUF
 port map (
   I => data_out_OBUF_112,
   O => data_out_112
);
data_out_OBUF_113_inst : OBUF
 port map (
   I => data_out_OBUF_113,
   O => data_out_113
);
data_out_OBUF_114_inst : OBUF
 port map (
   I => data_out_OBUF_114,
   O => data_out_114
);
data_out_OBUF_115_inst : OBUF
 port map (
   I => data_out_OBUF_115,
   O => data_out_115
);
data_out_OBUF_116_inst : OBUF
 port map (
   I => data_out_OBUF_116,
   O => data_out_116
);
data_out_OBUF_117_inst : OBUF
 port map (
   I => data_out_OBUF_117,
   O => data_out_117
);
data_out_OBUF_118_inst : OBUF
 port map (
   I => data_out_OBUF_118,
   O => data_out_118
);
data_out_OBUF_119_inst : OBUF
 port map (
   I => data_out_OBUF_119,
   O => data_out_119
);
data_out_OBUF_11_inst : OBUF
 port map (
   I => data_out_OBUF_11,
   O => data_out_11
);
data_out_OBUF_120_inst : OBUF
 port map (
   I => data_out_OBUF_120,
   O => data_out_120
);
data_out_OBUF_121_inst : OBUF
 port map (
   I => data_out_OBUF_121,
   O => data_out_121
);
data_out_OBUF_122_inst : OBUF
 port map (
   I => data_out_OBUF_122,
   O => data_out_122
);
data_out_OBUF_123_inst : OBUF
 port map (
   I => data_out_OBUF_123,
   O => data_out_123
);
data_out_OBUF_124_inst : OBUF
 port map (
   I => data_out_OBUF_124,
   O => data_out_124
);
data_out_OBUF_125_inst : OBUF
 port map (
   I => data_out_OBUF_125,
   O => data_out_125
);
data_out_OBUF_126_inst : OBUF
 port map (
   I => data_out_OBUF_126,
   O => data_out_126
);
data_out_OBUF_127_inst : OBUF
 port map (
   I => data_out_OBUF_127,
   O => data_out_127
);
data_out_OBUF_128_inst : OBUF
 port map (
   I => data_out_OBUF_128,
   O => data_out_128
);
data_out_OBUF_129_inst : OBUF
 port map (
   I => data_out_OBUF_129,
   O => data_out_129
);
data_out_OBUF_12_inst : OBUF
 port map (
   I => data_out_OBUF_12,
   O => data_out_12
);
data_out_OBUF_130_inst : OBUF
 port map (
   I => data_out_OBUF_130,
   O => data_out_130
);
data_out_OBUF_131_inst : OBUF
 port map (
   I => data_out_OBUF_131,
   O => data_out_131
);
data_out_OBUF_132_inst : OBUF
 port map (
   I => data_out_OBUF_132,
   O => data_out_132
);
data_out_OBUF_133_inst : OBUF
 port map (
   I => data_out_OBUF_133,
   O => data_out_133
);
data_out_OBUF_134_inst : OBUF
 port map (
   I => data_out_OBUF_134,
   O => data_out_134
);
data_out_OBUF_135_inst : OBUF
 port map (
   I => data_out_OBUF_135,
   O => data_out_135
);
data_out_OBUF_136_inst : OBUF
 port map (
   I => data_out_OBUF_136,
   O => data_out_136
);
data_out_OBUF_137_inst : OBUF
 port map (
   I => data_out_OBUF_137,
   O => data_out_137
);
data_out_OBUF_138_inst : OBUF
 port map (
   I => data_out_OBUF_138,
   O => data_out_138
);
data_out_OBUF_139_inst : OBUF
 port map (
   I => data_out_OBUF_139,
   O => data_out_139
);
data_out_OBUF_13_inst : OBUF
 port map (
   I => data_out_OBUF_13,
   O => data_out_13
);
data_out_OBUF_140_inst : OBUF
 port map (
   I => data_out_OBUF_140,
   O => data_out_140
);
data_out_OBUF_141_inst : OBUF
 port map (
   I => data_out_OBUF_141,
   O => data_out_141
);
data_out_OBUF_142_inst : OBUF
 port map (
   I => data_out_OBUF_142,
   O => data_out_142
);
data_out_OBUF_143_inst : OBUF
 port map (
   I => data_out_OBUF_143,
   O => data_out_143
);
data_out_OBUF_144_inst : OBUF
 port map (
   I => data_out_OBUF_144,
   O => data_out_144
);
data_out_OBUF_145_inst : OBUF
 port map (
   I => data_out_OBUF_145,
   O => data_out_145
);
data_out_OBUF_146_inst : OBUF
 port map (
   I => data_out_OBUF_146,
   O => data_out_146
);
data_out_OBUF_147_inst : OBUF
 port map (
   I => data_out_OBUF_147,
   O => data_out_147
);
data_out_OBUF_148_inst : OBUF
 port map (
   I => data_out_OBUF_148,
   O => data_out_148
);
data_out_OBUF_149_inst : OBUF
 port map (
   I => data_out_OBUF_149,
   O => data_out_149
);
data_out_OBUF_14_inst : OBUF
 port map (
   I => data_out_OBUF_14,
   O => data_out_14
);
data_out_OBUF_150_inst : OBUF
 port map (
   I => data_out_OBUF_150,
   O => data_out_150
);
data_out_OBUF_151_inst : OBUF
 port map (
   I => data_out_OBUF_151,
   O => data_out_151
);
data_out_OBUF_152_inst : OBUF
 port map (
   I => data_out_OBUF_152,
   O => data_out_152
);
data_out_OBUF_153_inst : OBUF
 port map (
   I => data_out_OBUF_153,
   O => data_out_153
);
data_out_OBUF_154_inst : OBUF
 port map (
   I => data_out_OBUF_154,
   O => data_out_154
);
data_out_OBUF_155_inst : OBUF
 port map (
   I => data_out_OBUF_155,
   O => data_out_155
);
data_out_OBUF_156_inst : OBUF
 port map (
   I => data_out_OBUF_156,
   O => data_out_156
);
data_out_OBUF_157_inst : OBUF
 port map (
   I => data_out_OBUF_157,
   O => data_out_157
);
data_out_OBUF_158_inst : OBUF
 port map (
   I => data_out_OBUF_158,
   O => data_out_158
);
data_out_OBUF_159_inst : OBUF
 port map (
   I => data_out_OBUF_159,
   O => data_out_159
);
data_out_OBUF_15_inst : OBUF
 port map (
   I => data_out_OBUF_15,
   O => data_out_15
);
data_out_OBUF_160_inst : OBUF
 port map (
   I => data_out_OBUF_160,
   O => data_out_160
);
data_out_OBUF_161_inst : OBUF
 port map (
   I => data_out_OBUF_161,
   O => data_out_161
);
data_out_OBUF_162_inst : OBUF
 port map (
   I => data_out_OBUF_162,
   O => data_out_162
);
data_out_OBUF_163_inst : OBUF
 port map (
   I => data_out_OBUF_163,
   O => data_out_163
);
data_out_OBUF_164_inst : OBUF
 port map (
   I => data_out_OBUF_164,
   O => data_out_164
);
data_out_OBUF_165_inst : OBUF
 port map (
   I => data_out_OBUF_165,
   O => data_out_165
);
data_out_OBUF_166_inst : OBUF
 port map (
   I => data_out_OBUF_166,
   O => data_out_166
);
data_out_OBUF_167_inst : OBUF
 port map (
   I => data_out_OBUF_167,
   O => data_out_167
);
data_out_OBUF_168_inst : OBUF
 port map (
   I => data_out_OBUF_168,
   O => data_out_168
);
data_out_OBUF_169_inst : OBUF
 port map (
   I => data_out_OBUF_169,
   O => data_out_169
);
data_out_OBUF_16_inst : OBUF
 port map (
   I => data_out_OBUF_16,
   O => data_out_16
);
data_out_OBUF_170_inst : OBUF
 port map (
   I => data_out_OBUF_170,
   O => data_out_170
);
data_out_OBUF_171_inst : OBUF
 port map (
   I => data_out_OBUF_171,
   O => data_out_171
);
data_out_OBUF_172_inst : OBUF
 port map (
   I => data_out_OBUF_172,
   O => data_out_172
);
data_out_OBUF_173_inst : OBUF
 port map (
   I => data_out_OBUF_173,
   O => data_out_173
);
data_out_OBUF_174_inst : OBUF
 port map (
   I => data_out_OBUF_174,
   O => data_out_174
);
data_out_OBUF_175_inst : OBUF
 port map (
   I => data_out_OBUF_175,
   O => data_out_175
);
data_out_OBUF_176_inst : OBUF
 port map (
   I => data_out_OBUF_176,
   O => data_out_176
);
data_out_OBUF_177_inst : OBUF
 port map (
   I => data_out_OBUF_177,
   O => data_out_177
);
data_out_OBUF_178_inst : OBUF
 port map (
   I => data_out_OBUF_178,
   O => data_out_178
);
data_out_OBUF_179_inst : OBUF
 port map (
   I => data_out_OBUF_179,
   O => data_out_179
);
data_out_OBUF_17_inst : OBUF
 port map (
   I => data_out_OBUF_17,
   O => data_out_17
);
data_out_OBUF_180_inst : OBUF
 port map (
   I => data_out_OBUF_180,
   O => data_out_180
);
data_out_OBUF_181_inst : OBUF
 port map (
   I => data_out_OBUF_181,
   O => data_out_181
);
data_out_OBUF_182_inst : OBUF
 port map (
   I => data_out_OBUF_182,
   O => data_out_182
);
data_out_OBUF_183_inst : OBUF
 port map (
   I => data_out_OBUF_183,
   O => data_out_183
);
data_out_OBUF_184_inst : OBUF
 port map (
   I => data_out_OBUF_184,
   O => data_out_184
);
data_out_OBUF_185_inst : OBUF
 port map (
   I => data_out_OBUF_185,
   O => data_out_185
);
data_out_OBUF_186_inst : OBUF
 port map (
   I => data_out_OBUF_186,
   O => data_out_186
);
data_out_OBUF_187_inst : OBUF
 port map (
   I => data_out_OBUF_187,
   O => data_out_187
);
data_out_OBUF_188_inst : OBUF
 port map (
   I => data_out_OBUF_188,
   O => data_out_188
);
data_out_OBUF_189_inst : OBUF
 port map (
   I => data_out_OBUF_189,
   O => data_out_189
);
data_out_OBUF_18_inst : OBUF
 port map (
   I => data_out_OBUF_18,
   O => data_out_18
);
data_out_OBUF_190_inst : OBUF
 port map (
   I => data_out_OBUF_190,
   O => data_out_190
);
data_out_OBUF_191_inst : OBUF
 port map (
   I => data_out_OBUF_191,
   O => data_out_191
);
data_out_OBUF_192_inst : OBUF
 port map (
   I => data_out_OBUF_192,
   O => data_out_192
);
data_out_OBUF_193_inst : OBUF
 port map (
   I => data_out_OBUF_193,
   O => data_out_193
);
data_out_OBUF_194_inst : OBUF
 port map (
   I => data_out_OBUF_194,
   O => data_out_194
);
data_out_OBUF_195_inst : OBUF
 port map (
   I => data_out_OBUF_195,
   O => data_out_195
);
data_out_OBUF_196_inst : OBUF
 port map (
   I => data_out_OBUF_196,
   O => data_out_196
);
data_out_OBUF_197_inst : OBUF
 port map (
   I => data_out_OBUF_197,
   O => data_out_197
);
data_out_OBUF_198_inst : OBUF
 port map (
   I => data_out_OBUF_198,
   O => data_out_198
);
data_out_OBUF_199_inst : OBUF
 port map (
   I => data_out_OBUF_199,
   O => data_out_199
);
data_out_OBUF_19_inst : OBUF
 port map (
   I => data_out_OBUF_19,
   O => data_out_19
);
data_out_OBUF_1_inst : OBUF
 port map (
   I => data_out_OBUF_1,
   O => data_out_1
);
data_out_OBUF_200_inst : OBUF
 port map (
   I => data_out_OBUF_200,
   O => data_out_200
);
data_out_OBUF_201_inst : OBUF
 port map (
   I => data_out_OBUF_201,
   O => data_out_201
);
data_out_OBUF_202_inst : OBUF
 port map (
   I => data_out_OBUF_202,
   O => data_out_202
);
data_out_OBUF_203_inst : OBUF
 port map (
   I => data_out_OBUF_203,
   O => data_out_203
);
data_out_OBUF_204_inst : OBUF
 port map (
   I => data_out_OBUF_204,
   O => data_out_204
);
data_out_OBUF_205_inst : OBUF
 port map (
   I => data_out_OBUF_205,
   O => data_out_205
);
data_out_OBUF_206_inst : OBUF
 port map (
   I => data_out_OBUF_206,
   O => data_out_206
);
data_out_OBUF_207_inst : OBUF
 port map (
   I => data_out_OBUF_207,
   O => data_out_207
);
data_out_OBUF_208_inst : OBUF
 port map (
   I => data_out_OBUF_208,
   O => data_out_208
);
data_out_OBUF_209_inst : OBUF
 port map (
   I => data_out_OBUF_209,
   O => data_out_209
);
data_out_OBUF_20_inst : OBUF
 port map (
   I => data_out_OBUF_20,
   O => data_out_20
);
data_out_OBUF_210_inst : OBUF
 port map (
   I => data_out_OBUF_210,
   O => data_out_210
);
data_out_OBUF_211_inst : OBUF
 port map (
   I => data_out_OBUF_211,
   O => data_out_211
);
data_out_OBUF_212_inst : OBUF
 port map (
   I => data_out_OBUF_212,
   O => data_out_212
);
data_out_OBUF_213_inst : OBUF
 port map (
   I => data_out_OBUF_213,
   O => data_out_213
);
data_out_OBUF_214_inst : OBUF
 port map (
   I => data_out_OBUF_214,
   O => data_out_214
);
data_out_OBUF_215_inst : OBUF
 port map (
   I => data_out_OBUF_215,
   O => data_out_215
);
data_out_OBUF_216_inst : OBUF
 port map (
   I => data_out_OBUF_216,
   O => data_out_216
);
data_out_OBUF_217_inst : OBUF
 port map (
   I => data_out_OBUF_217,
   O => data_out_217
);
data_out_OBUF_218_inst : OBUF
 port map (
   I => data_out_OBUF_218,
   O => data_out_218
);
data_out_OBUF_219_inst : OBUF
 port map (
   I => data_out_OBUF_219,
   O => data_out_219
);
data_out_OBUF_21_inst : OBUF
 port map (
   I => data_out_OBUF_21,
   O => data_out_21
);
data_out_OBUF_220_inst : OBUF
 port map (
   I => data_out_OBUF_220,
   O => data_out_220
);
data_out_OBUF_221_inst : OBUF
 port map (
   I => data_out_OBUF_221,
   O => data_out_221
);
data_out_OBUF_222_inst : OBUF
 port map (
   I => data_out_OBUF_222,
   O => data_out_222
);
data_out_OBUF_223_inst : OBUF
 port map (
   I => data_out_OBUF_223,
   O => data_out_223
);
data_out_OBUF_224_inst : OBUF
 port map (
   I => data_out_OBUF_224,
   O => data_out_224
);
data_out_OBUF_225_inst : OBUF
 port map (
   I => data_out_OBUF_225,
   O => data_out_225
);
data_out_OBUF_226_inst : OBUF
 port map (
   I => data_out_OBUF_226,
   O => data_out_226
);
data_out_OBUF_227_inst : OBUF
 port map (
   I => data_out_OBUF_227,
   O => data_out_227
);
data_out_OBUF_228_inst : OBUF
 port map (
   I => data_out_OBUF_228,
   O => data_out_228
);
data_out_OBUF_229_inst : OBUF
 port map (
   I => data_out_OBUF_229,
   O => data_out_229
);
data_out_OBUF_22_inst : OBUF
 port map (
   I => data_out_OBUF_22,
   O => data_out_22
);
data_out_OBUF_230_inst : OBUF
 port map (
   I => data_out_OBUF_230,
   O => data_out_230
);
data_out_OBUF_231_inst : OBUF
 port map (
   I => data_out_OBUF_231,
   O => data_out_231
);
data_out_OBUF_232_inst : OBUF
 port map (
   I => data_out_OBUF_232,
   O => data_out_232
);
data_out_OBUF_233_inst : OBUF
 port map (
   I => data_out_OBUF_233,
   O => data_out_233
);
data_out_OBUF_234_inst : OBUF
 port map (
   I => data_out_OBUF_234,
   O => data_out_234
);
data_out_OBUF_235_inst : OBUF
 port map (
   I => data_out_OBUF_235,
   O => data_out_235
);
data_out_OBUF_236_inst : OBUF
 port map (
   I => data_out_OBUF_236,
   O => data_out_236
);
data_out_OBUF_237_inst : OBUF
 port map (
   I => data_out_OBUF_237,
   O => data_out_237
);
data_out_OBUF_238_inst : OBUF
 port map (
   I => data_out_OBUF_238,
   O => data_out_238
);
data_out_OBUF_239_inst : OBUF
 port map (
   I => data_out_OBUF_239,
   O => data_out_239
);
data_out_OBUF_23_inst : OBUF
 port map (
   I => data_out_OBUF_23,
   O => data_out_23
);
data_out_OBUF_240_inst : OBUF
 port map (
   I => data_out_OBUF_240,
   O => data_out_240
);
data_out_OBUF_241_inst : OBUF
 port map (
   I => data_out_OBUF_241,
   O => data_out_241
);
data_out_OBUF_242_inst : OBUF
 port map (
   I => data_out_OBUF_242,
   O => data_out_242
);
data_out_OBUF_243_inst : OBUF
 port map (
   I => data_out_OBUF_243,
   O => data_out_243
);
data_out_OBUF_244_inst : OBUF
 port map (
   I => data_out_OBUF_244,
   O => data_out_244
);
data_out_OBUF_245_inst : OBUF
 port map (
   I => data_out_OBUF_245,
   O => data_out_245
);
data_out_OBUF_246_inst : OBUF
 port map (
   I => data_out_OBUF_246,
   O => data_out_246
);
data_out_OBUF_247_inst : OBUF
 port map (
   I => data_out_OBUF_247,
   O => data_out_247
);
data_out_OBUF_248_inst : OBUF
 port map (
   I => data_out_OBUF_248,
   O => data_out_248
);
data_out_OBUF_249_inst : OBUF
 port map (
   I => data_out_OBUF_249,
   O => data_out_249
);
data_out_OBUF_24_inst : OBUF
 port map (
   I => data_out_OBUF_24,
   O => data_out_24
);
data_out_OBUF_250_inst : OBUF
 port map (
   I => data_out_OBUF_250,
   O => data_out_250
);
data_out_OBUF_251_inst : OBUF
 port map (
   I => data_out_OBUF_251,
   O => data_out_251
);
data_out_OBUF_252_inst : OBUF
 port map (
   I => data_out_OBUF_252,
   O => data_out_252
);
data_out_OBUF_253_inst : OBUF
 port map (
   I => data_out_OBUF_253,
   O => data_out_253
);
data_out_OBUF_254_inst : OBUF
 port map (
   I => data_out_OBUF_254,
   O => data_out_254
);
data_out_OBUF_255_inst : OBUF
 port map (
   I => data_out_OBUF_255,
   O => data_out_255
);
data_out_OBUF_25_inst : OBUF
 port map (
   I => data_out_OBUF_25,
   O => data_out_25
);
data_out_OBUF_26_inst : OBUF
 port map (
   I => data_out_OBUF_26,
   O => data_out_26
);
data_out_OBUF_27_inst : OBUF
 port map (
   I => data_out_OBUF_27,
   O => data_out_27
);
data_out_OBUF_28_inst : OBUF
 port map (
   I => data_out_OBUF_28,
   O => data_out_28
);
data_out_OBUF_29_inst : OBUF
 port map (
   I => data_out_OBUF_29,
   O => data_out_29
);
data_out_OBUF_2_inst : OBUF
 port map (
   I => data_out_OBUF_2,
   O => data_out_2
);
data_out_OBUF_30_inst : OBUF
 port map (
   I => data_out_OBUF_30,
   O => data_out_30
);
data_out_OBUF_31_inst : OBUF
 port map (
   I => data_out_OBUF_31,
   O => data_out_31
);
data_out_OBUF_32_inst : OBUF
 port map (
   I => data_out_OBUF_32,
   O => data_out_32
);
data_out_OBUF_33_inst : OBUF
 port map (
   I => data_out_OBUF_33,
   O => data_out_33
);
data_out_OBUF_34_inst : OBUF
 port map (
   I => data_out_OBUF_34,
   O => data_out_34
);
data_out_OBUF_35_inst : OBUF
 port map (
   I => data_out_OBUF_35,
   O => data_out_35
);
data_out_OBUF_36_inst : OBUF
 port map (
   I => data_out_OBUF_36,
   O => data_out_36
);
data_out_OBUF_37_inst : OBUF
 port map (
   I => data_out_OBUF_37,
   O => data_out_37
);
data_out_OBUF_38_inst : OBUF
 port map (
   I => data_out_OBUF_38,
   O => data_out_38
);
data_out_OBUF_39_inst : OBUF
 port map (
   I => data_out_OBUF_39,
   O => data_out_39
);
data_out_OBUF_3_inst : OBUF
 port map (
   I => data_out_OBUF_3,
   O => data_out_3
);
data_out_OBUF_40_inst : OBUF
 port map (
   I => data_out_OBUF_40,
   O => data_out_40
);
data_out_OBUF_41_inst : OBUF
 port map (
   I => data_out_OBUF_41,
   O => data_out_41
);
data_out_OBUF_42_inst : OBUF
 port map (
   I => data_out_OBUF_42,
   O => data_out_42
);
data_out_OBUF_43_inst : OBUF
 port map (
   I => data_out_OBUF_43,
   O => data_out_43
);
data_out_OBUF_44_inst : OBUF
 port map (
   I => data_out_OBUF_44,
   O => data_out_44
);
data_out_OBUF_45_inst : OBUF
 port map (
   I => data_out_OBUF_45,
   O => data_out_45
);
data_out_OBUF_46_inst : OBUF
 port map (
   I => data_out_OBUF_46,
   O => data_out_46
);
data_out_OBUF_47_inst : OBUF
 port map (
   I => data_out_OBUF_47,
   O => data_out_47
);
data_out_OBUF_48_inst : OBUF
 port map (
   I => data_out_OBUF_48,
   O => data_out_48
);
data_out_OBUF_49_inst : OBUF
 port map (
   I => data_out_OBUF_49,
   O => data_out_49
);
data_out_OBUF_4_inst : OBUF
 port map (
   I => data_out_OBUF_4,
   O => data_out_4
);
data_out_OBUF_50_inst : OBUF
 port map (
   I => data_out_OBUF_50,
   O => data_out_50
);
data_out_OBUF_51_inst : OBUF
 port map (
   I => data_out_OBUF_51,
   O => data_out_51
);
data_out_OBUF_52_inst : OBUF
 port map (
   I => data_out_OBUF_52,
   O => data_out_52
);
data_out_OBUF_53_inst : OBUF
 port map (
   I => data_out_OBUF_53,
   O => data_out_53
);
data_out_OBUF_54_inst : OBUF
 port map (
   I => data_out_OBUF_54,
   O => data_out_54
);
data_out_OBUF_55_inst : OBUF
 port map (
   I => data_out_OBUF_55,
   O => data_out_55
);
data_out_OBUF_56_inst : OBUF
 port map (
   I => data_out_OBUF_56,
   O => data_out_56
);
data_out_OBUF_57_inst : OBUF
 port map (
   I => data_out_OBUF_57,
   O => data_out_57
);
data_out_OBUF_58_inst : OBUF
 port map (
   I => data_out_OBUF_58,
   O => data_out_58
);
data_out_OBUF_59_inst : OBUF
 port map (
   I => data_out_OBUF_59,
   O => data_out_59
);
data_out_OBUF_5_inst : OBUF
 port map (
   I => data_out_OBUF_5,
   O => data_out_5
);
data_out_OBUF_60_inst : OBUF
 port map (
   I => data_out_OBUF_60,
   O => data_out_60
);
data_out_OBUF_61_inst : OBUF
 port map (
   I => data_out_OBUF_61,
   O => data_out_61
);
data_out_OBUF_62_inst : OBUF
 port map (
   I => data_out_OBUF_62,
   O => data_out_62
);
data_out_OBUF_63_inst : OBUF
 port map (
   I => data_out_OBUF_63,
   O => data_out_63
);
data_out_OBUF_64_inst : OBUF
 port map (
   I => data_out_OBUF_64,
   O => data_out_64
);
data_out_OBUF_65_inst : OBUF
 port map (
   I => data_out_OBUF_65,
   O => data_out_65
);
data_out_OBUF_66_inst : OBUF
 port map (
   I => data_out_OBUF_66,
   O => data_out_66
);
data_out_OBUF_67_inst : OBUF
 port map (
   I => data_out_OBUF_67,
   O => data_out_67
);
data_out_OBUF_68_inst : OBUF
 port map (
   I => data_out_OBUF_68,
   O => data_out_68
);
data_out_OBUF_69_inst : OBUF
 port map (
   I => data_out_OBUF_69,
   O => data_out_69
);
data_out_OBUF_6_inst : OBUF
 port map (
   I => data_out_OBUF_6,
   O => data_out_6
);
data_out_OBUF_70_inst : OBUF
 port map (
   I => data_out_OBUF_70,
   O => data_out_70
);
data_out_OBUF_71_inst : OBUF
 port map (
   I => data_out_OBUF_71,
   O => data_out_71
);
data_out_OBUF_72_inst : OBUF
 port map (
   I => data_out_OBUF_72,
   O => data_out_72
);
data_out_OBUF_73_inst : OBUF
 port map (
   I => data_out_OBUF_73,
   O => data_out_73
);
data_out_OBUF_74_inst : OBUF
 port map (
   I => data_out_OBUF_74,
   O => data_out_74
);
data_out_OBUF_75_inst : OBUF
 port map (
   I => data_out_OBUF_75,
   O => data_out_75
);
data_out_OBUF_76_inst : OBUF
 port map (
   I => data_out_OBUF_76,
   O => data_out_76
);
data_out_OBUF_77_inst : OBUF
 port map (
   I => data_out_OBUF_77,
   O => data_out_77
);
data_out_OBUF_78_inst : OBUF
 port map (
   I => data_out_OBUF_78,
   O => data_out_78
);
data_out_OBUF_79_inst : OBUF
 port map (
   I => data_out_OBUF_79,
   O => data_out_79
);
data_out_OBUF_7_inst : OBUF
 port map (
   I => data_out_OBUF_7,
   O => data_out_7
);
data_out_OBUF_80_inst : OBUF
 port map (
   I => data_out_OBUF_80,
   O => data_out_80
);
data_out_OBUF_81_inst : OBUF
 port map (
   I => data_out_OBUF_81,
   O => data_out_81
);
data_out_OBUF_82_inst : OBUF
 port map (
   I => data_out_OBUF_82,
   O => data_out_82
);
data_out_OBUF_83_inst : OBUF
 port map (
   I => data_out_OBUF_83,
   O => data_out_83
);
data_out_OBUF_84_inst : OBUF
 port map (
   I => data_out_OBUF_84,
   O => data_out_84
);
data_out_OBUF_85_inst : OBUF
 port map (
   I => data_out_OBUF_85,
   O => data_out_85
);
data_out_OBUF_86_inst : OBUF
 port map (
   I => data_out_OBUF_86,
   O => data_out_86
);
data_out_OBUF_87_inst : OBUF
 port map (
   I => data_out_OBUF_87,
   O => data_out_87
);
data_out_OBUF_88_inst : OBUF
 port map (
   I => data_out_OBUF_88,
   O => data_out_88
);
data_out_OBUF_89_inst : OBUF
 port map (
   I => data_out_OBUF_89,
   O => data_out_89
);
data_out_OBUF_8_inst : OBUF
 port map (
   I => data_out_OBUF_8,
   O => data_out_8
);
data_out_OBUF_90_inst : OBUF
 port map (
   I => data_out_OBUF_90,
   O => data_out_90
);
data_out_OBUF_91_inst : OBUF
 port map (
   I => data_out_OBUF_91,
   O => data_out_91
);
data_out_OBUF_92_inst : OBUF
 port map (
   I => data_out_OBUF_92,
   O => data_out_92
);
data_out_OBUF_93_inst : OBUF
 port map (
   I => data_out_OBUF_93,
   O => data_out_93
);
data_out_OBUF_94_inst : OBUF
 port map (
   I => data_out_OBUF_94,
   O => data_out_94
);
data_out_OBUF_95_inst : OBUF
 port map (
   I => data_out_OBUF_95,
   O => data_out_95
);
data_out_OBUF_96_inst : OBUF
 port map (
   I => data_out_OBUF_96,
   O => data_out_96
);
data_out_OBUF_97_inst : OBUF
 port map (
   I => data_out_OBUF_97,
   O => data_out_97
);
data_out_OBUF_98_inst : OBUF
 port map (
   I => data_out_OBUF_98,
   O => data_out_98
);
data_out_OBUF_99_inst : OBUF
 port map (
   I => data_out_OBUF_99,
   O => data_out_99
);
data_out_OBUF_9_inst : OBUF
 port map (
   I => data_out_OBUF_9,
   O => data_out_9
);
data_ready_IBUF_inst : IBUF
 port map (
   I => data_ready,
   O => data_ready_IBUF
);
d_0_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => c_reg_n_0_0,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_128,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => d_0_i_1_n_0
);
d_10_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => c_reg_n_0_10,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_138,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => d_10_i_1_n_0
);
d_11_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => c_reg_n_0_11,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_139,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => d_11_i_1_n_0
);
d_12_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => c_reg_n_0_12,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_140,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => d_12_i_1_n_0
);
d_13_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => c_reg_n_0_13,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_141,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => d_13_i_1_n_0
);
d_14_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => c_reg_n_0_14,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_142,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => d_14_i_1_n_0
);
d_15_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => c_reg_n_0_15,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_143,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => d_15_i_1_n_0
);
d_16_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => c_reg_n_0_16,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_144,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => d_16_i_1_n_0
);
d_17_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => c_reg_n_0_17,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_145,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => d_17_i_1_n_0
);
d_18_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => c_reg_n_0_18,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_146,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => d_18_i_1_n_0
);
d_19_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => c_reg_n_0_19,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_147,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => d_19_i_1_n_0
);
d_1_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => c_reg_n_0_1,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_129,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => d_1_i_1_n_0
);
d_20_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => c_reg_n_0_20,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_148,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => d_20_i_1_n_0
);
d_21_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => c_reg_n_0_21,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_149,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => d_21_i_1_n_0
);
d_22_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => c_reg_n_0_22,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_150,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => d_22_i_1_n_0
);
d_23_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => c_reg_n_0_23,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_151,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => d_23_i_1_n_0
);
d_24_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => c_reg_n_0_24,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_152,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => d_24_i_1_n_0
);
d_25_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => c_reg_n_0_25,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_153,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => d_25_i_1_n_0
);
d_26_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => c_reg_n_0_26,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_154,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => d_26_i_1_n_0
);
d_27_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => c_reg_n_0_27,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_155,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => d_27_i_1_n_0
);
d_28_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => c_reg_n_0_28,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_156,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => d_28_i_1_n_0
);
d_29_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => c_reg_n_0_29,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_157,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => d_29_i_1_n_0
);
d_2_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => c_reg_n_0_2,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_130,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => d_2_i_1_n_0
);
d_30_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => c_reg_n_0_30,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_158,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => d_30_i_1_n_0
);
d_31_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => c_reg_n_0_31,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_159,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => d_31_i_1_n_0
);
d_3_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => c_reg_n_0_3,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_131,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => d_3_i_1_n_0
);
d_4_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => c_reg_n_0_4,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_132,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => d_4_i_1_n_0
);
d_5_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => c_reg_n_0_5,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_133,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => d_5_i_1_n_0
);
d_6_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => c_reg_n_0_6,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_134,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => d_6_i_1_n_0
);
d_7_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => c_reg_n_0_7,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_135,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => d_7_i_1_n_0
);
d_8_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => c_reg_n_0_8,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_136,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => d_8_i_1_n_0
);
d_9_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => c_reg_n_0_9,
   I1 => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0,
   I2 => data_out_OBUF_137,
   I3 => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0,
   O => d_9_i_1_n_0
);
d_reg_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => d_0_i_1_n_0,
   R => '0',
   Q => d_0
);
d_reg_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => d_10_i_1_n_0,
   R => '0',
   Q => d_10
);
d_reg_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => d_11_i_1_n_0,
   R => '0',
   Q => d_11
);
d_reg_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => d_12_i_1_n_0,
   R => '0',
   Q => d_12
);
d_reg_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => d_13_i_1_n_0,
   R => '0',
   Q => d_13
);
d_reg_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => d_14_i_1_n_0,
   R => '0',
   Q => d_14
);
d_reg_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => d_15_i_1_n_0,
   R => '0',
   Q => d_15
);
d_reg_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => d_16_i_1_n_0,
   R => '0',
   Q => d_16
);
d_reg_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => d_17_i_1_n_0,
   R => '0',
   Q => d_17
);
d_reg_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => d_18_i_1_n_0,
   R => '0',
   Q => d_18
);
d_reg_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => d_19_i_1_n_0,
   R => '0',
   Q => d_19
);
d_reg_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => d_1_i_1_n_0,
   R => '0',
   Q => d_1
);
d_reg_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => d_20_i_1_n_0,
   R => '0',
   Q => d_20
);
d_reg_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => d_21_i_1_n_0,
   R => '0',
   Q => d_21
);
d_reg_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => d_22_i_1_n_0,
   R => '0',
   Q => d_22
);
d_reg_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => d_23_i_1_n_0,
   R => '0',
   Q => d_23
);
d_reg_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => d_24_i_1_n_0,
   R => '0',
   Q => d_24
);
d_reg_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => d_25_i_1_n_0,
   R => '0',
   Q => d_25
);
d_reg_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => d_26_i_1_n_0,
   R => '0',
   Q => d_26
);
d_reg_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => d_27_i_1_n_0,
   R => '0',
   Q => d_27
);
d_reg_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => d_28_i_1_n_0,
   R => '0',
   Q => d_28
);
d_reg_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => d_29_i_1_n_0,
   R => '0',
   Q => d_29
);
d_reg_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => d_2_i_1_n_0,
   R => '0',
   Q => d_2
);
d_reg_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => d_30_i_1_n_0,
   R => '0',
   Q => d_30
);
d_reg_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => d_31_i_1_n_0,
   R => '0',
   Q => d_31
);
d_reg_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => d_3_i_1_n_0,
   R => '0',
   Q => d_3
);
d_reg_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => d_4_i_1_n_0,
   R => '0',
   Q => d_4
);
d_reg_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => d_5_i_1_n_0,
   R => '0',
   Q => d_5
);
d_reg_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => d_6_i_1_n_0,
   R => '0',
   Q => d_6
);
d_reg_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => d_7_i_1_n_0,
   R => '0',
   Q => d_7
);
d_reg_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => d_8_i_1_n_0,
   R => '0',
   Q => d_8
);
d_reg_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => d_9_i_1_n_0,
   R => '0',
   Q => d_9
);
e_0_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in15_0,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_96,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => e_0_i_1_n_0
);
e_10_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in15_10,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_106,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => e_10_i_1_n_0
);
e_11_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in15_11,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_107,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => e_11_i_1_n_0
);
e_11_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_11,
   I1 => T1_0_11,
   O => e_11_i_3_n_0
);
e_11_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_10,
   I1 => T1_0_10,
   O => e_11_i_4_n_0
);
e_11_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_9,
   I1 => T1_0_9,
   O => e_11_i_5_n_0
);
e_11_i_6 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_8,
   I1 => T1_0_8,
   O => e_11_i_6_n_0
);
e_12_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in15_12,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_108,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => e_12_i_1_n_0
);
e_13_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in15_13,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_109,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => e_13_i_1_n_0
);
e_14_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in15_14,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_110,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => e_14_i_1_n_0
);
e_15_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in15_15,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_111,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => e_15_i_1_n_0
);
e_15_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_15,
   I1 => T1_0_15,
   O => e_15_i_3_n_0
);
e_15_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_14,
   I1 => T1_0_14,
   O => e_15_i_4_n_0
);
e_15_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_13,
   I1 => T1_0_13,
   O => e_15_i_5_n_0
);
e_15_i_6 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_12,
   I1 => T1_0_12,
   O => e_15_i_6_n_0
);
e_16_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in15_16,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_112,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => e_16_i_1_n_0
);
e_17_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in15_17,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_113,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => e_17_i_1_n_0
);
e_18_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in15_18,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_114,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => e_18_i_1_n_0
);
e_19_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in15_19,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_115,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => e_19_i_1_n_0
);
e_19_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_19,
   I1 => T1_0_19,
   O => e_19_i_3_n_0
);
e_19_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_18,
   I1 => T1_0_18,
   O => e_19_i_4_n_0
);
e_19_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_17,
   I1 => T1_0_17,
   O => e_19_i_5_n_0
);
e_19_i_6 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_16,
   I1 => T1_0_16,
   O => e_19_i_6_n_0
);
e_1_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in15_1,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_97,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => e_1_i_1_n_0
);
e_20_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in15_20,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_116,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => e_20_i_1_n_0
);
e_21_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in15_21,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_117,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => e_21_i_1_n_0
);
e_22_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in15_22,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_118,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => e_22_i_1_n_0
);
e_23_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in15_23,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_119,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => e_23_i_1_n_0
);
e_23_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_23,
   I1 => T1_0_23,
   O => e_23_i_3_n_0
);
e_23_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_22,
   I1 => T1_0_22,
   O => e_23_i_4_n_0
);
e_23_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_21,
   I1 => T1_0_21,
   O => e_23_i_5_n_0
);
e_23_i_6 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_20,
   I1 => T1_0_20,
   O => e_23_i_6_n_0
);
e_24_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in15_24,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_120,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => e_24_i_1_n_0
);
e_25_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in15_25,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_121,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => e_25_i_1_n_0
);
e_26_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in15_26,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_122,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => e_26_i_1_n_0
);
e_27_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in15_27,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_123,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => e_27_i_1_n_0
);
e_27_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_27,
   I1 => T1_0_27,
   O => e_27_i_3_n_0
);
e_27_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_26,
   I1 => T1_0_26,
   O => e_27_i_4_n_0
);
e_27_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_25,
   I1 => T1_0_25,
   O => e_27_i_5_n_0
);
e_27_i_6 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_24,
   I1 => T1_0_24,
   O => e_27_i_6_n_0
);
e_28_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in15_28,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_124,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => e_28_i_1_n_0
);
e_29_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in15_29,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_125,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => e_29_i_1_n_0
);
e_2_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in15_2,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_98,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => e_2_i_1_n_0
);
e_30_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in15_30,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_126,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => e_30_i_1_n_0
);
e_31_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in15_31,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_127,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => e_31_i_1_n_0
);
e_31_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_31,
   I1 => T1_0_31,
   O => e_31_i_3_n_0
);
e_31_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_30,
   I1 => T1_0_30,
   O => e_31_i_4_n_0
);
e_31_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_29,
   I1 => T1_0_29,
   O => e_31_i_5_n_0
);
e_31_i_6 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_28,
   I1 => T1_0_28,
   O => e_31_i_6_n_0
);
e_3_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in15_3,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_99,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => e_3_i_1_n_0
);
e_3_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_3,
   I1 => T1_0_3,
   O => e_3_i_3_n_0
);
e_3_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_2,
   I1 => T1_0_2,
   O => e_3_i_4_n_0
);
e_3_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_1,
   I1 => T1_0_1,
   O => e_3_i_5_n_0
);
e_3_i_6 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_0,
   I1 => T1_0_0,
   O => e_3_i_6_n_0
);
e_4_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in15_4,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_100,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => e_4_i_1_n_0
);
e_5_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in15_5,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_101,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => e_5_i_1_n_0
);
e_6_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in15_6,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_102,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => e_6_i_1_n_0
);
e_7_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in15_7,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_103,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => e_7_i_1_n_0
);
e_7_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_7,
   I1 => T1_0_7,
   O => e_7_i_3_n_0
);
e_7_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_6,
   I1 => T1_0_6,
   O => e_7_i_4_n_0
);
e_7_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_5,
   I1 => T1_0_5,
   O => e_7_i_5_n_0
);
e_7_i_6 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_4,
   I1 => T1_0_4,
   O => e_7_i_6_n_0
);
e_8_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in15_8,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_104,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => e_8_i_1_n_0
);
e_9_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => in15_9,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_105,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => e_9_i_1_n_0
);
e_reg_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => e_0_i_1_n_0,
   R => '0',
   Q => ROTR11_out_11
);
e_reg_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => e_10_i_1_n_0,
   R => '0',
   Q => ROTR11_out_1
);
e_reg_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => e_11_i_1_n_0,
   R => '0',
   Q => ROTR11_out_32
);
e_reg_11_i_2 : CARRY4
 port map (
   CI => e_reg_7_i_2_n_0,
   CYINIT => '0',
   DI(0) => d_8,
   DI(1) => d_9,
   DI(2) => d_10,
   DI(3) => d_11,
   S(0) => e_11_i_6_n_0,
   S(1) => e_11_i_5_n_0,
   S(2) => e_11_i_4_n_0,
   S(3) => e_11_i_3_n_0,
   CO(0) => e_reg_11_i_2_n_3,
   CO(1) => e_reg_11_i_2_n_2,
   CO(2) => e_reg_11_i_2_n_1,
   CO(3) => e_reg_11_i_2_n_0,
   O(0) => in15_8,
   O(1) => in15_9,
   O(2) => in15_10,
   O(3) => in15_11
);
e_reg_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => e_12_i_1_n_0,
   R => '0',
   Q => ROTR11_out_31
);
e_reg_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => e_13_i_1_n_0,
   R => '0',
   Q => ROTR11_out_30
);
e_reg_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => e_14_i_1_n_0,
   R => '0',
   Q => ROTR11_out_29
);
e_reg_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => e_15_i_1_n_0,
   R => '0',
   Q => ROTR11_out_28
);
e_reg_15_i_2 : CARRY4
 port map (
   CI => e_reg_11_i_2_n_0,
   CYINIT => '0',
   DI(0) => d_12,
   DI(1) => d_13,
   DI(2) => d_14,
   DI(3) => d_15,
   S(0) => e_15_i_6_n_0,
   S(1) => e_15_i_5_n_0,
   S(2) => e_15_i_4_n_0,
   S(3) => e_15_i_3_n_0,
   CO(0) => e_reg_15_i_2_n_3,
   CO(1) => e_reg_15_i_2_n_2,
   CO(2) => e_reg_15_i_2_n_1,
   CO(3) => e_reg_15_i_2_n_0,
   O(0) => in15_12,
   O(1) => in15_13,
   O(2) => in15_14,
   O(3) => in15_15
);
e_reg_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => e_16_i_1_n_0,
   R => '0',
   Q => ROTR11_out_27
);
e_reg_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => e_17_i_1_n_0,
   R => '0',
   Q => ROTR11_out_26
);
e_reg_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => e_18_i_1_n_0,
   R => '0',
   Q => ROTR11_out_25
);
e_reg_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => e_19_i_1_n_0,
   R => '0',
   Q => ROTR11_out_24
);
e_reg_19_i_2 : CARRY4
 port map (
   CI => e_reg_15_i_2_n_0,
   CYINIT => '0',
   DI(0) => d_16,
   DI(1) => d_17,
   DI(2) => d_18,
   DI(3) => d_19,
   S(0) => e_19_i_6_n_0,
   S(1) => e_19_i_5_n_0,
   S(2) => e_19_i_4_n_0,
   S(3) => e_19_i_3_n_0,
   CO(0) => e_reg_19_i_2_n_3,
   CO(1) => e_reg_19_i_2_n_2,
   CO(2) => e_reg_19_i_2_n_1,
   CO(3) => e_reg_19_i_2_n_0,
   O(0) => in15_16,
   O(1) => in15_17,
   O(2) => in15_18,
   O(3) => in15_19
);
e_reg_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => e_1_i_1_n_0,
   R => '0',
   Q => ROTR11_out_10
);
e_reg_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => e_20_i_1_n_0,
   R => '0',
   Q => ROTR11_out_23
);
e_reg_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => e_21_i_1_n_0,
   R => '0',
   Q => ROTR11_out_22
);
e_reg_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => e_22_i_1_n_0,
   R => '0',
   Q => ROTR11_out_21
);
e_reg_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => e_23_i_1_n_0,
   R => '0',
   Q => ROTR11_out_20
);
e_reg_23_i_2 : CARRY4
 port map (
   CI => e_reg_19_i_2_n_0,
   CYINIT => '0',
   DI(0) => d_20,
   DI(1) => d_21,
   DI(2) => d_22,
   DI(3) => d_23,
   S(0) => e_23_i_6_n_0,
   S(1) => e_23_i_5_n_0,
   S(2) => e_23_i_4_n_0,
   S(3) => e_23_i_3_n_0,
   CO(0) => e_reg_23_i_2_n_3,
   CO(1) => e_reg_23_i_2_n_2,
   CO(2) => e_reg_23_i_2_n_1,
   CO(3) => e_reg_23_i_2_n_0,
   O(0) => in15_20,
   O(1) => in15_21,
   O(2) => in15_22,
   O(3) => in15_23
);
e_reg_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => e_24_i_1_n_0,
   R => '0',
   Q => ROTR11_out_19
);
e_reg_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => e_25_i_1_n_0,
   R => '0',
   Q => ROTR11_out_18
);
e_reg_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => e_26_i_1_n_0,
   R => '0',
   Q => ROTR11_out_17
);
e_reg_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => e_27_i_1_n_0,
   R => '0',
   Q => ROTR11_out_16
);
e_reg_27_i_2 : CARRY4
 port map (
   CI => e_reg_23_i_2_n_0,
   CYINIT => '0',
   DI(0) => d_24,
   DI(1) => d_25,
   DI(2) => d_26,
   DI(3) => d_27,
   S(0) => e_27_i_6_n_0,
   S(1) => e_27_i_5_n_0,
   S(2) => e_27_i_4_n_0,
   S(3) => e_27_i_3_n_0,
   CO(0) => e_reg_27_i_2_n_3,
   CO(1) => e_reg_27_i_2_n_2,
   CO(2) => e_reg_27_i_2_n_1,
   CO(3) => e_reg_27_i_2_n_0,
   O(0) => in15_24,
   O(1) => in15_25,
   O(2) => in15_26,
   O(3) => in15_27
);
e_reg_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => e_28_i_1_n_0,
   R => '0',
   Q => ROTR11_out_15
);
e_reg_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => e_29_i_1_n_0,
   R => '0',
   Q => ROTR11_out_14
);
e_reg_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => e_2_i_1_n_0,
   R => '0',
   Q => ROTR11_out_9
);
e_reg_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => e_30_i_1_n_0,
   R => '0',
   Q => ROTR11_out_13
);
e_reg_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => e_31_i_1_n_0,
   R => '0',
   Q => ROTR11_out_12
);
e_reg_31_i_2 : CARRY4
 port map (
   CI => e_reg_27_i_2_n_0,
   CYINIT => '0',
   DI(0) => d_28,
   DI(1) => d_29,
   DI(2) => d_30,
   DI(3) => '0',
   S(0) => e_31_i_6_n_0,
   S(1) => e_31_i_5_n_0,
   S(2) => e_31_i_4_n_0,
   S(3) => e_31_i_3_n_0,
   CO(0) => e_reg_31_i_2_n_3,
   CO(1) => e_reg_31_i_2_n_2,
   CO(2) => e_reg_31_i_2_n_1,
   CO(3) => NLW_e_reg_31_i_2_CO_UNCONNECTED_3,
   O(0) => in15_28,
   O(1) => in15_29,
   O(2) => in15_30,
   O(3) => in15_31
);
e_reg_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => e_3_i_1_n_0,
   R => '0',
   Q => ROTR11_out_8
);
e_reg_3_i_2 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => d_0,
   DI(1) => d_1,
   DI(2) => d_2,
   DI(3) => d_3,
   S(0) => e_3_i_6_n_0,
   S(1) => e_3_i_5_n_0,
   S(2) => e_3_i_4_n_0,
   S(3) => e_3_i_3_n_0,
   CO(0) => e_reg_3_i_2_n_3,
   CO(1) => e_reg_3_i_2_n_2,
   CO(2) => e_reg_3_i_2_n_1,
   CO(3) => e_reg_3_i_2_n_0,
   O(0) => in15_0,
   O(1) => in15_1,
   O(2) => in15_2,
   O(3) => in15_3
);
e_reg_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => e_4_i_1_n_0,
   R => '0',
   Q => ROTR11_out_7
);
e_reg_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => e_5_i_1_n_0,
   R => '0',
   Q => ROTR11_out_6
);
e_reg_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => e_6_i_1_n_0,
   R => '0',
   Q => ROTR11_out_5
);
e_reg_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => e_7_i_1_n_0,
   R => '0',
   Q => ROTR11_out_4
);
e_reg_7_i_2 : CARRY4
 port map (
   CI => e_reg_3_i_2_n_0,
   CYINIT => '0',
   DI(0) => d_4,
   DI(1) => d_5,
   DI(2) => d_6,
   DI(3) => d_7,
   S(0) => e_7_i_6_n_0,
   S(1) => e_7_i_5_n_0,
   S(2) => e_7_i_4_n_0,
   S(3) => e_7_i_3_n_0,
   CO(0) => e_reg_7_i_2_n_3,
   CO(1) => e_reg_7_i_2_n_2,
   CO(2) => e_reg_7_i_2_n_1,
   CO(3) => e_reg_7_i_2_n_0,
   O(0) => in15_4,
   O(1) => in15_5,
   O(2) => in15_6,
   O(3) => in15_7
);
e_reg_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => e_8_i_1_n_0,
   R => '0',
   Q => ROTR11_out_3
);
e_reg_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => e_9_i_1_n_0,
   R => '0',
   Q => ROTR11_out_2
);
finished_OBUF_inst : OBUF
 port map (
   I => finished_OBUF,
   O => finished
);
FSM_onehot_CURRENT_STATE_0_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_0,
   I1 => rst_IBUF,
   O => FSM_onehot_CURRENT_STATE_0_i_1_n_0
);
FSM_onehot_CURRENT_STATE_10_i_1 : LUT2
  generic map(
   INIT => X"e"
  )
 port map (
   I0 => finished_OBUF,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   O => FSM_onehot_CURRENT_STATE_10_i_1_n_0
);
FSM_onehot_CURRENT_STATE_11_i_1 : LUT4
  generic map(
   INIT => X"a8aa"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_8,
   I1 => FSM_onehot_CURRENT_STATE_11_i_2_n_0,
   I2 => FSM_onehot_CURRENT_STATE_11_i_3_n_0,
   I3 => FSM_onehot_CURRENT_STATE_11_i_4_n_0,
   O => FSM_onehot_CURRENT_STATE_11_i_1_n_0
);
FSM_onehot_CURRENT_STATE_11_i_2 : LUT5
  generic map(
   INIT => X"fffffffe"
  )
 port map (
   I0 => HASH_02_COUNTER_7,
   I1 => HASH_02_COUNTER_28,
   I2 => HASH_02_COUNTER_16,
   I3 => HASH_02_COUNTER_17,
   I4 => FSM_onehot_CURRENT_STATE_11_i_5_n_0,
   O => FSM_onehot_CURRENT_STATE_11_i_2_n_0
);
FSM_onehot_CURRENT_STATE_11_i_3 : LUT5
  generic map(
   INIT => X"fffffffe"
  )
 port map (
   I0 => HASH_02_COUNTER_3,
   I1 => HASH_02_COUNTER_29,
   I2 => HASH_02_COUNTER_5,
   I3 => HASH_02_COUNTER_18,
   I4 => FSM_onehot_CURRENT_STATE_11_i_6_n_0,
   O => FSM_onehot_CURRENT_STATE_11_i_3_n_0
);
FSM_onehot_CURRENT_STATE_11_i_4 : LUT6
  generic map(
   INIT => X"0000000000040000"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_11_i_7_n_0,
   I1 => FSM_onehot_CURRENT_STATE_11_i_8_n_0,
   I2 => FSM_onehot_CURRENT_STATE_11_i_9_n_0,
   I3 => HASH_02_COUNTER_0,
   I4 => HASH_02_COUNTER_6,
   I5 => HASH_02_COUNTER_12,
   O => FSM_onehot_CURRENT_STATE_11_i_4_n_0
);
FSM_onehot_CURRENT_STATE_11_i_5 : LUT4
  generic map(
   INIT => X"fffe"
  )
 port map (
   I0 => HASH_02_COUNTER_30,
   I1 => HASH_02_COUNTER_19,
   I2 => HASH_02_COUNTER_23,
   I3 => HASH_02_COUNTER_8,
   O => FSM_onehot_CURRENT_STATE_11_i_5_n_0
);
FSM_onehot_CURRENT_STATE_11_i_6 : LUT4
  generic map(
   INIT => X"fffe"
  )
 port map (
   I0 => HASH_02_COUNTER_20,
   I1 => HASH_02_COUNTER_11,
   I2 => HASH_02_COUNTER_25,
   I3 => HASH_02_COUNTER_2,
   O => FSM_onehot_CURRENT_STATE_11_i_6_n_0
);
FSM_onehot_CURRENT_STATE_11_i_7 : LUT4
  generic map(
   INIT => X"fffe"
  )
 port map (
   I0 => HASH_02_COUNTER_27,
   I1 => HASH_02_COUNTER_26,
   I2 => HASH_02_COUNTER_24,
   I3 => HASH_02_COUNTER_15,
   O => FSM_onehot_CURRENT_STATE_11_i_7_n_0
);
FSM_onehot_CURRENT_STATE_11_i_8 : LUT4
  generic map(
   INIT => X"0001"
  )
 port map (
   I0 => HASH_02_COUNTER_22,
   I1 => HASH_02_COUNTER_13,
   I2 => HASH_02_COUNTER_14,
   I3 => HASH_02_COUNTER_1,
   O => FSM_onehot_CURRENT_STATE_11_i_8_n_0
);
FSM_onehot_CURRENT_STATE_11_i_9 : LUT4
  generic map(
   INIT => X"fffe"
  )
 port map (
   I0 => HASH_02_COUNTER_21,
   I1 => HASH_02_COUNTER_10,
   I2 => HASH_02_COUNTER_9,
   I3 => HASH_02_COUNTER_4,
   O => FSM_onehot_CURRENT_STATE_11_i_9_n_0
);
FSM_onehot_CURRENT_STATE_11_rep_i_1 : LUT4
  generic map(
   INIT => X"a8aa"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_8,
   I1 => FSM_onehot_CURRENT_STATE_11_i_2_n_0,
   I2 => FSM_onehot_CURRENT_STATE_11_i_3_n_0,
   I3 => FSM_onehot_CURRENT_STATE_11_i_4_n_0,
   O => FSM_onehot_CURRENT_STATE_11_rep_i_1_n_0
);
FSM_onehot_CURRENT_STATE_1_i_1 : LUT4
  generic map(
   INIT => X"4f44"
  )
 port map (
   I0 => data_ready_IBUF,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_1,
   I2 => rst_IBUF,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_0,
   O => FSM_onehot_CURRENT_STATE_1_i_1_n_0
);
FSM_onehot_CURRENT_STATE_2_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => data_ready_IBUF,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_1,
   O => FSM_onehot_CURRENT_STATE_2_i_1_n_0
);
FSM_onehot_CURRENT_STATE_8_i_1 : LUT2
  generic map(
   INIT => X"e"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_12,
   O => FSM_onehot_CURRENT_STATE_8_i_1_n_0
);
FSM_onehot_CURRENT_STATE_9_i_1 : LUT4
  generic map(
   INIT => X"0200"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_8,
   I1 => FSM_onehot_CURRENT_STATE_11_i_2_n_0,
   I2 => FSM_onehot_CURRENT_STATE_11_i_3_n_0,
   I3 => FSM_onehot_CURRENT_STATE_11_i_4_n_0,
   O => FSM_onehot_CURRENT_STATE_9_i_1_n_0
);
FSM_onehot_CURRENT_STATE_reg_0 : FDPE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => '1',
   D => FSM_onehot_CURRENT_STATE_0_i_1_n_0,
   PRE => rst_IBUF,
   Q => FSM_onehot_CURRENT_STATE_reg_n_0_0
);
FSM_onehot_CURRENT_STATE_reg_10 : FDCE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => '1',
   CLR => rst_IBUF,
   D => FSM_onehot_CURRENT_STATE_10_i_1_n_0,
   Q => finished_OBUF
);
FSM_onehot_CURRENT_STATE_reg_11 : FDCE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => '1',
   CLR => rst_IBUF,
   D => FSM_onehot_CURRENT_STATE_11_i_1_n_0,
   Q => FSM_onehot_CURRENT_STATE_reg_n_0_11
);
FSM_onehot_CURRENT_STATE_reg_11_rep : FDCE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => '1',
   CLR => rst_IBUF,
   D => FSM_onehot_CURRENT_STATE_11_rep_i_1_n_0,
   Q => FSM_onehot_CURRENT_STATE_reg_11_rep_n_0
);
FSM_onehot_CURRENT_STATE_reg_12 : FDCE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => '1',
   CLR => rst_IBUF,
   D => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   Q => FSM_onehot_CURRENT_STATE_reg_n_0_12
);
FSM_onehot_CURRENT_STATE_reg_1 : FDCE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => '1',
   CLR => rst_IBUF,
   D => FSM_onehot_CURRENT_STATE_1_i_1_n_0,
   Q => FSM_onehot_CURRENT_STATE_reg_n_0_1
);
FSM_onehot_CURRENT_STATE_reg_2 : FDCE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => '1',
   CLR => rst_IBUF,
   D => FSM_onehot_CURRENT_STATE_2_i_1_n_0,
   Q => M_0
);
FSM_onehot_CURRENT_STATE_reg_3 : FDCE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => '1',
   CLR => rst_IBUF,
   D => M_0,
   Q => W_0
);
FSM_onehot_CURRENT_STATE_reg_4 : FDCE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => '1',
   CLR => rst_IBUF,
   D => W_0,
   Q => W_16
);
FSM_onehot_CURRENT_STATE_reg_5 : FDCE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => '1',
   CLR => rst_IBUF,
   D => W_16,
   Q => W_32
);
FSM_onehot_CURRENT_STATE_reg_6 : FDCE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => '1',
   CLR => rst_IBUF,
   D => W_32,
   Q => W_48
);
FSM_onehot_CURRENT_STATE_reg_7 : FDCE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => '1',
   CLR => rst_IBUF,
   D => W_48,
   Q => FSM_onehot_CURRENT_STATE_reg_n_0_7
);
FSM_onehot_CURRENT_STATE_reg_7_rep : FDCE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => '1',
   CLR => rst_IBUF,
   D => W_48,
   Q => FSM_onehot_CURRENT_STATE_reg_7_rep_n_0
);
FSM_onehot_CURRENT_STATE_reg_8 : FDCE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => '1',
   CLR => rst_IBUF,
   D => FSM_onehot_CURRENT_STATE_8_i_1_n_0,
   Q => FSM_onehot_CURRENT_STATE_reg_n_0_8
);
FSM_onehot_CURRENT_STATE_reg_9 : FDCE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => '1',
   CLR => rst_IBUF,
   D => FSM_onehot_CURRENT_STATE_9_i_1_n_0,
   Q => FSM_onehot_CURRENT_STATE_reg_n_0_9
);
f_0_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => ROTR11_out_11,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_64,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => f_0_i_1_n_0
);
f_10_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => ROTR11_out_1,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_74,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => f_10_i_1_n_0
);
f_11_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => ROTR11_out_32,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_75,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => f_11_i_1_n_0
);
f_12_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => ROTR11_out_31,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_76,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => f_12_i_1_n_0
);
f_13_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => ROTR11_out_30,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_77,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => f_13_i_1_n_0
);
f_14_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => ROTR11_out_29,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_78,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => f_14_i_1_n_0
);
f_15_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => ROTR11_out_28,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_79,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => f_15_i_1_n_0
);
f_16_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => ROTR11_out_27,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_80,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => f_16_i_1_n_0
);
f_17_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => ROTR11_out_26,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_81,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => f_17_i_1_n_0
);
f_18_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => ROTR11_out_25,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_82,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => f_18_i_1_n_0
);
f_19_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => ROTR11_out_24,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_83,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => f_19_i_1_n_0
);
f_1_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => ROTR11_out_10,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_65,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => f_1_i_1_n_0
);
f_20_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => ROTR11_out_23,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_84,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => f_20_i_1_n_0
);
f_21_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => ROTR11_out_22,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_85,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => f_21_i_1_n_0
);
f_22_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => ROTR11_out_21,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_86,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => f_22_i_1_n_0
);
f_23_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => ROTR11_out_20,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_87,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => f_23_i_1_n_0
);
f_24_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => ROTR11_out_19,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_88,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => f_24_i_1_n_0
);
f_25_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => ROTR11_out_18,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_89,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => f_25_i_1_n_0
);
f_26_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => ROTR11_out_17,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_90,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => f_26_i_1_n_0
);
f_27_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => ROTR11_out_16,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_91,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => f_27_i_1_n_0
);
f_28_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => ROTR11_out_15,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_92,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => f_28_i_1_n_0
);
f_29_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => ROTR11_out_14,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_93,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => f_29_i_1_n_0
);
f_2_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => ROTR11_out_9,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_66,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => f_2_i_1_n_0
);
f_30_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => ROTR11_out_13,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_94,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => f_30_i_1_n_0
);
f_31_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => ROTR11_out_12,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_95,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => f_31_i_1_n_0
);
f_3_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => ROTR11_out_8,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_67,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => f_3_i_1_n_0
);
f_4_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => ROTR11_out_7,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_68,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => f_4_i_1_n_0
);
f_5_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => ROTR11_out_6,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_69,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => f_5_i_1_n_0
);
f_6_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => ROTR11_out_5,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_70,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => f_6_i_1_n_0
);
f_7_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => ROTR11_out_4,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_71,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => f_7_i_1_n_0
);
f_8_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => ROTR11_out_3,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_72,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => f_8_i_1_n_0
);
f_9_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => ROTR11_out_2,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_73,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => f_9_i_1_n_0
);
f_reg_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => f_0_i_1_n_0,
   R => '0',
   Q => f_reg_n_0_0
);
f_reg_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => f_10_i_1_n_0,
   R => '0',
   Q => f_reg_n_0_10
);
f_reg_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => f_11_i_1_n_0,
   R => '0',
   Q => f_reg_n_0_11
);
f_reg_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => f_12_i_1_n_0,
   R => '0',
   Q => f_reg_n_0_12
);
f_reg_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => f_13_i_1_n_0,
   R => '0',
   Q => f_reg_n_0_13
);
f_reg_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => f_14_i_1_n_0,
   R => '0',
   Q => f_reg_n_0_14
);
f_reg_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => f_15_i_1_n_0,
   R => '0',
   Q => f_reg_n_0_15
);
f_reg_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => f_16_i_1_n_0,
   R => '0',
   Q => f_reg_n_0_16
);
f_reg_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => f_17_i_1_n_0,
   R => '0',
   Q => f_reg_n_0_17
);
f_reg_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => f_18_i_1_n_0,
   R => '0',
   Q => f_reg_n_0_18
);
f_reg_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => f_19_i_1_n_0,
   R => '0',
   Q => f_reg_n_0_19
);
f_reg_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => f_1_i_1_n_0,
   R => '0',
   Q => f_reg_n_0_1
);
f_reg_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => f_20_i_1_n_0,
   R => '0',
   Q => f_reg_n_0_20
);
f_reg_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => f_21_i_1_n_0,
   R => '0',
   Q => f_reg_n_0_21
);
f_reg_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => f_22_i_1_n_0,
   R => '0',
   Q => f_reg_n_0_22
);
f_reg_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => f_23_i_1_n_0,
   R => '0',
   Q => f_reg_n_0_23
);
f_reg_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => f_24_i_1_n_0,
   R => '0',
   Q => f_reg_n_0_24
);
f_reg_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => f_25_i_1_n_0,
   R => '0',
   Q => f_reg_n_0_25
);
f_reg_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => f_26_i_1_n_0,
   R => '0',
   Q => f_reg_n_0_26
);
f_reg_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => f_27_i_1_n_0,
   R => '0',
   Q => f_reg_n_0_27
);
f_reg_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => f_28_i_1_n_0,
   R => '0',
   Q => f_reg_n_0_28
);
f_reg_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => f_29_i_1_n_0,
   R => '0',
   Q => f_reg_n_0_29
);
f_reg_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => f_2_i_1_n_0,
   R => '0',
   Q => f_reg_n_0_2
);
f_reg_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => f_30_i_1_n_0,
   R => '0',
   Q => f_reg_n_0_30
);
f_reg_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => f_31_i_1_n_0,
   R => '0',
   Q => f_reg_n_0_31
);
f_reg_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => f_3_i_1_n_0,
   R => '0',
   Q => f_reg_n_0_3
);
f_reg_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => f_4_i_1_n_0,
   R => '0',
   Q => f_reg_n_0_4
);
f_reg_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => f_5_i_1_n_0,
   R => '0',
   Q => f_reg_n_0_5
);
f_reg_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => f_6_i_1_n_0,
   R => '0',
   Q => f_reg_n_0_6
);
f_reg_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => f_7_i_1_n_0,
   R => '0',
   Q => f_reg_n_0_7
);
f_reg_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => f_8_i_1_n_0,
   R => '0',
   Q => f_reg_n_0_8
);
f_reg_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => f_9_i_1_n_0,
   R => '0',
   Q => f_reg_n_0_9
);
g0_b0 : LUT6
  generic map(
   INIT => X"62d85ba9fa114abe"
  )
 port map (
   I0 => HASH_02_COUNTER_0,
   I1 => HASH_02_COUNTER_1,
   I2 => HASH_02_COUNTER_2,
   I3 => HASH_02_COUNTER_3,
   I4 => HASH_02_COUNTER_4,
   I5 => HASH_02_COUNTER_5,
   O => g0_b0_n_0
);
g0_b1 : LUT6
  generic map(
   INIT => X"f3f10a68b9b66c14"
  )
 port map (
   I0 => HASH_02_COUNTER_0,
   I1 => HASH_02_COUNTER_1,
   I2 => HASH_02_COUNTER_2,
   I3 => HASH_02_COUNTER_3,
   I4 => HASH_02_COUNTER_4,
   I5 => HASH_02_COUNTER_5,
   O => g0_b1_n_0
);
g0_b10 : LUT6
  generic map(
   INIT => X"309e628c0e365c83"
  )
 port map (
   I0 => HASH_02_COUNTER_0,
   I1 => HASH_02_COUNTER_1,
   I2 => HASH_02_COUNTER_2,
   I3 => HASH_02_COUNTER_3,
   I4 => HASH_02_COUNTER_4,
   I5 => HASH_02_COUNTER_5,
   O => g0_b10_n_0
);
g0_b11 : LUT6
  generic map(
   INIT => X"b4fa15ed98d51b8d"
  )
 port map (
   I0 => HASH_02_COUNTER_0,
   I1 => HASH_02_COUNTER_1,
   I2 => HASH_02_COUNTER_2,
   I3 => HASH_02_COUNTER_3,
   I4 => HASH_02_COUNTER_4,
   I5 => HASH_02_COUNTER_5,
   O => g0_b11_n_0
);
g0_b12 : LUT6
  generic map(
   INIT => X"940c48102904baac"
  )
 port map (
   I0 => HASH_02_COUNTER_0,
   I1 => HASH_02_COUNTER_1,
   I2 => HASH_02_COUNTER_2,
   I3 => HASH_02_COUNTER_3,
   I4 => HASH_02_COUNTER_4,
   I5 => HASH_02_COUNTER_5,
   O => g0_b12_n_0
);
g0_b13 : LUT6
  generic map(
   INIT => X"f6aed396cc59a905"
  )
 port map (
   I0 => HASH_02_COUNTER_0,
   I1 => HASH_02_COUNTER_1,
   I2 => HASH_02_COUNTER_2,
   I3 => HASH_02_COUNTER_3,
   I4 => HASH_02_COUNTER_4,
   I5 => HASH_02_COUNTER_5,
   O => g0_b13_n_0
);
g0_b14 : LUT6
  generic map(
   INIT => X"b6c71b544b039a9e"
  )
 port map (
   I0 => HASH_02_COUNTER_0,
   I1 => HASH_02_COUNTER_1,
   I2 => HASH_02_COUNTER_2,
   I3 => HASH_02_COUNTER_3,
   I4 => HASH_02_COUNTER_4,
   I5 => HASH_02_COUNTER_5,
   O => g0_b14_n_0
);
g0_b15 : LUT6
  generic map(
   INIT => X"5169954022eca55c"
  )
 port map (
   I0 => HASH_02_COUNTER_0,
   I1 => HASH_02_COUNTER_1,
   I2 => HASH_02_COUNTER_2,
   I3 => HASH_02_COUNTER_3,
   I4 => HASH_02_COUNTER_4,
   I5 => HASH_02_COUNTER_5,
   O => g0_b15_n_0
);
g0_b16 : LUT6
  generic map(
   INIT => X"cb022503ae95876a"
  )
 port map (
   I0 => HASH_02_COUNTER_0,
   I1 => HASH_02_COUNTER_1,
   I2 => HASH_02_COUNTER_2,
   I3 => HASH_02_COUNTER_3,
   I4 => HASH_02_COUNTER_4,
   I5 => HASH_02_COUNTER_5,
   O => g0_b16_n_0
);
g0_b17 : LUT6
  generic map(
   INIT => X"1982d7f36503b353"
  )
 port map (
   I0 => HASH_02_COUNTER_0,
   I1 => HASH_02_COUNTER_1,
   I2 => HASH_02_COUNTER_2,
   I3 => HASH_02_COUNTER_3,
   I4 => HASH_02_COUNTER_4,
   I5 => HASH_02_COUNTER_5,
   O => g0_b17_n_0
);
g0_b18 : LUT6
  generic map(
   INIT => X"1bd34905212a79da"
  )
 port map (
   I0 => HASH_02_COUNTER_0,
   I1 => HASH_02_COUNTER_1,
   I2 => HASH_02_COUNTER_2,
   I3 => HASH_02_COUNTER_3,
   I4 => HASH_02_COUNTER_4,
   I5 => HASH_02_COUNTER_5,
   O => g0_b18_n_0
);
g0_b19 : LUT6
  generic map(
   INIT => X"55f4ef3ec99bf8c1"
  )
 port map (
   I0 => HASH_02_COUNTER_0,
   I1 => HASH_02_COUNTER_1,
   I2 => HASH_02_COUNTER_2,
   I3 => HASH_02_COUNTER_3,
   I4 => HASH_02_COUNTER_4,
   I5 => HASH_02_COUNTER_5,
   O => g0_b19_n_0
);
g0_b2 : LUT6
  generic map(
   INIT => X"474d60d5aa5ef4cc"
  )
 port map (
   I0 => HASH_02_COUNTER_0,
   I1 => HASH_02_COUNTER_1,
   I2 => HASH_02_COUNTER_2,
   I3 => HASH_02_COUNTER_3,
   I4 => HASH_02_COUNTER_4,
   I5 => HASH_02_COUNTER_5,
   O => g0_b2_n_0
);
g0_b20 : LUT6
  generic map(
   INIT => X"f07a338b0be3f4fa"
  )
 port map (
   I0 => HASH_02_COUNTER_0,
   I1 => HASH_02_COUNTER_1,
   I2 => HASH_02_COUNTER_2,
   I3 => HASH_02_COUNTER_3,
   I4 => HASH_02_COUNTER_4,
   I5 => HASH_02_COUNTER_5,
   O => g0_b20_n_0
);
g0_b21 : LUT6
  generic map(
   INIT => X"d28b89adb3f2146a"
  )
 port map (
   I0 => HASH_02_COUNTER_0,
   I1 => HASH_02_COUNTER_1,
   I2 => HASH_02_COUNTER_2,
   I3 => HASH_02_COUNTER_3,
   I4 => HASH_02_COUNTER_4,
   I5 => HASH_02_COUNTER_5,
   O => g0_b21_n_0
);
g0_b22 : LUT6
  generic map(
   INIT => X"ec248ce058b46034"
  )
 port map (
   I0 => HASH_02_COUNTER_0,
   I1 => HASH_02_COUNTER_1,
   I2 => HASH_02_COUNTER_2,
   I3 => HASH_02_COUNTER_3,
   I4 => HASH_02_COUNTER_4,
   I5 => HASH_02_COUNTER_5,
   O => g0_b22_n_0
);
g0_b23 : LUT6
  generic map(
   INIT => X"5f69314170d7f22d"
  )
 port map (
   I0 => HASH_02_COUNTER_0,
   I1 => HASH_02_COUNTER_1,
   I2 => HASH_02_COUNTER_2,
   I3 => HASH_02_COUNTER_3,
   I4 => HASH_02_COUNTER_4,
   I5 => HASH_02_COUNTER_5,
   O => g0_b23_n_0
);
g0_b24 : LUT6
  generic map(
   INIT => X"0055185d2816c8be"
  )
 port map (
   I0 => HASH_02_COUNTER_0,
   I1 => HASH_02_COUNTER_1,
   I2 => HASH_02_COUNTER_2,
   I3 => HASH_02_COUNTER_3,
   I4 => HASH_02_COUNTER_4,
   I5 => HASH_02_COUNTER_5,
   O => g0_b24_n_0
);
g0_b25 : LUT6
  generic map(
   INIT => X"c0662dab58a652c1"
  )
 port map (
   I0 => HASH_02_COUNTER_0,
   I1 => HASH_02_COUNTER_1,
   I2 => HASH_02_COUNTER_2,
   I3 => HASH_02_COUNTER_3,
   I4 => HASH_02_COUNTER_4,
   I5 => HASH_02_COUNTER_5,
   O => g0_b25_n_0
);
g0_b26 : LUT6
  generic map(
   INIT => X"ed2e6837f8df0c04"
  )
 port map (
   I0 => HASH_02_COUNTER_0,
   I1 => HASH_02_COUNTER_1,
   I2 => HASH_02_COUNTER_2,
   I3 => HASH_02_COUNTER_3,
   I4 => HASH_02_COUNTER_4,
   I5 => HASH_02_COUNTER_5,
   O => g0_b26_n_0
);
g0_b27 : LUT6
  generic map(
   INIT => X"4af302060b7641b8"
  )
 port map (
   I0 => HASH_02_COUNTER_0,
   I1 => HASH_02_COUNTER_1,
   I2 => HASH_02_COUNTER_2,
   I3 => HASH_02_COUNTER_3,
   I4 => HASH_02_COUNTER_4,
   I5 => HASH_02_COUNTER_5,
   O => g0_b27_n_0
);
g0_b28 : LUT6
  generic map(
   INIT => X"535bf0a8adc05b76"
  )
 port map (
   I0 => HASH_02_COUNTER_0,
   I1 => HASH_02_COUNTER_1,
   I2 => HASH_02_COUNTER_2,
   I3 => HASH_02_COUNTER_3,
   I4 => HASH_02_COUNTER_4,
   I5 => HASH_02_COUNTER_5,
   O => g0_b28_n_0
);
g0_b29 : LUT6
  generic map(
   INIT => X"639c43330e9b149e"
  )
 port map (
   I0 => HASH_02_COUNTER_0,
   I1 => HASH_02_COUNTER_1,
   I2 => HASH_02_COUNTER_2,
   I3 => HASH_02_COUNTER_3,
   I4 => HASH_02_COUNTER_4,
   I5 => HASH_02_COUNTER_5,
   O => g0_b29_n_0
);
g0_b3 : LUT6
  generic map(
   INIT => X"3b66126606f82515"
  )
 port map (
   I0 => HASH_02_COUNTER_0,
   I1 => HASH_02_COUNTER_1,
   I2 => HASH_02_COUNTER_2,
   I3 => HASH_02_COUNTER_3,
   I4 => HASH_02_COUNTER_4,
   I5 => HASH_02_COUNTER_5,
   O => g0_b3_n_0
);
g0_b30 : LUT6
  generic map(
   INIT => X"83e07c3c30e3992b"
  )
 port map (
   I0 => HASH_02_COUNTER_0,
   I1 => HASH_02_COUNTER_1,
   I2 => HASH_02_COUNTER_2,
   I3 => HASH_02_COUNTER_3,
   I4 => HASH_02_COUNTER_4,
   I5 => HASH_02_COUNTER_5,
   O => g0_b30_n_0
);
g0_b31 : LUT6
  generic map(
   INIT => X"fc007fc03f03e1cc"
  )
 port map (
   I0 => HASH_02_COUNTER_0,
   I1 => HASH_02_COUNTER_1,
   I2 => HASH_02_COUNTER_2,
   I3 => HASH_02_COUNTER_3,
   I4 => HASH_02_COUNTER_4,
   I5 => HASH_02_COUNTER_5,
   O => g0_b31_n_0
);
g0_b4 : LUT6
  generic map(
   INIT => X"d499943e51c0b5b3"
  )
 port map (
   I0 => HASH_02_COUNTER_0,
   I1 => HASH_02_COUNTER_1,
   I2 => HASH_02_COUNTER_2,
   I3 => HASH_02_COUNTER_3,
   I4 => HASH_02_COUNTER_4,
   I5 => HASH_02_COUNTER_5,
   O => g0_b4_n_0
);
g0_b5 : LUT6
  generic map(
   INIT => X"f398ad669230f468"
  )
 port map (
   I0 => HASH_02_COUNTER_0,
   I1 => HASH_02_COUNTER_1,
   I2 => HASH_02_COUNTER_2,
   I3 => HASH_02_COUNTER_3,
   I4 => HASH_02_COUNTER_4,
   I5 => HASH_02_COUNTER_5,
   O => g0_b5_n_0
);
g0_b6 : LUT6
  generic map(
   INIT => X"f3e48614ffddb8b4"
  )
 port map (
   I0 => HASH_02_COUNTER_0,
   I1 => HASH_02_COUNTER_1,
   I2 => HASH_02_COUNTER_2,
   I3 => HASH_02_COUNTER_3,
   I4 => HASH_02_COUNTER_4,
   I5 => HASH_02_COUNTER_5,
   O => g0_b6_n_0
);
g0_b7 : LUT6
  generic map(
   INIT => X"f19849a51cef6def"
  )
 port map (
   I0 => HASH_02_COUNTER_0,
   I1 => HASH_02_COUNTER_1,
   I2 => HASH_02_COUNTER_2,
   I3 => HASH_02_COUNTER_3,
   I4 => HASH_02_COUNTER_4,
   I5 => HASH_02_COUNTER_5,
   O => g0_b7_n_0
);
g0_b8 : LUT6
  generic map(
   INIT => X"52854c5efd4fbe2d"
  )
 port map (
   I0 => HASH_02_COUNTER_0,
   I1 => HASH_02_COUNTER_1,
   I2 => HASH_02_COUNTER_2,
   I3 => HASH_02_COUNTER_3,
   I4 => HASH_02_COUNTER_4,
   I5 => HASH_02_COUNTER_5,
   O => g0_b8_n_0
);
g0_b9 : LUT6
  generic map(
   INIT => X"5be426315e0243dd"
  )
 port map (
   I0 => HASH_02_COUNTER_0,
   I1 => HASH_02_COUNTER_1,
   I2 => HASH_02_COUNTER_2,
   I3 => HASH_02_COUNTER_3,
   I4 => HASH_02_COUNTER_4,
   I5 => HASH_02_COUNTER_5,
   O => g0_b9_n_0
);
g_0_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => f_reg_n_0_0,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_32,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => g_0_i_1_n_0
);
g_10_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => f_reg_n_0_10,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_42,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => g_10_i_1_n_0
);
g_11_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => f_reg_n_0_11,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_43,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => g_11_i_1_n_0
);
g_12_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => f_reg_n_0_12,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_44,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => g_12_i_1_n_0
);
g_13_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => f_reg_n_0_13,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_45,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => g_13_i_1_n_0
);
g_14_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => f_reg_n_0_14,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_46,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => g_14_i_1_n_0
);
g_15_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => f_reg_n_0_15,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_47,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => g_15_i_1_n_0
);
g_16_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => f_reg_n_0_16,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_48,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => g_16_i_1_n_0
);
g_17_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => f_reg_n_0_17,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_49,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => g_17_i_1_n_0
);
g_18_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => f_reg_n_0_18,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_50,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => g_18_i_1_n_0
);
g_19_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => f_reg_n_0_19,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_51,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => g_19_i_1_n_0
);
g_1_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => f_reg_n_0_1,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_33,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => g_1_i_1_n_0
);
g_20_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => f_reg_n_0_20,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_52,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => g_20_i_1_n_0
);
g_21_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => f_reg_n_0_21,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_53,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => g_21_i_1_n_0
);
g_22_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => f_reg_n_0_22,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_54,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => g_22_i_1_n_0
);
g_23_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => f_reg_n_0_23,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_55,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => g_23_i_1_n_0
);
g_24_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => f_reg_n_0_24,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_56,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => g_24_i_1_n_0
);
g_25_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => f_reg_n_0_25,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_57,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => g_25_i_1_n_0
);
g_26_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => f_reg_n_0_26,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_58,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => g_26_i_1_n_0
);
g_27_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => f_reg_n_0_27,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_59,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => g_27_i_1_n_0
);
g_28_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => f_reg_n_0_28,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_60,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => g_28_i_1_n_0
);
g_29_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => f_reg_n_0_29,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_61,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => g_29_i_1_n_0
);
g_2_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => f_reg_n_0_2,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_34,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => g_2_i_1_n_0
);
g_30_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => f_reg_n_0_30,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_62,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => g_30_i_1_n_0
);
g_31_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => f_reg_n_0_31,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_63,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => g_31_i_1_n_0
);
g_3_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => f_reg_n_0_3,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_35,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => g_3_i_1_n_0
);
g_4_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => f_reg_n_0_4,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_36,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => g_4_i_1_n_0
);
g_5_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => f_reg_n_0_5,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_37,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => g_5_i_1_n_0
);
g_6_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => f_reg_n_0_6,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_38,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => g_6_i_1_n_0
);
g_7_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => f_reg_n_0_7,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_39,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => g_7_i_1_n_0
);
g_8_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => f_reg_n_0_8,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_40,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => g_8_i_1_n_0
);
g_9_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => f_reg_n_0_9,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_41,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => g_9_i_1_n_0
);
g_reg_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => g_0_i_1_n_0,
   R => '0',
   Q => g_reg_n_0_0
);
g_reg_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => g_10_i_1_n_0,
   R => '0',
   Q => g_reg_n_0_10
);
g_reg_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => g_11_i_1_n_0,
   R => '0',
   Q => g_reg_n_0_11
);
g_reg_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => g_12_i_1_n_0,
   R => '0',
   Q => g_reg_n_0_12
);
g_reg_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => g_13_i_1_n_0,
   R => '0',
   Q => g_reg_n_0_13
);
g_reg_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => g_14_i_1_n_0,
   R => '0',
   Q => g_reg_n_0_14
);
g_reg_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => g_15_i_1_n_0,
   R => '0',
   Q => g_reg_n_0_15
);
g_reg_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => g_16_i_1_n_0,
   R => '0',
   Q => g_reg_n_0_16
);
g_reg_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => g_17_i_1_n_0,
   R => '0',
   Q => g_reg_n_0_17
);
g_reg_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => g_18_i_1_n_0,
   R => '0',
   Q => g_reg_n_0_18
);
g_reg_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => g_19_i_1_n_0,
   R => '0',
   Q => g_reg_n_0_19
);
g_reg_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => g_1_i_1_n_0,
   R => '0',
   Q => g_reg_n_0_1
);
g_reg_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => g_20_i_1_n_0,
   R => '0',
   Q => g_reg_n_0_20
);
g_reg_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => g_21_i_1_n_0,
   R => '0',
   Q => g_reg_n_0_21
);
g_reg_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => g_22_i_1_n_0,
   R => '0',
   Q => g_reg_n_0_22
);
g_reg_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => g_23_i_1_n_0,
   R => '0',
   Q => g_reg_n_0_23
);
g_reg_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => g_24_i_1_n_0,
   R => '0',
   Q => g_reg_n_0_24
);
g_reg_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => g_25_i_1_n_0,
   R => '0',
   Q => g_reg_n_0_25
);
g_reg_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => g_26_i_1_n_0,
   R => '0',
   Q => g_reg_n_0_26
);
g_reg_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => g_27_i_1_n_0,
   R => '0',
   Q => g_reg_n_0_27
);
g_reg_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => g_28_i_1_n_0,
   R => '0',
   Q => g_reg_n_0_28
);
g_reg_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => g_29_i_1_n_0,
   R => '0',
   Q => g_reg_n_0_29
);
g_reg_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => g_2_i_1_n_0,
   R => '0',
   Q => g_reg_n_0_2
);
g_reg_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => g_30_i_1_n_0,
   R => '0',
   Q => g_reg_n_0_30
);
g_reg_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => g_31_i_1_n_0,
   R => '0',
   Q => g_reg_n_0_31
);
g_reg_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => g_3_i_1_n_0,
   R => '0',
   Q => g_reg_n_0_3
);
g_reg_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => g_4_i_1_n_0,
   R => '0',
   Q => g_reg_n_0_4
);
g_reg_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => g_5_i_1_n_0,
   R => '0',
   Q => g_reg_n_0_5
);
g_reg_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => g_6_i_1_n_0,
   R => '0',
   Q => g_reg_n_0_6
);
g_reg_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => g_7_i_1_n_0,
   R => '0',
   Q => g_reg_n_0_7
);
g_reg_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => g_8_i_1_n_0,
   R => '0',
   Q => g_reg_n_0_8
);
g_reg_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => g_9_i_1_n_0,
   R => '0',
   Q => g_reg_n_0_9
);
HASH_02_COUNTER_0_i_1 : LUT1
  generic map(
   INIT => X"1"
  )
 port map (
   I0 => HASH_02_COUNTER_0,
   O => HASH_02_COUNTER_0_i_1_n_0
);
HASH_02_COUNTER_30_i_1 : LUT4
  generic map(
   INIT => X"000e"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_0,
   I1 => FSM_onehot_CURRENT_STATE_9_i_1_n_0,
   I2 => rst_IBUF,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_12,
   O => HASH_02_COUNTER_30_i_1_n_0
);
HASH_02_COUNTER_30_i_2 : LUT4
  generic map(
   INIT => X"5554"
  )
 port map (
   I0 => rst_IBUF,
   I1 => FSM_onehot_CURRENT_STATE_9_i_1_n_0,
   I2 => FSM_onehot_CURRENT_STATE_reg_n_0_0,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_12,
   O => HASH_02_COUNTER_30_i_2_n_0
);
HASH_02_COUNTER_reg_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HASH_02_COUNTER_30_i_2_n_0,
   D => HASH_02_COUNTER_0_i_1_n_0,
   R => HASH_02_COUNTER_30_i_1_n_0,
   Q => HASH_02_COUNTER_0
);
HASH_02_COUNTER_reg_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HASH_02_COUNTER_30_i_2_n_0,
   D => in32_10,
   R => HASH_02_COUNTER_30_i_1_n_0,
   Q => HASH_02_COUNTER_10
);
HASH_02_COUNTER_reg_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HASH_02_COUNTER_30_i_2_n_0,
   D => in32_11,
   R => HASH_02_COUNTER_30_i_1_n_0,
   Q => HASH_02_COUNTER_11
);
HASH_02_COUNTER_reg_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HASH_02_COUNTER_30_i_2_n_0,
   D => in32_12,
   R => HASH_02_COUNTER_30_i_1_n_0,
   Q => HASH_02_COUNTER_12
);
HASH_02_COUNTER_reg_12_i_1 : CARRY4
 port map (
   CI => HASH_02_COUNTER_reg_8_i_1_n_0,
   CYINIT => '0',
   DI(0) => '0',
   DI(1) => '0',
   DI(2) => '0',
   DI(3) => '0',
   S(0) => HASH_02_COUNTER_9,
   S(1) => HASH_02_COUNTER_10,
   S(2) => HASH_02_COUNTER_11,
   S(3) => HASH_02_COUNTER_12,
   CO(0) => HASH_02_COUNTER_reg_12_i_1_n_3,
   CO(1) => HASH_02_COUNTER_reg_12_i_1_n_2,
   CO(2) => HASH_02_COUNTER_reg_12_i_1_n_1,
   CO(3) => HASH_02_COUNTER_reg_12_i_1_n_0,
   O(0) => in32_9,
   O(1) => in32_10,
   O(2) => in32_11,
   O(3) => in32_12
);
HASH_02_COUNTER_reg_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HASH_02_COUNTER_30_i_2_n_0,
   D => in32_13,
   R => HASH_02_COUNTER_30_i_1_n_0,
   Q => HASH_02_COUNTER_13
);
HASH_02_COUNTER_reg_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HASH_02_COUNTER_30_i_2_n_0,
   D => in32_14,
   R => HASH_02_COUNTER_30_i_1_n_0,
   Q => HASH_02_COUNTER_14
);
HASH_02_COUNTER_reg_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HASH_02_COUNTER_30_i_2_n_0,
   D => in32_15,
   R => HASH_02_COUNTER_30_i_1_n_0,
   Q => HASH_02_COUNTER_15
);
HASH_02_COUNTER_reg_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HASH_02_COUNTER_30_i_2_n_0,
   D => in32_16,
   R => HASH_02_COUNTER_30_i_1_n_0,
   Q => HASH_02_COUNTER_16
);
HASH_02_COUNTER_reg_16_i_1 : CARRY4
 port map (
   CI => HASH_02_COUNTER_reg_12_i_1_n_0,
   CYINIT => '0',
   DI(0) => '0',
   DI(1) => '0',
   DI(2) => '0',
   DI(3) => '0',
   S(0) => HASH_02_COUNTER_13,
   S(1) => HASH_02_COUNTER_14,
   S(2) => HASH_02_COUNTER_15,
   S(3) => HASH_02_COUNTER_16,
   CO(0) => HASH_02_COUNTER_reg_16_i_1_n_3,
   CO(1) => HASH_02_COUNTER_reg_16_i_1_n_2,
   CO(2) => HASH_02_COUNTER_reg_16_i_1_n_1,
   CO(3) => HASH_02_COUNTER_reg_16_i_1_n_0,
   O(0) => in32_13,
   O(1) => in32_14,
   O(2) => in32_15,
   O(3) => in32_16
);
HASH_02_COUNTER_reg_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HASH_02_COUNTER_30_i_2_n_0,
   D => in32_17,
   R => HASH_02_COUNTER_30_i_1_n_0,
   Q => HASH_02_COUNTER_17
);
HASH_02_COUNTER_reg_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HASH_02_COUNTER_30_i_2_n_0,
   D => in32_18,
   R => HASH_02_COUNTER_30_i_1_n_0,
   Q => HASH_02_COUNTER_18
);
HASH_02_COUNTER_reg_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HASH_02_COUNTER_30_i_2_n_0,
   D => in32_19,
   R => HASH_02_COUNTER_30_i_1_n_0,
   Q => HASH_02_COUNTER_19
);
HASH_02_COUNTER_reg_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HASH_02_COUNTER_30_i_2_n_0,
   D => in32_1,
   R => HASH_02_COUNTER_30_i_1_n_0,
   Q => HASH_02_COUNTER_1
);
HASH_02_COUNTER_reg_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HASH_02_COUNTER_30_i_2_n_0,
   D => in32_20,
   R => HASH_02_COUNTER_30_i_1_n_0,
   Q => HASH_02_COUNTER_20
);
HASH_02_COUNTER_reg_20_i_1 : CARRY4
 port map (
   CI => HASH_02_COUNTER_reg_16_i_1_n_0,
   CYINIT => '0',
   DI(0) => '0',
   DI(1) => '0',
   DI(2) => '0',
   DI(3) => '0',
   S(0) => HASH_02_COUNTER_17,
   S(1) => HASH_02_COUNTER_18,
   S(2) => HASH_02_COUNTER_19,
   S(3) => HASH_02_COUNTER_20,
   CO(0) => HASH_02_COUNTER_reg_20_i_1_n_3,
   CO(1) => HASH_02_COUNTER_reg_20_i_1_n_2,
   CO(2) => HASH_02_COUNTER_reg_20_i_1_n_1,
   CO(3) => HASH_02_COUNTER_reg_20_i_1_n_0,
   O(0) => in32_17,
   O(1) => in32_18,
   O(2) => in32_19,
   O(3) => in32_20
);
HASH_02_COUNTER_reg_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HASH_02_COUNTER_30_i_2_n_0,
   D => in32_21,
   R => HASH_02_COUNTER_30_i_1_n_0,
   Q => HASH_02_COUNTER_21
);
HASH_02_COUNTER_reg_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HASH_02_COUNTER_30_i_2_n_0,
   D => in32_22,
   R => HASH_02_COUNTER_30_i_1_n_0,
   Q => HASH_02_COUNTER_22
);
HASH_02_COUNTER_reg_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HASH_02_COUNTER_30_i_2_n_0,
   D => in32_23,
   R => HASH_02_COUNTER_30_i_1_n_0,
   Q => HASH_02_COUNTER_23
);
HASH_02_COUNTER_reg_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HASH_02_COUNTER_30_i_2_n_0,
   D => in32_24,
   R => HASH_02_COUNTER_30_i_1_n_0,
   Q => HASH_02_COUNTER_24
);
HASH_02_COUNTER_reg_24_i_1 : CARRY4
 port map (
   CI => HASH_02_COUNTER_reg_20_i_1_n_0,
   CYINIT => '0',
   DI(0) => '0',
   DI(1) => '0',
   DI(2) => '0',
   DI(3) => '0',
   S(0) => HASH_02_COUNTER_21,
   S(1) => HASH_02_COUNTER_22,
   S(2) => HASH_02_COUNTER_23,
   S(3) => HASH_02_COUNTER_24,
   CO(0) => HASH_02_COUNTER_reg_24_i_1_n_3,
   CO(1) => HASH_02_COUNTER_reg_24_i_1_n_2,
   CO(2) => HASH_02_COUNTER_reg_24_i_1_n_1,
   CO(3) => HASH_02_COUNTER_reg_24_i_1_n_0,
   O(0) => in32_21,
   O(1) => in32_22,
   O(2) => in32_23,
   O(3) => in32_24
);
HASH_02_COUNTER_reg_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HASH_02_COUNTER_30_i_2_n_0,
   D => in32_25,
   R => HASH_02_COUNTER_30_i_1_n_0,
   Q => HASH_02_COUNTER_25
);
HASH_02_COUNTER_reg_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HASH_02_COUNTER_30_i_2_n_0,
   D => in32_26,
   R => HASH_02_COUNTER_30_i_1_n_0,
   Q => HASH_02_COUNTER_26
);
HASH_02_COUNTER_reg_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HASH_02_COUNTER_30_i_2_n_0,
   D => in32_27,
   R => HASH_02_COUNTER_30_i_1_n_0,
   Q => HASH_02_COUNTER_27
);
HASH_02_COUNTER_reg_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HASH_02_COUNTER_30_i_2_n_0,
   D => in32_28,
   R => HASH_02_COUNTER_30_i_1_n_0,
   Q => HASH_02_COUNTER_28
);
HASH_02_COUNTER_reg_28_i_1 : CARRY4
 port map (
   CI => HASH_02_COUNTER_reg_24_i_1_n_0,
   CYINIT => '0',
   DI(0) => '0',
   DI(1) => '0',
   DI(2) => '0',
   DI(3) => '0',
   S(0) => HASH_02_COUNTER_25,
   S(1) => HASH_02_COUNTER_26,
   S(2) => HASH_02_COUNTER_27,
   S(3) => HASH_02_COUNTER_28,
   CO(0) => HASH_02_COUNTER_reg_28_i_1_n_3,
   CO(1) => HASH_02_COUNTER_reg_28_i_1_n_2,
   CO(2) => HASH_02_COUNTER_reg_28_i_1_n_1,
   CO(3) => HASH_02_COUNTER_reg_28_i_1_n_0,
   O(0) => in32_25,
   O(1) => in32_26,
   O(2) => in32_27,
   O(3) => in32_28
);
HASH_02_COUNTER_reg_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HASH_02_COUNTER_30_i_2_n_0,
   D => in32_29,
   R => HASH_02_COUNTER_30_i_1_n_0,
   Q => HASH_02_COUNTER_29
);
HASH_02_COUNTER_reg_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HASH_02_COUNTER_30_i_2_n_0,
   D => in32_2,
   R => HASH_02_COUNTER_30_i_1_n_0,
   Q => HASH_02_COUNTER_2
);
HASH_02_COUNTER_reg_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HASH_02_COUNTER_30_i_2_n_0,
   D => in32_30,
   R => HASH_02_COUNTER_30_i_1_n_0,
   Q => HASH_02_COUNTER_30
);
HASH_02_COUNTER_reg_30_i_3 : CARRY4
 port map (
   CI => HASH_02_COUNTER_reg_28_i_1_n_0,
   CYINIT => '0',
   DI(0) => '0',
   DI(1) => '0',
   DI(2) => '0',
   DI(3) => '0',
   S(0) => HASH_02_COUNTER_29,
   S(1) => HASH_02_COUNTER_30,
   S(2) => '0',
   S(3) => '0',
   CO(0) => HASH_02_COUNTER_reg_30_i_3_n_3,
   CO(1) => NLW_HASH_02_COUNTER_reg_30_i_3_CO_UNCONNECTED_1,
   CO(2) => NLW_HASH_02_COUNTER_reg_30_i_3_CO_UNCONNECTED_2,
   CO(3) => NLW_HASH_02_COUNTER_reg_30_i_3_CO_UNCONNECTED_3,
   O(0) => in32_29,
   O(1) => in32_30,
   O(2) => NLW_HASH_02_COUNTER_reg_30_i_3_O_UNCONNECTED_2,
   O(3) => NLW_HASH_02_COUNTER_reg_30_i_3_O_UNCONNECTED_3
);
HASH_02_COUNTER_reg_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HASH_02_COUNTER_30_i_2_n_0,
   D => in32_3,
   R => HASH_02_COUNTER_30_i_1_n_0,
   Q => HASH_02_COUNTER_3
);
HASH_02_COUNTER_reg_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HASH_02_COUNTER_30_i_2_n_0,
   D => in32_4,
   R => HASH_02_COUNTER_30_i_1_n_0,
   Q => HASH_02_COUNTER_4
);
HASH_02_COUNTER_reg_4_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => HASH_02_COUNTER_0,
   DI(0) => '0',
   DI(1) => '0',
   DI(2) => '0',
   DI(3) => '0',
   S(0) => HASH_02_COUNTER_1,
   S(1) => HASH_02_COUNTER_2,
   S(2) => HASH_02_COUNTER_3,
   S(3) => HASH_02_COUNTER_4,
   CO(0) => HASH_02_COUNTER_reg_4_i_1_n_3,
   CO(1) => HASH_02_COUNTER_reg_4_i_1_n_2,
   CO(2) => HASH_02_COUNTER_reg_4_i_1_n_1,
   CO(3) => HASH_02_COUNTER_reg_4_i_1_n_0,
   O(0) => in32_1,
   O(1) => in32_2,
   O(2) => in32_3,
   O(3) => in32_4
);
HASH_02_COUNTER_reg_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HASH_02_COUNTER_30_i_2_n_0,
   D => in32_5,
   R => HASH_02_COUNTER_30_i_1_n_0,
   Q => HASH_02_COUNTER_5
);
HASH_02_COUNTER_reg_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HASH_02_COUNTER_30_i_2_n_0,
   D => in32_6,
   R => HASH_02_COUNTER_30_i_1_n_0,
   Q => HASH_02_COUNTER_6
);
HASH_02_COUNTER_reg_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HASH_02_COUNTER_30_i_2_n_0,
   D => in32_7,
   R => HASH_02_COUNTER_30_i_1_n_0,
   Q => HASH_02_COUNTER_7
);
HASH_02_COUNTER_reg_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HASH_02_COUNTER_30_i_2_n_0,
   D => in32_8,
   R => HASH_02_COUNTER_30_i_1_n_0,
   Q => HASH_02_COUNTER_8
);
HASH_02_COUNTER_reg_8_i_1 : CARRY4
 port map (
   CI => HASH_02_COUNTER_reg_4_i_1_n_0,
   CYINIT => '0',
   DI(0) => '0',
   DI(1) => '0',
   DI(2) => '0',
   DI(3) => '0',
   S(0) => HASH_02_COUNTER_5,
   S(1) => HASH_02_COUNTER_6,
   S(2) => HASH_02_COUNTER_7,
   S(3) => HASH_02_COUNTER_8,
   CO(0) => HASH_02_COUNTER_reg_8_i_1_n_3,
   CO(1) => HASH_02_COUNTER_reg_8_i_1_n_2,
   CO(2) => HASH_02_COUNTER_reg_8_i_1_n_1,
   CO(3) => HASH_02_COUNTER_reg_8_i_1_n_0,
   O(0) => in32_5,
   O(1) => in32_6,
   O(2) => in32_7,
   O(3) => in32_8
);
HASH_02_COUNTER_reg_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HASH_02_COUNTER_30_i_2_n_0,
   D => in32_9,
   R => HASH_02_COUNTER_30_i_1_n_0,
   Q => HASH_02_COUNTER_9
);
HV_0_0_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in23_0,
   O => HV_0_0_i_1_n_0
);
HV_0_10_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in23_10,
   O => HV_0_10_i_1_n_0
);
HV_0_11_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR2_out_2,
   I1 => data_out_OBUF_235,
   O => HV_0_11_i_2_n_0
);
HV_0_11_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR2_out_3,
   I1 => data_out_OBUF_234,
   O => HV_0_11_i_3_n_0
);
HV_0_11_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR2_out_4,
   I1 => data_out_OBUF_233,
   O => HV_0_11_i_4_n_0
);
HV_0_11_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR2_out_5,
   I1 => data_out_OBUF_232,
   O => HV_0_11_i_5_n_0
);
HV_0_12_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR2_out_30,
   I1 => data_out_OBUF_239,
   O => HV_0_12_i_2_n_0
);
HV_0_12_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR2_out_31,
   I1 => data_out_OBUF_238,
   O => HV_0_12_i_3_n_0
);
HV_0_12_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR2_out_32,
   I1 => data_out_OBUF_237,
   O => HV_0_12_i_4_n_0
);
HV_0_12_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR2_out_1,
   I1 => data_out_OBUF_236,
   O => HV_0_12_i_5_n_0
);
HV_0_13_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in23_13,
   O => HV_0_13_i_1_n_0
);
HV_0_14_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in23_14,
   O => HV_0_14_i_1_n_0
);
HV_0_15_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in23_15,
   O => HV_0_15_i_1_n_0
);
HV_0_16_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in23_16,
   O => HV_0_16_i_1_n_0
);
HV_0_18_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR2_out_26,
   I1 => data_out_OBUF_243,
   O => HV_0_18_i_2_n_0
);
HV_0_18_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR2_out_27,
   I1 => data_out_OBUF_242,
   O => HV_0_18_i_3_n_0
);
HV_0_18_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR2_out_28,
   I1 => data_out_OBUF_241,
   O => HV_0_18_i_4_n_0
);
HV_0_18_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR2_out_29,
   I1 => data_out_OBUF_240,
   O => HV_0_18_i_5_n_0
);
HV_0_19_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in23_19,
   O => HV_0_19_i_1_n_0
);
HV_0_1_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in23_1,
   O => HV_0_1_i_1_n_0
);
HV_0_23_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR2_out_22,
   I1 => data_out_OBUF_247,
   O => HV_0_23_i_2_n_0
);
HV_0_23_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR2_out_23,
   I1 => data_out_OBUF_246,
   O => HV_0_23_i_3_n_0
);
HV_0_23_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR2_out_24,
   I1 => data_out_OBUF_245,
   O => HV_0_23_i_4_n_0
);
HV_0_23_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR2_out_25,
   I1 => data_out_OBUF_244,
   O => HV_0_23_i_5_n_0
);
HV_0_25_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in23_25,
   O => HV_0_25_i_1_n_0
);
HV_0_26_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR2_out_18,
   I1 => data_out_OBUF_251,
   O => HV_0_26_i_2_n_0
);
HV_0_26_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR2_out_19,
   I1 => data_out_OBUF_250,
   O => HV_0_26_i_3_n_0
);
HV_0_26_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR2_out_20,
   I1 => data_out_OBUF_249,
   O => HV_0_26_i_4_n_0
);
HV_0_26_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR2_out_21,
   I1 => data_out_OBUF_248,
   O => HV_0_26_i_5_n_0
);
HV_0_27_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in23_27,
   O => HV_0_27_i_1_n_0
);
HV_0_29_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in23_29,
   O => HV_0_29_i_1_n_0
);
HV_0_2_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in23_2,
   O => HV_0_2_i_1_n_0
);
HV_0_30_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in23_30,
   O => HV_0_30_i_1_n_0
);
HV_0_31_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR2_out_14,
   I1 => data_out_OBUF_255,
   O => HV_0_31_i_2_n_0
);
HV_0_31_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR2_out_15,
   I1 => data_out_OBUF_254,
   O => HV_0_31_i_3_n_0
);
HV_0_31_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR2_out_16,
   I1 => data_out_OBUF_253,
   O => HV_0_31_i_4_n_0
);
HV_0_31_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR2_out_17,
   I1 => data_out_OBUF_252,
   O => HV_0_31_i_5_n_0
);
HV_0_3_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR2_out_10,
   I1 => data_out_OBUF_227,
   O => HV_0_3_i_2_n_0
);
HV_0_3_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR2_out_11,
   I1 => data_out_OBUF_226,
   O => HV_0_3_i_3_n_0
);
HV_0_3_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR2_out_12,
   I1 => data_out_OBUF_225,
   O => HV_0_3_i_4_n_0
);
HV_0_3_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR2_out_13,
   I1 => data_out_OBUF_224,
   O => HV_0_3_i_5_n_0
);
HV_0_5_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in23_5,
   O => HV_0_5_i_1_n_0
);
HV_0_6_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in23_6,
   O => HV_0_6_i_1_n_0
);
HV_0_7_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR2_out_6,
   I1 => data_out_OBUF_231,
   O => HV_0_7_i_2_n_0
);
HV_0_7_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR2_out_7,
   I1 => data_out_OBUF_230,
   O => HV_0_7_i_3_n_0
);
HV_0_7_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR2_out_8,
   I1 => data_out_OBUF_229,
   O => HV_0_7_i_4_n_0
);
HV_0_7_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR2_out_9,
   I1 => data_out_OBUF_228,
   O => HV_0_7_i_5_n_0
);
HV_0_9_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in23_9,
   O => HV_0_9_i_1_n_0
);
HV_1_0_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in25_0,
   O => HV_1_0_i_1_n_0
);
HV_1_10_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in25_10,
   O => HV_1_10_i_1_n_0
);
HV_1_11_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in25_11,
   O => HV_1_11_i_1_n_0
);
HV_1_13_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in25_13,
   O => HV_1_13_i_1_n_0
);
HV_1_14_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => b_reg_n_0_15,
   I1 => data_out_OBUF_207,
   O => HV_1_14_i_2_n_0
);
HV_1_14_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => b_reg_n_0_14,
   I1 => data_out_OBUF_206,
   O => HV_1_14_i_3_n_0
);
HV_1_14_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => b_reg_n_0_13,
   I1 => data_out_OBUF_205,
   O => HV_1_14_i_4_n_0
);
HV_1_14_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => b_reg_n_0_12,
   I1 => data_out_OBUF_204,
   O => HV_1_14_i_5_n_0
);
HV_1_15_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in25_15,
   O => HV_1_15_i_1_n_0
);
HV_1_16_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in25_16,
   O => HV_1_16_i_1_n_0
);
HV_1_17_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in25_17,
   O => HV_1_17_i_1_n_0
);
HV_1_18_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in25_18,
   O => HV_1_18_i_1_n_0
);
HV_1_19_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => b_reg_n_0_19,
   I1 => data_out_OBUF_211,
   O => HV_1_19_i_2_n_0
);
HV_1_19_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => b_reg_n_0_18,
   I1 => data_out_OBUF_210,
   O => HV_1_19_i_3_n_0
);
HV_1_19_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => b_reg_n_0_17,
   I1 => data_out_OBUF_209,
   O => HV_1_19_i_4_n_0
);
HV_1_19_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => b_reg_n_0_16,
   I1 => data_out_OBUF_208,
   O => HV_1_19_i_5_n_0
);
HV_1_21_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in25_21,
   O => HV_1_21_i_1_n_0
);
HV_1_22_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in25_22,
   O => HV_1_22_i_1_n_0
);
HV_1_23_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => b_reg_n_0_23,
   I1 => data_out_OBUF_215,
   O => HV_1_23_i_2_n_0
);
HV_1_23_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => b_reg_n_0_22,
   I1 => data_out_OBUF_214,
   O => HV_1_23_i_3_n_0
);
HV_1_23_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => b_reg_n_0_21,
   I1 => data_out_OBUF_213,
   O => HV_1_23_i_4_n_0
);
HV_1_23_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => b_reg_n_0_20,
   I1 => data_out_OBUF_212,
   O => HV_1_23_i_5_n_0
);
HV_1_24_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in25_24,
   O => HV_1_24_i_1_n_0
);
HV_1_25_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in25_25,
   O => HV_1_25_i_1_n_0
);
HV_1_26_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => b_reg_n_0_27,
   I1 => data_out_OBUF_219,
   O => HV_1_26_i_2_n_0
);
HV_1_26_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => b_reg_n_0_26,
   I1 => data_out_OBUF_218,
   O => HV_1_26_i_3_n_0
);
HV_1_26_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => b_reg_n_0_25,
   I1 => data_out_OBUF_217,
   O => HV_1_26_i_4_n_0
);
HV_1_26_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => b_reg_n_0_24,
   I1 => data_out_OBUF_216,
   O => HV_1_26_i_5_n_0
);
HV_1_27_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in25_27,
   O => HV_1_27_i_1_n_0
);
HV_1_28_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in25_28,
   O => HV_1_28_i_1_n_0
);
HV_1_29_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in25_29,
   O => HV_1_29_i_1_n_0
);
HV_1_2_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in25_2,
   O => HV_1_2_i_1_n_0
);
HV_1_30_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => data_out_OBUF_223,
   I1 => b_reg_n_0_31,
   O => HV_1_30_i_2_n_0
);
HV_1_30_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => b_reg_n_0_30,
   I1 => data_out_OBUF_222,
   O => HV_1_30_i_3_n_0
);
HV_1_30_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => b_reg_n_0_29,
   I1 => data_out_OBUF_221,
   O => HV_1_30_i_4_n_0
);
HV_1_30_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => b_reg_n_0_28,
   I1 => data_out_OBUF_220,
   O => HV_1_30_i_5_n_0
);
HV_1_31_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in25_31,
   O => HV_1_31_i_1_n_0
);
HV_1_3_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => b_reg_n_0_3,
   I1 => data_out_OBUF_195,
   O => HV_1_3_i_2_n_0
);
HV_1_3_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => b_reg_n_0_2,
   I1 => data_out_OBUF_194,
   O => HV_1_3_i_3_n_0
);
HV_1_3_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => b_reg_n_0_1,
   I1 => data_out_OBUF_193,
   O => HV_1_3_i_4_n_0
);
HV_1_3_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => b_reg_n_0_0,
   I1 => data_out_OBUF_192,
   O => HV_1_3_i_5_n_0
);
HV_1_6_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => b_reg_n_0_7,
   I1 => data_out_OBUF_199,
   O => HV_1_6_i_2_n_0
);
HV_1_6_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => b_reg_n_0_6,
   I1 => data_out_OBUF_198,
   O => HV_1_6_i_3_n_0
);
HV_1_6_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => b_reg_n_0_5,
   I1 => data_out_OBUF_197,
   O => HV_1_6_i_4_n_0
);
HV_1_6_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => b_reg_n_0_4,
   I1 => data_out_OBUF_196,
   O => HV_1_6_i_5_n_0
);
HV_1_7_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in25_7,
   O => HV_1_7_i_1_n_0
);
HV_1_8_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => b_reg_n_0_11,
   I1 => data_out_OBUF_203,
   O => HV_1_8_i_2_n_0
);
HV_1_8_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => b_reg_n_0_10,
   I1 => data_out_OBUF_202,
   O => HV_1_8_i_3_n_0
);
HV_1_8_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => b_reg_n_0_9,
   I1 => data_out_OBUF_201,
   O => HV_1_8_i_4_n_0
);
HV_1_8_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => b_reg_n_0_8,
   I1 => data_out_OBUF_200,
   O => HV_1_8_i_5_n_0
);
HV_1_9_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in25_9,
   O => HV_1_9_i_1_n_0
);
HV_2_11_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => c_reg_n_0_11,
   I1 => data_out_OBUF_171,
   O => HV_2_11_i_2_n_0
);
HV_2_11_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => c_reg_n_0_10,
   I1 => data_out_OBUF_170,
   O => HV_2_11_i_3_n_0
);
HV_2_11_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => c_reg_n_0_9,
   I1 => data_out_OBUF_169,
   O => HV_2_11_i_4_n_0
);
HV_2_11_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => c_reg_n_0_8,
   I1 => data_out_OBUF_168,
   O => HV_2_11_i_5_n_0
);
HV_2_12_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in26_12,
   O => HV_2_12_i_1_n_0
);
HV_2_13_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in26_13,
   O => HV_2_13_i_1_n_0
);
HV_2_14_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in26_14,
   O => HV_2_14_i_1_n_0
);
HV_2_15_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in26_15,
   O => HV_2_15_i_1_n_0
);
HV_2_16_i_10 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => c_reg_n_0_12,
   I1 => data_out_OBUF_172,
   O => HV_2_16_i_10_n_0
);
HV_2_16_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => c_reg_n_0_19,
   I1 => data_out_OBUF_179,
   O => HV_2_16_i_3_n_0
);
HV_2_16_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => c_reg_n_0_18,
   I1 => data_out_OBUF_178,
   O => HV_2_16_i_4_n_0
);
HV_2_16_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => c_reg_n_0_17,
   I1 => data_out_OBUF_177,
   O => HV_2_16_i_5_n_0
);
HV_2_16_i_6 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => c_reg_n_0_16,
   I1 => data_out_OBUF_176,
   O => HV_2_16_i_6_n_0
);
HV_2_16_i_7 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => c_reg_n_0_15,
   I1 => data_out_OBUF_175,
   O => HV_2_16_i_7_n_0
);
HV_2_16_i_8 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => c_reg_n_0_14,
   I1 => data_out_OBUF_174,
   O => HV_2_16_i_8_n_0
);
HV_2_16_i_9 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => c_reg_n_0_13,
   I1 => data_out_OBUF_173,
   O => HV_2_16_i_9_n_0
);
HV_2_17_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in26_17,
   O => HV_2_17_i_1_n_0
);
HV_2_18_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in26_18,
   O => HV_2_18_i_1_n_0
);
HV_2_19_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in26_19,
   O => HV_2_19_i_1_n_0
);
HV_2_1_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in26_1,
   O => HV_2_1_i_1_n_0
);
HV_2_21_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in26_21,
   O => HV_2_21_i_1_n_0
);
HV_2_22_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in26_22,
   O => HV_2_22_i_1_n_0
);
HV_2_23_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => c_reg_n_0_23,
   I1 => data_out_OBUF_183,
   O => HV_2_23_i_2_n_0
);
HV_2_23_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => c_reg_n_0_22,
   I1 => data_out_OBUF_182,
   O => HV_2_23_i_3_n_0
);
HV_2_23_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => c_reg_n_0_21,
   I1 => data_out_OBUF_181,
   O => HV_2_23_i_4_n_0
);
HV_2_23_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => c_reg_n_0_20,
   I1 => data_out_OBUF_180,
   O => HV_2_23_i_5_n_0
);
HV_2_25_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => c_reg_n_0_27,
   I1 => data_out_OBUF_187,
   O => HV_2_25_i_2_n_0
);
HV_2_25_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => c_reg_n_0_26,
   I1 => data_out_OBUF_186,
   O => HV_2_25_i_3_n_0
);
HV_2_25_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => c_reg_n_0_25,
   I1 => data_out_OBUF_185,
   O => HV_2_25_i_4_n_0
);
HV_2_25_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => c_reg_n_0_24,
   I1 => data_out_OBUF_184,
   O => HV_2_25_i_5_n_0
);
HV_2_26_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in26_26,
   O => HV_2_26_i_1_n_0
);
HV_2_27_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in26_27,
   O => HV_2_27_i_1_n_0
);
HV_2_28_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in26_28,
   O => HV_2_28_i_1_n_0
);
HV_2_29_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in26_29,
   O => HV_2_29_i_1_n_0
);
HV_2_31_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => data_out_OBUF_191,
   I1 => c_reg_n_0_31,
   O => HV_2_31_i_2_n_0
);
HV_2_31_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => c_reg_n_0_30,
   I1 => data_out_OBUF_190,
   O => HV_2_31_i_3_n_0
);
HV_2_31_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => c_reg_n_0_29,
   I1 => data_out_OBUF_189,
   O => HV_2_31_i_4_n_0
);
HV_2_31_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => c_reg_n_0_28,
   I1 => data_out_OBUF_188,
   O => HV_2_31_i_5_n_0
);
HV_2_3_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => c_reg_n_0_3,
   I1 => data_out_OBUF_163,
   O => HV_2_3_i_2_n_0
);
HV_2_3_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => c_reg_n_0_2,
   I1 => data_out_OBUF_162,
   O => HV_2_3_i_3_n_0
);
HV_2_3_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => c_reg_n_0_1,
   I1 => data_out_OBUF_161,
   O => HV_2_3_i_4_n_0
);
HV_2_3_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => c_reg_n_0_0,
   I1 => data_out_OBUF_160,
   O => HV_2_3_i_5_n_0
);
HV_2_4_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in26_4,
   O => HV_2_4_i_1_n_0
);
HV_2_5_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in26_5,
   O => HV_2_5_i_1_n_0
);
HV_2_6_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in26_6,
   O => HV_2_6_i_1_n_0
);
HV_2_7_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => c_reg_n_0_7,
   I1 => data_out_OBUF_167,
   O => HV_2_7_i_2_n_0
);
HV_2_7_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => c_reg_n_0_6,
   I1 => data_out_OBUF_166,
   O => HV_2_7_i_3_n_0
);
HV_2_7_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => c_reg_n_0_5,
   I1 => data_out_OBUF_165,
   O => HV_2_7_i_4_n_0
);
HV_2_7_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => c_reg_n_0_4,
   I1 => data_out_OBUF_164,
   O => HV_2_7_i_5_n_0
);
HV_2_8_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in26_8,
   O => HV_2_8_i_1_n_0
);
HV_2_9_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in26_9,
   O => HV_2_9_i_1_n_0
);
HV_3_10_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in27_10,
   O => HV_3_10_i_1_n_0
);
HV_3_11_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_11,
   I1 => data_out_OBUF_139,
   O => HV_3_11_i_2_n_0
);
HV_3_11_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_10,
   I1 => data_out_OBUF_138,
   O => HV_3_11_i_3_n_0
);
HV_3_11_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_9,
   I1 => data_out_OBUF_137,
   O => HV_3_11_i_4_n_0
);
HV_3_11_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_8,
   I1 => data_out_OBUF_136,
   O => HV_3_11_i_5_n_0
);
HV_3_12_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in27_12,
   O => HV_3_12_i_1_n_0
);
HV_3_13_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in27_13,
   O => HV_3_13_i_1_n_0
);
HV_3_14_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in27_14,
   O => HV_3_14_i_1_n_0
);
HV_3_15_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in27_15,
   O => HV_3_15_i_1_n_0
);
HV_3_15_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_15,
   I1 => data_out_OBUF_143,
   O => HV_3_15_i_3_n_0
);
HV_3_15_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_14,
   I1 => data_out_OBUF_142,
   O => HV_3_15_i_4_n_0
);
HV_3_15_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_13,
   I1 => data_out_OBUF_141,
   O => HV_3_15_i_5_n_0
);
HV_3_15_i_6 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_12,
   I1 => data_out_OBUF_140,
   O => HV_3_15_i_6_n_0
);
HV_3_16_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in27_16,
   O => HV_3_16_i_1_n_0
);
HV_3_17_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in27_17,
   O => HV_3_17_i_1_n_0
);
HV_3_18_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in27_18,
   O => HV_3_18_i_1_n_0
);
HV_3_19_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in27_19,
   O => HV_3_19_i_1_n_0
);
HV_3_1_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in27_1,
   O => HV_3_1_i_1_n_0
);
HV_3_22_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in27_22,
   O => HV_3_22_i_1_n_0
);
HV_3_23_i_10 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_16,
   I1 => data_out_OBUF_144,
   O => HV_3_23_i_10_n_0
);
HV_3_23_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_23,
   I1 => data_out_OBUF_151,
   O => HV_3_23_i_3_n_0
);
HV_3_23_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_22,
   I1 => data_out_OBUF_150,
   O => HV_3_23_i_4_n_0
);
HV_3_23_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_21,
   I1 => data_out_OBUF_149,
   O => HV_3_23_i_5_n_0
);
HV_3_23_i_6 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_20,
   I1 => data_out_OBUF_148,
   O => HV_3_23_i_6_n_0
);
HV_3_23_i_7 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_19,
   I1 => data_out_OBUF_147,
   O => HV_3_23_i_7_n_0
);
HV_3_23_i_8 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_18,
   I1 => data_out_OBUF_146,
   O => HV_3_23_i_8_n_0
);
HV_3_23_i_9 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_17,
   I1 => data_out_OBUF_145,
   O => HV_3_23_i_9_n_0
);
HV_3_24_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in27_24,
   O => HV_3_24_i_1_n_0
);
HV_3_26_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in27_26,
   O => HV_3_26_i_1_n_0
);
HV_3_27_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_27,
   I1 => data_out_OBUF_155,
   O => HV_3_27_i_2_n_0
);
HV_3_27_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_26,
   I1 => data_out_OBUF_154,
   O => HV_3_27_i_3_n_0
);
HV_3_27_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_25,
   I1 => data_out_OBUF_153,
   O => HV_3_27_i_4_n_0
);
HV_3_27_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_24,
   I1 => data_out_OBUF_152,
   O => HV_3_27_i_5_n_0
);
HV_3_29_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in27_29,
   O => HV_3_29_i_1_n_0
);
HV_3_2_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_3,
   I1 => data_out_OBUF_131,
   O => HV_3_2_i_2_n_0
);
HV_3_2_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_2,
   I1 => data_out_OBUF_130,
   O => HV_3_2_i_3_n_0
);
HV_3_2_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_1,
   I1 => data_out_OBUF_129,
   O => HV_3_2_i_4_n_0
);
HV_3_2_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_0,
   I1 => data_out_OBUF_128,
   O => HV_3_2_i_5_n_0
);
HV_3_30_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => data_out_OBUF_159,
   I1 => d_31,
   O => HV_3_30_i_2_n_0
);
HV_3_30_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_30,
   I1 => data_out_OBUF_158,
   O => HV_3_30_i_3_n_0
);
HV_3_30_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_29,
   I1 => data_out_OBUF_157,
   O => HV_3_30_i_4_n_0
);
HV_3_30_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_28,
   I1 => data_out_OBUF_156,
   O => HV_3_30_i_5_n_0
);
HV_3_31_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in27_31,
   O => HV_3_31_i_1_n_0
);
HV_3_3_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in27_3,
   O => HV_3_3_i_1_n_0
);
HV_3_4_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in27_4,
   O => HV_3_4_i_1_n_0
);
HV_3_5_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in27_5,
   O => HV_3_5_i_1_n_0
);
HV_3_7_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_7,
   I1 => data_out_OBUF_135,
   O => HV_3_7_i_2_n_0
);
HV_3_7_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_6,
   I1 => data_out_OBUF_134,
   O => HV_3_7_i_3_n_0
);
HV_3_7_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_5,
   I1 => data_out_OBUF_133,
   O => HV_3_7_i_4_n_0
);
HV_3_7_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => d_4,
   I1 => data_out_OBUF_132,
   O => HV_3_7_i_5_n_0
);
HV_3_8_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in27_8,
   O => HV_3_8_i_1_n_0
);
HV_4_0_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in28_0,
   O => HV_4_0_i_1_n_0
);
HV_4_11_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR11_out_32,
   I1 => data_out_OBUF_107,
   O => HV_4_11_i_2_n_0
);
HV_4_11_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR11_out_1,
   I1 => data_out_OBUF_106,
   O => HV_4_11_i_3_n_0
);
HV_4_11_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR11_out_2,
   I1 => data_out_OBUF_105,
   O => HV_4_11_i_4_n_0
);
HV_4_11_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR11_out_3,
   I1 => data_out_OBUF_104,
   O => HV_4_11_i_5_n_0
);
HV_4_12_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in28_12,
   O => HV_4_12_i_1_n_0
);
HV_4_14_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in28_14,
   O => HV_4_14_i_1_n_0
);
HV_4_15_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR11_out_28,
   I1 => data_out_OBUF_111,
   O => HV_4_15_i_2_n_0
);
HV_4_15_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR11_out_29,
   I1 => data_out_OBUF_110,
   O => HV_4_15_i_3_n_0
);
HV_4_15_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR11_out_30,
   I1 => data_out_OBUF_109,
   O => HV_4_15_i_4_n_0
);
HV_4_15_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR11_out_31,
   I1 => data_out_OBUF_108,
   O => HV_4_15_i_5_n_0
);
HV_4_16_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR11_out_24,
   I1 => data_out_OBUF_115,
   O => HV_4_16_i_2_n_0
);
HV_4_16_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR11_out_25,
   I1 => data_out_OBUF_114,
   O => HV_4_16_i_3_n_0
);
HV_4_16_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR11_out_26,
   I1 => data_out_OBUF_113,
   O => HV_4_16_i_4_n_0
);
HV_4_16_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR11_out_27,
   I1 => data_out_OBUF_112,
   O => HV_4_16_i_5_n_0
);
HV_4_17_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in28_17,
   O => HV_4_17_i_1_n_0
);
HV_4_18_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in28_18,
   O => HV_4_18_i_1_n_0
);
HV_4_19_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in28_19,
   O => HV_4_19_i_1_n_0
);
HV_4_1_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in28_1,
   O => HV_4_1_i_1_n_0
);
HV_4_23_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR11_out_20,
   I1 => data_out_OBUF_119,
   O => HV_4_23_i_2_n_0
);
HV_4_23_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR11_out_21,
   I1 => data_out_OBUF_118,
   O => HV_4_23_i_3_n_0
);
HV_4_23_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR11_out_22,
   I1 => data_out_OBUF_117,
   O => HV_4_23_i_4_n_0
);
HV_4_23_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR11_out_23,
   I1 => data_out_OBUF_116,
   O => HV_4_23_i_5_n_0
);
HV_4_24_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in28_24,
   O => HV_4_24_i_1_n_0
);
HV_4_27_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR11_out_16,
   I1 => data_out_OBUF_123,
   O => HV_4_27_i_2_n_0
);
HV_4_27_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR11_out_17,
   I1 => data_out_OBUF_122,
   O => HV_4_27_i_3_n_0
);
HV_4_27_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR11_out_18,
   I1 => data_out_OBUF_121,
   O => HV_4_27_i_4_n_0
);
HV_4_27_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR11_out_19,
   I1 => data_out_OBUF_120,
   O => HV_4_27_i_5_n_0
);
HV_4_28_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in28_28,
   O => HV_4_28_i_1_n_0
);
HV_4_2_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in28_2,
   O => HV_4_2_i_1_n_0
);
HV_4_30_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in28_30,
   O => HV_4_30_i_1_n_0
);
HV_4_31_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => data_out_OBUF_127,
   I1 => ROTR11_out_12,
   O => HV_4_31_i_2_n_0
);
HV_4_31_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR11_out_13,
   I1 => data_out_OBUF_126,
   O => HV_4_31_i_3_n_0
);
HV_4_31_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR11_out_14,
   I1 => data_out_OBUF_125,
   O => HV_4_31_i_4_n_0
);
HV_4_31_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR11_out_15,
   I1 => data_out_OBUF_124,
   O => HV_4_31_i_5_n_0
);
HV_4_3_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in28_3,
   O => HV_4_3_i_1_n_0
);
HV_4_4_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in28_4,
   O => HV_4_4_i_1_n_0
);
HV_4_5_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in28_5,
   O => HV_4_5_i_1_n_0
);
HV_4_6_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in28_6,
   O => HV_4_6_i_1_n_0
);
HV_4_7_i_10 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR11_out_11,
   I1 => data_out_OBUF_96,
   O => HV_4_7_i_10_n_0
);
HV_4_7_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR11_out_4,
   I1 => data_out_OBUF_103,
   O => HV_4_7_i_3_n_0
);
HV_4_7_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR11_out_5,
   I1 => data_out_OBUF_102,
   O => HV_4_7_i_4_n_0
);
HV_4_7_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR11_out_6,
   I1 => data_out_OBUF_101,
   O => HV_4_7_i_5_n_0
);
HV_4_7_i_6 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR11_out_7,
   I1 => data_out_OBUF_100,
   O => HV_4_7_i_6_n_0
);
HV_4_7_i_7 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR11_out_8,
   I1 => data_out_OBUF_99,
   O => HV_4_7_i_7_n_0
);
HV_4_7_i_8 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR11_out_9,
   I1 => data_out_OBUF_98,
   O => HV_4_7_i_8_n_0
);
HV_4_7_i_9 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => ROTR11_out_10,
   I1 => data_out_OBUF_97,
   O => HV_4_7_i_9_n_0
);
HV_4_9_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in28_9,
   O => HV_4_9_i_1_n_0
);
HV_5_10_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => f_reg_n_0_11,
   I1 => data_out_OBUF_75,
   O => HV_5_10_i_2_n_0
);
HV_5_10_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => f_reg_n_0_10,
   I1 => data_out_OBUF_74,
   O => HV_5_10_i_3_n_0
);
HV_5_10_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => f_reg_n_0_9,
   I1 => data_out_OBUF_73,
   O => HV_5_10_i_4_n_0
);
HV_5_10_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => f_reg_n_0_8,
   I1 => data_out_OBUF_72,
   O => HV_5_10_i_5_n_0
);
HV_5_11_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in29_11,
   O => HV_5_11_i_1_n_0
);
HV_5_13_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in29_13,
   O => HV_5_13_i_1_n_0
);
HV_5_14_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in29_14,
   O => HV_5_14_i_1_n_0
);
HV_5_15_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => f_reg_n_0_15,
   I1 => data_out_OBUF_79,
   O => HV_5_15_i_2_n_0
);
HV_5_15_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => f_reg_n_0_14,
   I1 => data_out_OBUF_78,
   O => HV_5_15_i_3_n_0
);
HV_5_15_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => f_reg_n_0_13,
   I1 => data_out_OBUF_77,
   O => HV_5_15_i_4_n_0
);
HV_5_15_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => f_reg_n_0_12,
   I1 => data_out_OBUF_76,
   O => HV_5_15_i_5_n_0
);
HV_5_16_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in29_16,
   O => HV_5_16_i_1_n_0
);
HV_5_18_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in29_18,
   O => HV_5_18_i_1_n_0
);
HV_5_19_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => f_reg_n_0_19,
   I1 => data_out_OBUF_83,
   O => HV_5_19_i_2_n_0
);
HV_5_19_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => f_reg_n_0_18,
   I1 => data_out_OBUF_82,
   O => HV_5_19_i_3_n_0
);
HV_5_19_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => f_reg_n_0_17,
   I1 => data_out_OBUF_81,
   O => HV_5_19_i_4_n_0
);
HV_5_19_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => f_reg_n_0_16,
   I1 => data_out_OBUF_80,
   O => HV_5_19_i_5_n_0
);
HV_5_1_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => f_reg_n_0_3,
   I1 => data_out_OBUF_67,
   O => HV_5_1_i_2_n_0
);
HV_5_1_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => f_reg_n_0_2,
   I1 => data_out_OBUF_66,
   O => HV_5_1_i_3_n_0
);
HV_5_1_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => f_reg_n_0_1,
   I1 => data_out_OBUF_65,
   O => HV_5_1_i_4_n_0
);
HV_5_1_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => f_reg_n_0_0,
   I1 => data_out_OBUF_64,
   O => HV_5_1_i_5_n_0
);
HV_5_23_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => f_reg_n_0_23,
   I1 => data_out_OBUF_87,
   O => HV_5_23_i_2_n_0
);
HV_5_23_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => f_reg_n_0_22,
   I1 => data_out_OBUF_86,
   O => HV_5_23_i_3_n_0
);
HV_5_23_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => f_reg_n_0_21,
   I1 => data_out_OBUF_85,
   O => HV_5_23_i_4_n_0
);
HV_5_23_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => f_reg_n_0_20,
   I1 => data_out_OBUF_84,
   O => HV_5_23_i_5_n_0
);
HV_5_24_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in29_24,
   O => HV_5_24_i_1_n_0
);
HV_5_25_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in29_25,
   O => HV_5_25_i_1_n_0
);
HV_5_26_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => f_reg_n_0_27,
   I1 => data_out_OBUF_91,
   O => HV_5_26_i_2_n_0
);
HV_5_26_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => f_reg_n_0_26,
   I1 => data_out_OBUF_90,
   O => HV_5_26_i_3_n_0
);
HV_5_26_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => f_reg_n_0_25,
   I1 => data_out_OBUF_89,
   O => HV_5_26_i_4_n_0
);
HV_5_26_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => f_reg_n_0_24,
   I1 => data_out_OBUF_88,
   O => HV_5_26_i_5_n_0
);
HV_5_27_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in29_27,
   O => HV_5_27_i_1_n_0
);
HV_5_28_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in29_28,
   O => HV_5_28_i_1_n_0
);
HV_5_2_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in29_2,
   O => HV_5_2_i_1_n_0
);
HV_5_30_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => data_out_OBUF_95,
   I1 => f_reg_n_0_31,
   O => HV_5_30_i_2_n_0
);
HV_5_30_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => f_reg_n_0_30,
   I1 => data_out_OBUF_94,
   O => HV_5_30_i_3_n_0
);
HV_5_30_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => f_reg_n_0_29,
   I1 => data_out_OBUF_93,
   O => HV_5_30_i_4_n_0
);
HV_5_30_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => f_reg_n_0_28,
   I1 => data_out_OBUF_92,
   O => HV_5_30_i_5_n_0
);
HV_5_31_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in29_31,
   O => HV_5_31_i_1_n_0
);
HV_5_3_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in29_3,
   O => HV_5_3_i_1_n_0
);
HV_5_6_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => f_reg_n_0_7,
   I1 => data_out_OBUF_71,
   O => HV_5_6_i_2_n_0
);
HV_5_6_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => f_reg_n_0_6,
   I1 => data_out_OBUF_70,
   O => HV_5_6_i_3_n_0
);
HV_5_6_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => f_reg_n_0_5,
   I1 => data_out_OBUF_69,
   O => HV_5_6_i_4_n_0
);
HV_5_6_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => f_reg_n_0_4,
   I1 => data_out_OBUF_68,
   O => HV_5_6_i_5_n_0
);
HV_5_7_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in29_7,
   O => HV_5_7_i_1_n_0
);
HV_6_0_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in30_0,
   O => HV_6_0_i_1_n_0
);
HV_6_10_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => g_reg_n_0_11,
   I1 => data_out_OBUF_43,
   O => HV_6_10_i_2_n_0
);
HV_6_10_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => g_reg_n_0_10,
   I1 => data_out_OBUF_42,
   O => HV_6_10_i_3_n_0
);
HV_6_10_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => g_reg_n_0_9,
   I1 => data_out_OBUF_41,
   O => HV_6_10_i_4_n_0
);
HV_6_10_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => g_reg_n_0_8,
   I1 => data_out_OBUF_40,
   O => HV_6_10_i_5_n_0
);
HV_6_11_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in30_11,
   O => HV_6_11_i_1_n_0
);
HV_6_12_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in30_12,
   O => HV_6_12_i_1_n_0
);
HV_6_13_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => g_reg_n_0_15,
   I1 => data_out_OBUF_47,
   O => HV_6_13_i_2_n_0
);
HV_6_13_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => g_reg_n_0_14,
   I1 => data_out_OBUF_46,
   O => HV_6_13_i_3_n_0
);
HV_6_13_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => g_reg_n_0_13,
   I1 => data_out_OBUF_45,
   O => HV_6_13_i_4_n_0
);
HV_6_13_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => g_reg_n_0_12,
   I1 => data_out_OBUF_44,
   O => HV_6_13_i_5_n_0
);
HV_6_14_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in30_14,
   O => HV_6_14_i_1_n_0
);
HV_6_15_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in30_15,
   O => HV_6_15_i_1_n_0
);
HV_6_16_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in30_16,
   O => HV_6_16_i_1_n_0
);
HV_6_17_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in30_17,
   O => HV_6_17_i_1_n_0
);
HV_6_19_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => g_reg_n_0_19,
   I1 => data_out_OBUF_51,
   O => HV_6_19_i_2_n_0
);
HV_6_19_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => g_reg_n_0_18,
   I1 => data_out_OBUF_50,
   O => HV_6_19_i_3_n_0
);
HV_6_19_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => g_reg_n_0_17,
   I1 => data_out_OBUF_49,
   O => HV_6_19_i_4_n_0
);
HV_6_19_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => g_reg_n_0_16,
   I1 => data_out_OBUF_48,
   O => HV_6_19_i_5_n_0
);
HV_6_1_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in30_1,
   O => HV_6_1_i_1_n_0
);
HV_6_22_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => g_reg_n_0_23,
   I1 => data_out_OBUF_55,
   O => HV_6_22_i_2_n_0
);
HV_6_22_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => g_reg_n_0_22,
   I1 => data_out_OBUF_54,
   O => HV_6_22_i_3_n_0
);
HV_6_22_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => g_reg_n_0_21,
   I1 => data_out_OBUF_53,
   O => HV_6_22_i_4_n_0
);
HV_6_22_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => g_reg_n_0_20,
   I1 => data_out_OBUF_52,
   O => HV_6_22_i_5_n_0
);
HV_6_23_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in30_23,
   O => HV_6_23_i_1_n_0
);
HV_6_24_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in30_24,
   O => HV_6_24_i_1_n_0
);
HV_6_25_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in30_25,
   O => HV_6_25_i_1_n_0
);
HV_6_26_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in30_26,
   O => HV_6_26_i_1_n_0
);
HV_6_27_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in30_27,
   O => HV_6_27_i_1_n_0
);
HV_6_28_i_1 : LUT3
  generic map(
   INIT => X"32"
  )
 port map (
   I0 => M_0,
   I1 => rst_IBUF,
   I2 => FSM_onehot_CURRENT_STATE_reg_n_0_0,
   O => HV_6_28_i_1_n_0
);
HV_6_28_i_2 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in30_28,
   O => HV_6_28_i_2_n_0
);
HV_6_2_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => g_reg_n_0_3,
   I1 => data_out_OBUF_35,
   O => HV_6_2_i_2_n_0
);
HV_6_2_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => g_reg_n_0_2,
   I1 => data_out_OBUF_34,
   O => HV_6_2_i_3_n_0
);
HV_6_2_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => g_reg_n_0_1,
   I1 => data_out_OBUF_33,
   O => HV_6_2_i_4_n_0
);
HV_6_2_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => g_reg_n_0_0,
   I1 => data_out_OBUF_32,
   O => HV_6_2_i_5_n_0
);
HV_6_31_i_1 : LUT4
  generic map(
   INIT => X"0302"
  )
 port map (
   I0 => M_0,
   I1 => rst_IBUF,
   I2 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_0,
   O => HV_6_31_i_1_n_0
);
HV_6_31_i_10 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => g_reg_n_0_26,
   I1 => data_out_OBUF_58,
   O => HV_6_31_i_10_n_0
);
HV_6_31_i_11 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => g_reg_n_0_25,
   I1 => data_out_OBUF_57,
   O => HV_6_31_i_11_n_0
);
HV_6_31_i_12 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => g_reg_n_0_24,
   I1 => data_out_OBUF_56,
   O => HV_6_31_i_12_n_0
);
HV_6_31_i_2 : LUT4
  generic map(
   INIT => X"3332"
  )
 port map (
   I0 => M_0,
   I1 => rst_IBUF,
   I2 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_0,
   O => HV_reg_0_0
);
HV_6_31_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => data_out_OBUF_63,
   I1 => g_reg_n_0_31,
   O => HV_6_31_i_5_n_0
);
HV_6_31_i_6 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => g_reg_n_0_30,
   I1 => data_out_OBUF_62,
   O => HV_6_31_i_6_n_0
);
HV_6_31_i_7 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => g_reg_n_0_29,
   I1 => data_out_OBUF_61,
   O => HV_6_31_i_7_n_0
);
HV_6_31_i_8 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => g_reg_n_0_28,
   I1 => data_out_OBUF_60,
   O => HV_6_31_i_8_n_0
);
HV_6_31_i_9 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => g_reg_n_0_27,
   I1 => data_out_OBUF_59,
   O => HV_6_31_i_9_n_0
);
HV_6_3_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in30_3,
   O => HV_6_3_i_1_n_0
);
HV_6_5_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in30_5,
   O => HV_6_5_i_1_n_0
);
HV_6_6_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => g_reg_n_0_7,
   I1 => data_out_OBUF_39,
   O => HV_6_6_i_2_n_0
);
HV_6_6_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => g_reg_n_0_6,
   I1 => data_out_OBUF_38,
   O => HV_6_6_i_3_n_0
);
HV_6_6_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => g_reg_n_0_5,
   I1 => data_out_OBUF_37,
   O => HV_6_6_i_4_n_0
);
HV_6_6_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => g_reg_n_0_4,
   I1 => data_out_OBUF_36,
   O => HV_6_6_i_5_n_0
);
HV_6_7_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in30_7,
   O => HV_6_7_i_1_n_0
);
HV_6_8_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in30_8,
   O => HV_6_8_i_1_n_0
);
HV_7_0_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in31_0,
   O => HV_7_0_i_1_n_0
);
HV_7_10_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in31_10,
   O => HV_7_10_i_1_n_0
);
HV_7_11_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in31_11,
   O => HV_7_11_i_1_n_0
);
HV_7_13_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => h_15,
   I1 => data_out_OBUF_15,
   O => HV_7_13_i_2_n_0
);
HV_7_13_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => h_14,
   I1 => data_out_OBUF_14,
   O => HV_7_13_i_3_n_0
);
HV_7_13_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => h_13,
   I1 => data_out_OBUF_13,
   O => HV_7_13_i_4_n_0
);
HV_7_13_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => h_12,
   I1 => data_out_OBUF_12,
   O => HV_7_13_i_5_n_0
);
HV_7_14_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in31_14,
   O => HV_7_14_i_1_n_0
);
HV_7_15_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in31_15,
   O => HV_7_15_i_1_n_0
);
HV_7_19_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => h_19,
   I1 => data_out_OBUF_19,
   O => HV_7_19_i_2_n_0
);
HV_7_19_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => h_18,
   I1 => data_out_OBUF_18,
   O => HV_7_19_i_3_n_0
);
HV_7_19_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => h_17,
   I1 => data_out_OBUF_17,
   O => HV_7_19_i_4_n_0
);
HV_7_19_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => h_16,
   I1 => data_out_OBUF_16,
   O => HV_7_19_i_5_n_0
);
HV_7_20_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => h_23,
   I1 => data_out_OBUF_23,
   O => HV_7_20_i_2_n_0
);
HV_7_20_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => h_22,
   I1 => data_out_OBUF_22,
   O => HV_7_20_i_3_n_0
);
HV_7_20_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => h_21,
   I1 => data_out_OBUF_21,
   O => HV_7_20_i_4_n_0
);
HV_7_20_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => h_20,
   I1 => data_out_OBUF_20,
   O => HV_7_20_i_5_n_0
);
HV_7_21_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in31_21,
   O => HV_7_21_i_1_n_0
);
HV_7_22_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in31_22,
   O => HV_7_22_i_1_n_0
);
HV_7_23_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in31_23,
   O => HV_7_23_i_1_n_0
);
HV_7_24_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in31_24,
   O => HV_7_24_i_1_n_0
);
HV_7_25_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in31_25,
   O => HV_7_25_i_1_n_0
);
HV_7_26_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => h_27,
   I1 => data_out_OBUF_27,
   O => HV_7_26_i_2_n_0
);
HV_7_26_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => h_26,
   I1 => data_out_OBUF_26,
   O => HV_7_26_i_3_n_0
);
HV_7_26_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => h_25,
   I1 => data_out_OBUF_25,
   O => HV_7_26_i_4_n_0
);
HV_7_26_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => h_24,
   I1 => data_out_OBUF_24,
   O => HV_7_26_i_5_n_0
);
HV_7_27_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in31_27,
   O => HV_7_27_i_1_n_0
);
HV_7_28_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in31_28,
   O => HV_7_28_i_1_n_0
);
HV_7_2_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => h_3,
   I1 => data_out_OBUF_3,
   O => HV_7_2_i_2_n_0
);
HV_7_2_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => h_2,
   I1 => data_out_OBUF_2,
   O => HV_7_2_i_3_n_0
);
HV_7_2_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => h_1,
   I1 => data_out_OBUF_1,
   O => HV_7_2_i_4_n_0
);
HV_7_2_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => h_0,
   I1 => data_out_OBUF_0,
   O => HV_7_2_i_5_n_0
);
HV_7_30_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in31_30,
   O => HV_7_30_i_1_n_0
);
HV_7_31_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => h_31,
   I1 => data_out_OBUF_31,
   O => HV_7_31_i_2_n_0
);
HV_7_31_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => h_30,
   I1 => data_out_OBUF_30,
   O => HV_7_31_i_3_n_0
);
HV_7_31_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => h_29,
   I1 => data_out_OBUF_29,
   O => HV_7_31_i_4_n_0
);
HV_7_31_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => h_28,
   I1 => data_out_OBUF_28,
   O => HV_7_31_i_5_n_0
);
HV_7_3_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in31_3,
   O => HV_7_3_i_1_n_0
);
HV_7_4_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in31_4,
   O => HV_7_4_i_1_n_0
);
HV_7_7_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => h_7,
   I1 => data_out_OBUF_7,
   O => HV_7_7_i_2_n_0
);
HV_7_7_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => h_6,
   I1 => data_out_OBUF_6,
   O => HV_7_7_i_3_n_0
);
HV_7_7_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => h_5,
   I1 => data_out_OBUF_5,
   O => HV_7_7_i_4_n_0
);
HV_7_7_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => h_4,
   I1 => data_out_OBUF_4,
   O => HV_7_7_i_5_n_0
);
HV_7_8_i_1 : LUT2
  generic map(
   INIT => X"8"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_9,
   I1 => in31_8,
   O => HV_7_8_i_1_n_0
);
HV_7_9_i_2 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => h_11,
   I1 => data_out_OBUF_11,
   O => HV_7_9_i_2_n_0
);
HV_7_9_i_3 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => h_10,
   I1 => data_out_OBUF_10,
   O => HV_7_9_i_3_n_0
);
HV_7_9_i_4 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => h_9,
   I1 => data_out_OBUF_9,
   O => HV_7_9_i_4_n_0
);
HV_7_9_i_5 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => h_8,
   I1 => data_out_OBUF_8,
   O => HV_7_9_i_5_n_0
);
HV_reg_0_0 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_0_0_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_224
);
HV_reg_0_10 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_0_10_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_234
);
HV_reg_0_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in23_11,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_235
);
HV_reg_0_11_i_1 : CARRY4
 port map (
   CI => HV_reg_0_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => ROTR2_out_5,
   DI(1) => ROTR2_out_4,
   DI(2) => ROTR2_out_3,
   DI(3) => ROTR2_out_2,
   S(0) => HV_0_11_i_5_n_0,
   S(1) => HV_0_11_i_4_n_0,
   S(2) => HV_0_11_i_3_n_0,
   S(3) => HV_0_11_i_2_n_0,
   CO(0) => HV_reg_0_11_i_1_n_3,
   CO(1) => HV_reg_0_11_i_1_n_2,
   CO(2) => HV_reg_0_11_i_1_n_1,
   CO(3) => HV_reg_0_11_i_1_n_0,
   O(0) => in23_8,
   O(1) => in23_9,
   O(2) => in23_10,
   O(3) => in23_11
);
HV_reg_0_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in23_12,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_236
);
HV_reg_0_12_i_1 : CARRY4
 port map (
   CI => HV_reg_0_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => ROTR2_out_1,
   DI(1) => ROTR2_out_32,
   DI(2) => ROTR2_out_31,
   DI(3) => ROTR2_out_30,
   S(0) => HV_0_12_i_5_n_0,
   S(1) => HV_0_12_i_4_n_0,
   S(2) => HV_0_12_i_3_n_0,
   S(3) => HV_0_12_i_2_n_0,
   CO(0) => HV_reg_0_12_i_1_n_3,
   CO(1) => HV_reg_0_12_i_1_n_2,
   CO(2) => HV_reg_0_12_i_1_n_1,
   CO(3) => HV_reg_0_12_i_1_n_0,
   O(0) => in23_12,
   O(1) => in23_13,
   O(2) => in23_14,
   O(3) => in23_15
);
HV_reg_0_13 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_0_13_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_237
);
HV_reg_0_14 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_0_14_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_238
);
HV_reg_0_15 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_0_15_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_239
);
HV_reg_0_16 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_0_16_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_240
);
HV_reg_0_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in23_17,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_241
);
HV_reg_0_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in23_18,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_242
);
HV_reg_0_18_i_1 : CARRY4
 port map (
   CI => HV_reg_0_12_i_1_n_0,
   CYINIT => '0',
   DI(0) => ROTR2_out_29,
   DI(1) => ROTR2_out_28,
   DI(2) => ROTR2_out_27,
   DI(3) => ROTR2_out_26,
   S(0) => HV_0_18_i_5_n_0,
   S(1) => HV_0_18_i_4_n_0,
   S(2) => HV_0_18_i_3_n_0,
   S(3) => HV_0_18_i_2_n_0,
   CO(0) => HV_reg_0_18_i_1_n_3,
   CO(1) => HV_reg_0_18_i_1_n_2,
   CO(2) => HV_reg_0_18_i_1_n_1,
   CO(3) => HV_reg_0_18_i_1_n_0,
   O(0) => in23_16,
   O(1) => in23_17,
   O(2) => in23_18,
   O(3) => in23_19
);
HV_reg_0_19 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_0_19_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_243
);
HV_reg_0_1 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_0_1_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_225
);
HV_reg_0_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in23_20,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_244
);
HV_reg_0_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in23_21,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_245
);
HV_reg_0_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in23_22,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_246
);
HV_reg_0_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in23_23,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_247
);
HV_reg_0_23_i_1 : CARRY4
 port map (
   CI => HV_reg_0_18_i_1_n_0,
   CYINIT => '0',
   DI(0) => ROTR2_out_25,
   DI(1) => ROTR2_out_24,
   DI(2) => ROTR2_out_23,
   DI(3) => ROTR2_out_22,
   S(0) => HV_0_23_i_5_n_0,
   S(1) => HV_0_23_i_4_n_0,
   S(2) => HV_0_23_i_3_n_0,
   S(3) => HV_0_23_i_2_n_0,
   CO(0) => HV_reg_0_23_i_1_n_3,
   CO(1) => HV_reg_0_23_i_1_n_2,
   CO(2) => HV_reg_0_23_i_1_n_1,
   CO(3) => HV_reg_0_23_i_1_n_0,
   O(0) => in23_20,
   O(1) => in23_21,
   O(2) => in23_22,
   O(3) => in23_23
);
HV_reg_0_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in23_24,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_248
);
HV_reg_0_25 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_0_25_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_249
);
HV_reg_0_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in23_26,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_250
);
HV_reg_0_26_i_1 : CARRY4
 port map (
   CI => HV_reg_0_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => ROTR2_out_21,
   DI(1) => ROTR2_out_20,
   DI(2) => ROTR2_out_19,
   DI(3) => ROTR2_out_18,
   S(0) => HV_0_26_i_5_n_0,
   S(1) => HV_0_26_i_4_n_0,
   S(2) => HV_0_26_i_3_n_0,
   S(3) => HV_0_26_i_2_n_0,
   CO(0) => HV_reg_0_26_i_1_n_3,
   CO(1) => HV_reg_0_26_i_1_n_2,
   CO(2) => HV_reg_0_26_i_1_n_1,
   CO(3) => HV_reg_0_26_i_1_n_0,
   O(0) => in23_24,
   O(1) => in23_25,
   O(2) => in23_26,
   O(3) => in23_27
);
HV_reg_0_27 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_0_27_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_251
);
HV_reg_0_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in23_28,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_252
);
HV_reg_0_29 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_0_29_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_253
);
HV_reg_0_2 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_0_2_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_226
);
HV_reg_0_30 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_0_30_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_254
);
HV_reg_0_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in23_31,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_255
);
HV_reg_0_31_i_1 : CARRY4
 port map (
   CI => HV_reg_0_26_i_1_n_0,
   CYINIT => '0',
   DI(0) => ROTR2_out_17,
   DI(1) => ROTR2_out_16,
   DI(2) => ROTR2_out_15,
   DI(3) => '0',
   S(0) => HV_0_31_i_5_n_0,
   S(1) => HV_0_31_i_4_n_0,
   S(2) => HV_0_31_i_3_n_0,
   S(3) => HV_0_31_i_2_n_0,
   CO(0) => HV_reg_0_31_i_1_n_3,
   CO(1) => HV_reg_0_31_i_1_n_2,
   CO(2) => HV_reg_0_31_i_1_n_1,
   CO(3) => NLW_HV_reg_0_31_i_1_CO_UNCONNECTED_3,
   O(0) => in23_28,
   O(1) => in23_29,
   O(2) => in23_30,
   O(3) => in23_31
);
HV_reg_0_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in23_3,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_227
);
HV_reg_0_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => ROTR2_out_13,
   DI(1) => ROTR2_out_12,
   DI(2) => ROTR2_out_11,
   DI(3) => ROTR2_out_10,
   S(0) => HV_0_3_i_5_n_0,
   S(1) => HV_0_3_i_4_n_0,
   S(2) => HV_0_3_i_3_n_0,
   S(3) => HV_0_3_i_2_n_0,
   CO(0) => HV_reg_0_3_i_1_n_3,
   CO(1) => HV_reg_0_3_i_1_n_2,
   CO(2) => HV_reg_0_3_i_1_n_1,
   CO(3) => HV_reg_0_3_i_1_n_0,
   O(0) => in23_0,
   O(1) => in23_1,
   O(2) => in23_2,
   O(3) => in23_3
);
HV_reg_0_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in23_4,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_228
);
HV_reg_0_5 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_0_5_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_229
);
HV_reg_0_6 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_0_6_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_230
);
HV_reg_0_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in23_7,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_231
);
HV_reg_0_7_i_1 : CARRY4
 port map (
   CI => HV_reg_0_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => ROTR2_out_9,
   DI(1) => ROTR2_out_8,
   DI(2) => ROTR2_out_7,
   DI(3) => ROTR2_out_6,
   S(0) => HV_0_7_i_5_n_0,
   S(1) => HV_0_7_i_4_n_0,
   S(2) => HV_0_7_i_3_n_0,
   S(3) => HV_0_7_i_2_n_0,
   CO(0) => HV_reg_0_7_i_1_n_3,
   CO(1) => HV_reg_0_7_i_1_n_2,
   CO(2) => HV_reg_0_7_i_1_n_1,
   CO(3) => HV_reg_0_7_i_1_n_0,
   O(0) => in23_4,
   O(1) => in23_5,
   O(2) => in23_6,
   O(3) => in23_7
);
HV_reg_0_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in23_8,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_232
);
HV_reg_0_9 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_0_9_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_233
);
HV_reg_1_0 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_1_0_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_192
);
HV_reg_1_10 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_1_10_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_202
);
HV_reg_1_11 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_1_11_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_203
);
HV_reg_1_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in25_12,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_204
);
HV_reg_1_13 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_1_13_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_205
);
HV_reg_1_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in25_14,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_206
);
HV_reg_1_14_i_1 : CARRY4
 port map (
   CI => HV_reg_1_8_i_1_n_0,
   CYINIT => '0',
   DI(0) => b_reg_n_0_12,
   DI(1) => b_reg_n_0_13,
   DI(2) => b_reg_n_0_14,
   DI(3) => b_reg_n_0_15,
   S(0) => HV_1_14_i_5_n_0,
   S(1) => HV_1_14_i_4_n_0,
   S(2) => HV_1_14_i_3_n_0,
   S(3) => HV_1_14_i_2_n_0,
   CO(0) => HV_reg_1_14_i_1_n_3,
   CO(1) => HV_reg_1_14_i_1_n_2,
   CO(2) => HV_reg_1_14_i_1_n_1,
   CO(3) => HV_reg_1_14_i_1_n_0,
   O(0) => in25_12,
   O(1) => in25_13,
   O(2) => in25_14,
   O(3) => in25_15
);
HV_reg_1_15 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_1_15_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_207
);
HV_reg_1_16 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_1_16_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_208
);
HV_reg_1_17 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_1_17_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_209
);
HV_reg_1_18 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_1_18_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_210
);
HV_reg_1_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in25_19,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_211
);
HV_reg_1_19_i_1 : CARRY4
 port map (
   CI => HV_reg_1_14_i_1_n_0,
   CYINIT => '0',
   DI(0) => b_reg_n_0_16,
   DI(1) => b_reg_n_0_17,
   DI(2) => b_reg_n_0_18,
   DI(3) => b_reg_n_0_19,
   S(0) => HV_1_19_i_5_n_0,
   S(1) => HV_1_19_i_4_n_0,
   S(2) => HV_1_19_i_3_n_0,
   S(3) => HV_1_19_i_2_n_0,
   CO(0) => HV_reg_1_19_i_1_n_3,
   CO(1) => HV_reg_1_19_i_1_n_2,
   CO(2) => HV_reg_1_19_i_1_n_1,
   CO(3) => HV_reg_1_19_i_1_n_0,
   O(0) => in25_16,
   O(1) => in25_17,
   O(2) => in25_18,
   O(3) => in25_19
);
HV_reg_1_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in25_1,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_193
);
HV_reg_1_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in25_20,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_212
);
HV_reg_1_21 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_1_21_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_213
);
HV_reg_1_22 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_1_22_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_214
);
HV_reg_1_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in25_23,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_215
);
HV_reg_1_23_i_1 : CARRY4
 port map (
   CI => HV_reg_1_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => b_reg_n_0_20,
   DI(1) => b_reg_n_0_21,
   DI(2) => b_reg_n_0_22,
   DI(3) => b_reg_n_0_23,
   S(0) => HV_1_23_i_5_n_0,
   S(1) => HV_1_23_i_4_n_0,
   S(2) => HV_1_23_i_3_n_0,
   S(3) => HV_1_23_i_2_n_0,
   CO(0) => HV_reg_1_23_i_1_n_3,
   CO(1) => HV_reg_1_23_i_1_n_2,
   CO(2) => HV_reg_1_23_i_1_n_1,
   CO(3) => HV_reg_1_23_i_1_n_0,
   O(0) => in25_20,
   O(1) => in25_21,
   O(2) => in25_22,
   O(3) => in25_23
);
HV_reg_1_24 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_1_24_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_216
);
HV_reg_1_25 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_1_25_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_217
);
HV_reg_1_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in25_26,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_218
);
HV_reg_1_26_i_1 : CARRY4
 port map (
   CI => HV_reg_1_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => b_reg_n_0_24,
   DI(1) => b_reg_n_0_25,
   DI(2) => b_reg_n_0_26,
   DI(3) => b_reg_n_0_27,
   S(0) => HV_1_26_i_5_n_0,
   S(1) => HV_1_26_i_4_n_0,
   S(2) => HV_1_26_i_3_n_0,
   S(3) => HV_1_26_i_2_n_0,
   CO(0) => HV_reg_1_26_i_1_n_3,
   CO(1) => HV_reg_1_26_i_1_n_2,
   CO(2) => HV_reg_1_26_i_1_n_1,
   CO(3) => HV_reg_1_26_i_1_n_0,
   O(0) => in25_24,
   O(1) => in25_25,
   O(2) => in25_26,
   O(3) => in25_27
);
HV_reg_1_27 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_1_27_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_219
);
HV_reg_1_28 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_1_28_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_220
);
HV_reg_1_29 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_1_29_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_221
);
HV_reg_1_2 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_1_2_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_194
);
HV_reg_1_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in25_30,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_222
);
HV_reg_1_30_i_1 : CARRY4
 port map (
   CI => HV_reg_1_26_i_1_n_0,
   CYINIT => '0',
   DI(0) => b_reg_n_0_28,
   DI(1) => b_reg_n_0_29,
   DI(2) => b_reg_n_0_30,
   DI(3) => '0',
   S(0) => HV_1_30_i_5_n_0,
   S(1) => HV_1_30_i_4_n_0,
   S(2) => HV_1_30_i_3_n_0,
   S(3) => HV_1_30_i_2_n_0,
   CO(0) => HV_reg_1_30_i_1_n_3,
   CO(1) => HV_reg_1_30_i_1_n_2,
   CO(2) => HV_reg_1_30_i_1_n_1,
   CO(3) => NLW_HV_reg_1_30_i_1_CO_UNCONNECTED_3,
   O(0) => in25_28,
   O(1) => in25_29,
   O(2) => in25_30,
   O(3) => in25_31
);
HV_reg_1_31 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_1_31_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_223
);
HV_reg_1_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in25_3,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_195
);
HV_reg_1_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => b_reg_n_0_0,
   DI(1) => b_reg_n_0_1,
   DI(2) => b_reg_n_0_2,
   DI(3) => b_reg_n_0_3,
   S(0) => HV_1_3_i_5_n_0,
   S(1) => HV_1_3_i_4_n_0,
   S(2) => HV_1_3_i_3_n_0,
   S(3) => HV_1_3_i_2_n_0,
   CO(0) => HV_reg_1_3_i_1_n_3,
   CO(1) => HV_reg_1_3_i_1_n_2,
   CO(2) => HV_reg_1_3_i_1_n_1,
   CO(3) => HV_reg_1_3_i_1_n_0,
   O(0) => in25_0,
   O(1) => in25_1,
   O(2) => in25_2,
   O(3) => in25_3
);
HV_reg_1_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in25_4,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_196
);
HV_reg_1_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in25_5,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_197
);
HV_reg_1_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in25_6,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_198
);
HV_reg_1_6_i_1 : CARRY4
 port map (
   CI => HV_reg_1_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => b_reg_n_0_4,
   DI(1) => b_reg_n_0_5,
   DI(2) => b_reg_n_0_6,
   DI(3) => b_reg_n_0_7,
   S(0) => HV_1_6_i_5_n_0,
   S(1) => HV_1_6_i_4_n_0,
   S(2) => HV_1_6_i_3_n_0,
   S(3) => HV_1_6_i_2_n_0,
   CO(0) => HV_reg_1_6_i_1_n_3,
   CO(1) => HV_reg_1_6_i_1_n_2,
   CO(2) => HV_reg_1_6_i_1_n_1,
   CO(3) => HV_reg_1_6_i_1_n_0,
   O(0) => in25_4,
   O(1) => in25_5,
   O(2) => in25_6,
   O(3) => in25_7
);
HV_reg_1_7 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_1_7_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_199
);
HV_reg_1_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in25_8,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_200
);
HV_reg_1_8_i_1 : CARRY4
 port map (
   CI => HV_reg_1_6_i_1_n_0,
   CYINIT => '0',
   DI(0) => b_reg_n_0_8,
   DI(1) => b_reg_n_0_9,
   DI(2) => b_reg_n_0_10,
   DI(3) => b_reg_n_0_11,
   S(0) => HV_1_8_i_5_n_0,
   S(1) => HV_1_8_i_4_n_0,
   S(2) => HV_1_8_i_3_n_0,
   S(3) => HV_1_8_i_2_n_0,
   CO(0) => HV_reg_1_8_i_1_n_3,
   CO(1) => HV_reg_1_8_i_1_n_2,
   CO(2) => HV_reg_1_8_i_1_n_1,
   CO(3) => HV_reg_1_8_i_1_n_0,
   O(0) => in25_8,
   O(1) => in25_9,
   O(2) => in25_10,
   O(3) => in25_11
);
HV_reg_1_9 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_1_9_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_201
);
HV_reg_2_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in26_0,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_160
);
HV_reg_2_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in26_10,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_170
);
HV_reg_2_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in26_11,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_171
);
HV_reg_2_11_i_1 : CARRY4
 port map (
   CI => HV_reg_2_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => c_reg_n_0_8,
   DI(1) => c_reg_n_0_9,
   DI(2) => c_reg_n_0_10,
   DI(3) => c_reg_n_0_11,
   S(0) => HV_2_11_i_5_n_0,
   S(1) => HV_2_11_i_4_n_0,
   S(2) => HV_2_11_i_3_n_0,
   S(3) => HV_2_11_i_2_n_0,
   CO(0) => HV_reg_2_11_i_1_n_3,
   CO(1) => HV_reg_2_11_i_1_n_2,
   CO(2) => HV_reg_2_11_i_1_n_1,
   CO(3) => HV_reg_2_11_i_1_n_0,
   O(0) => in26_8,
   O(1) => in26_9,
   O(2) => in26_10,
   O(3) => in26_11
);
HV_reg_2_12 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_2_12_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_172
);
HV_reg_2_13 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_2_13_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_173
);
HV_reg_2_14 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_2_14_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_174
);
HV_reg_2_15 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_2_15_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_175
);
HV_reg_2_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in26_16,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_176
);
HV_reg_2_16_i_1 : CARRY4
 port map (
   CI => HV_reg_2_16_i_2_n_0,
   CYINIT => '0',
   DI(0) => c_reg_n_0_16,
   DI(1) => c_reg_n_0_17,
   DI(2) => c_reg_n_0_18,
   DI(3) => c_reg_n_0_19,
   S(0) => HV_2_16_i_6_n_0,
   S(1) => HV_2_16_i_5_n_0,
   S(2) => HV_2_16_i_4_n_0,
   S(3) => HV_2_16_i_3_n_0,
   CO(0) => HV_reg_2_16_i_1_n_3,
   CO(1) => HV_reg_2_16_i_1_n_2,
   CO(2) => HV_reg_2_16_i_1_n_1,
   CO(3) => HV_reg_2_16_i_1_n_0,
   O(0) => in26_16,
   O(1) => in26_17,
   O(2) => in26_18,
   O(3) => in26_19
);
HV_reg_2_16_i_2 : CARRY4
 port map (
   CI => HV_reg_2_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => c_reg_n_0_12,
   DI(1) => c_reg_n_0_13,
   DI(2) => c_reg_n_0_14,
   DI(3) => c_reg_n_0_15,
   S(0) => HV_2_16_i_10_n_0,
   S(1) => HV_2_16_i_9_n_0,
   S(2) => HV_2_16_i_8_n_0,
   S(3) => HV_2_16_i_7_n_0,
   CO(0) => HV_reg_2_16_i_2_n_3,
   CO(1) => HV_reg_2_16_i_2_n_2,
   CO(2) => HV_reg_2_16_i_2_n_1,
   CO(3) => HV_reg_2_16_i_2_n_0,
   O(0) => in26_12,
   O(1) => in26_13,
   O(2) => in26_14,
   O(3) => in26_15
);
HV_reg_2_17 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_2_17_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_177
);
HV_reg_2_18 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_2_18_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_178
);
HV_reg_2_19 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_2_19_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_179
);
HV_reg_2_1 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_2_1_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_161
);
HV_reg_2_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in26_20,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_180
);
HV_reg_2_21 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_2_21_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_181
);
HV_reg_2_22 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_2_22_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_182
);
HV_reg_2_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in26_23,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_183
);
HV_reg_2_23_i_1 : CARRY4
 port map (
   CI => HV_reg_2_16_i_1_n_0,
   CYINIT => '0',
   DI(0) => c_reg_n_0_20,
   DI(1) => c_reg_n_0_21,
   DI(2) => c_reg_n_0_22,
   DI(3) => c_reg_n_0_23,
   S(0) => HV_2_23_i_5_n_0,
   S(1) => HV_2_23_i_4_n_0,
   S(2) => HV_2_23_i_3_n_0,
   S(3) => HV_2_23_i_2_n_0,
   CO(0) => HV_reg_2_23_i_1_n_3,
   CO(1) => HV_reg_2_23_i_1_n_2,
   CO(2) => HV_reg_2_23_i_1_n_1,
   CO(3) => HV_reg_2_23_i_1_n_0,
   O(0) => in26_20,
   O(1) => in26_21,
   O(2) => in26_22,
   O(3) => in26_23
);
HV_reg_2_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in26_24,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_184
);
HV_reg_2_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in26_25,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_185
);
HV_reg_2_25_i_1 : CARRY4
 port map (
   CI => HV_reg_2_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => c_reg_n_0_24,
   DI(1) => c_reg_n_0_25,
   DI(2) => c_reg_n_0_26,
   DI(3) => c_reg_n_0_27,
   S(0) => HV_2_25_i_5_n_0,
   S(1) => HV_2_25_i_4_n_0,
   S(2) => HV_2_25_i_3_n_0,
   S(3) => HV_2_25_i_2_n_0,
   CO(0) => HV_reg_2_25_i_1_n_3,
   CO(1) => HV_reg_2_25_i_1_n_2,
   CO(2) => HV_reg_2_25_i_1_n_1,
   CO(3) => HV_reg_2_25_i_1_n_0,
   O(0) => in26_24,
   O(1) => in26_25,
   O(2) => in26_26,
   O(3) => in26_27
);
HV_reg_2_26 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_2_26_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_186
);
HV_reg_2_27 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_2_27_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_187
);
HV_reg_2_28 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_2_28_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_188
);
HV_reg_2_29 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_2_29_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_189
);
HV_reg_2_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in26_2,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_162
);
HV_reg_2_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in26_30,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_190
);
HV_reg_2_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in26_31,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_191
);
HV_reg_2_31_i_1 : CARRY4
 port map (
   CI => HV_reg_2_25_i_1_n_0,
   CYINIT => '0',
   DI(0) => c_reg_n_0_28,
   DI(1) => c_reg_n_0_29,
   DI(2) => c_reg_n_0_30,
   DI(3) => '0',
   S(0) => HV_2_31_i_5_n_0,
   S(1) => HV_2_31_i_4_n_0,
   S(2) => HV_2_31_i_3_n_0,
   S(3) => HV_2_31_i_2_n_0,
   CO(0) => HV_reg_2_31_i_1_n_3,
   CO(1) => HV_reg_2_31_i_1_n_2,
   CO(2) => HV_reg_2_31_i_1_n_1,
   CO(3) => NLW_HV_reg_2_31_i_1_CO_UNCONNECTED_3,
   O(0) => in26_28,
   O(1) => in26_29,
   O(2) => in26_30,
   O(3) => in26_31
);
HV_reg_2_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in26_3,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_163
);
HV_reg_2_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => c_reg_n_0_0,
   DI(1) => c_reg_n_0_1,
   DI(2) => c_reg_n_0_2,
   DI(3) => c_reg_n_0_3,
   S(0) => HV_2_3_i_5_n_0,
   S(1) => HV_2_3_i_4_n_0,
   S(2) => HV_2_3_i_3_n_0,
   S(3) => HV_2_3_i_2_n_0,
   CO(0) => HV_reg_2_3_i_1_n_3,
   CO(1) => HV_reg_2_3_i_1_n_2,
   CO(2) => HV_reg_2_3_i_1_n_1,
   CO(3) => HV_reg_2_3_i_1_n_0,
   O(0) => in26_0,
   O(1) => in26_1,
   O(2) => in26_2,
   O(3) => in26_3
);
HV_reg_2_4 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_2_4_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_164
);
HV_reg_2_5 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_2_5_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_165
);
HV_reg_2_6 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_2_6_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_166
);
HV_reg_2_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in26_7,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_167
);
HV_reg_2_7_i_1 : CARRY4
 port map (
   CI => HV_reg_2_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => c_reg_n_0_4,
   DI(1) => c_reg_n_0_5,
   DI(2) => c_reg_n_0_6,
   DI(3) => c_reg_n_0_7,
   S(0) => HV_2_7_i_5_n_0,
   S(1) => HV_2_7_i_4_n_0,
   S(2) => HV_2_7_i_3_n_0,
   S(3) => HV_2_7_i_2_n_0,
   CO(0) => HV_reg_2_7_i_1_n_3,
   CO(1) => HV_reg_2_7_i_1_n_2,
   CO(2) => HV_reg_2_7_i_1_n_1,
   CO(3) => HV_reg_2_7_i_1_n_0,
   O(0) => in26_4,
   O(1) => in26_5,
   O(2) => in26_6,
   O(3) => in26_7
);
HV_reg_2_8 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_2_8_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_168
);
HV_reg_2_9 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_2_9_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_169
);
HV_reg_3_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in27_0,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_128
);
HV_reg_3_10 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_3_10_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_138
);
HV_reg_3_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in27_11,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_139
);
HV_reg_3_11_i_1 : CARRY4
 port map (
   CI => HV_reg_3_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => d_8,
   DI(1) => d_9,
   DI(2) => d_10,
   DI(3) => d_11,
   S(0) => HV_3_11_i_5_n_0,
   S(1) => HV_3_11_i_4_n_0,
   S(2) => HV_3_11_i_3_n_0,
   S(3) => HV_3_11_i_2_n_0,
   CO(0) => HV_reg_3_11_i_1_n_3,
   CO(1) => HV_reg_3_11_i_1_n_2,
   CO(2) => HV_reg_3_11_i_1_n_1,
   CO(3) => HV_reg_3_11_i_1_n_0,
   O(0) => in27_8,
   O(1) => in27_9,
   O(2) => in27_10,
   O(3) => in27_11
);
HV_reg_3_12 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_3_12_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_140
);
HV_reg_3_13 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_3_13_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_141
);
HV_reg_3_14 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_3_14_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_142
);
HV_reg_3_15 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_3_15_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_143
);
HV_reg_3_15_i_2 : CARRY4
 port map (
   CI => HV_reg_3_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => d_12,
   DI(1) => d_13,
   DI(2) => d_14,
   DI(3) => d_15,
   S(0) => HV_3_15_i_6_n_0,
   S(1) => HV_3_15_i_5_n_0,
   S(2) => HV_3_15_i_4_n_0,
   S(3) => HV_3_15_i_3_n_0,
   CO(0) => HV_reg_3_15_i_2_n_3,
   CO(1) => HV_reg_3_15_i_2_n_2,
   CO(2) => HV_reg_3_15_i_2_n_1,
   CO(3) => HV_reg_3_15_i_2_n_0,
   O(0) => in27_12,
   O(1) => in27_13,
   O(2) => in27_14,
   O(3) => in27_15
);
HV_reg_3_16 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_3_16_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_144
);
HV_reg_3_17 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_3_17_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_145
);
HV_reg_3_18 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_3_18_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_146
);
HV_reg_3_19 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_3_19_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_147
);
HV_reg_3_1 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_3_1_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_129
);
HV_reg_3_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in27_20,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_148
);
HV_reg_3_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in27_21,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_149
);
HV_reg_3_22 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_3_22_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_150
);
HV_reg_3_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in27_23,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_151
);
HV_reg_3_23_i_1 : CARRY4
 port map (
   CI => HV_reg_3_23_i_2_n_0,
   CYINIT => '0',
   DI(0) => d_20,
   DI(1) => d_21,
   DI(2) => d_22,
   DI(3) => d_23,
   S(0) => HV_3_23_i_6_n_0,
   S(1) => HV_3_23_i_5_n_0,
   S(2) => HV_3_23_i_4_n_0,
   S(3) => HV_3_23_i_3_n_0,
   CO(0) => HV_reg_3_23_i_1_n_3,
   CO(1) => HV_reg_3_23_i_1_n_2,
   CO(2) => HV_reg_3_23_i_1_n_1,
   CO(3) => HV_reg_3_23_i_1_n_0,
   O(0) => in27_20,
   O(1) => in27_21,
   O(2) => in27_22,
   O(3) => in27_23
);
HV_reg_3_23_i_2 : CARRY4
 port map (
   CI => HV_reg_3_15_i_2_n_0,
   CYINIT => '0',
   DI(0) => d_16,
   DI(1) => d_17,
   DI(2) => d_18,
   DI(3) => d_19,
   S(0) => HV_3_23_i_10_n_0,
   S(1) => HV_3_23_i_9_n_0,
   S(2) => HV_3_23_i_8_n_0,
   S(3) => HV_3_23_i_7_n_0,
   CO(0) => HV_reg_3_23_i_2_n_3,
   CO(1) => HV_reg_3_23_i_2_n_2,
   CO(2) => HV_reg_3_23_i_2_n_1,
   CO(3) => HV_reg_3_23_i_2_n_0,
   O(0) => in27_16,
   O(1) => in27_17,
   O(2) => in27_18,
   O(3) => in27_19
);
HV_reg_3_24 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_3_24_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_152
);
HV_reg_3_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in27_25,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_153
);
HV_reg_3_26 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_3_26_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_154
);
HV_reg_3_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in27_27,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_155
);
HV_reg_3_27_i_1 : CARRY4
 port map (
   CI => HV_reg_3_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => d_24,
   DI(1) => d_25,
   DI(2) => d_26,
   DI(3) => d_27,
   S(0) => HV_3_27_i_5_n_0,
   S(1) => HV_3_27_i_4_n_0,
   S(2) => HV_3_27_i_3_n_0,
   S(3) => HV_3_27_i_2_n_0,
   CO(0) => HV_reg_3_27_i_1_n_3,
   CO(1) => HV_reg_3_27_i_1_n_2,
   CO(2) => HV_reg_3_27_i_1_n_1,
   CO(3) => HV_reg_3_27_i_1_n_0,
   O(0) => in27_24,
   O(1) => in27_25,
   O(2) => in27_26,
   O(3) => in27_27
);
HV_reg_3_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in27_28,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_156
);
HV_reg_3_29 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_3_29_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_157
);
HV_reg_3_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in27_2,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_130
);
HV_reg_3_2_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => d_0,
   DI(1) => d_1,
   DI(2) => d_2,
   DI(3) => d_3,
   S(0) => HV_3_2_i_5_n_0,
   S(1) => HV_3_2_i_4_n_0,
   S(2) => HV_3_2_i_3_n_0,
   S(3) => HV_3_2_i_2_n_0,
   CO(0) => HV_reg_3_2_i_1_n_3,
   CO(1) => HV_reg_3_2_i_1_n_2,
   CO(2) => HV_reg_3_2_i_1_n_1,
   CO(3) => HV_reg_3_2_i_1_n_0,
   O(0) => in27_0,
   O(1) => in27_1,
   O(2) => in27_2,
   O(3) => in27_3
);
HV_reg_3_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in27_30,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_158
);
HV_reg_3_30_i_1 : CARRY4
 port map (
   CI => HV_reg_3_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => d_28,
   DI(1) => d_29,
   DI(2) => d_30,
   DI(3) => '0',
   S(0) => HV_3_30_i_5_n_0,
   S(1) => HV_3_30_i_4_n_0,
   S(2) => HV_3_30_i_3_n_0,
   S(3) => HV_3_30_i_2_n_0,
   CO(0) => HV_reg_3_30_i_1_n_3,
   CO(1) => HV_reg_3_30_i_1_n_2,
   CO(2) => HV_reg_3_30_i_1_n_1,
   CO(3) => NLW_HV_reg_3_30_i_1_CO_UNCONNECTED_3,
   O(0) => in27_28,
   O(1) => in27_29,
   O(2) => in27_30,
   O(3) => in27_31
);
HV_reg_3_31 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_3_31_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_159
);
HV_reg_3_3 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_3_3_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_131
);
HV_reg_3_4 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_3_4_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_132
);
HV_reg_3_5 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_3_5_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_133
);
HV_reg_3_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in27_6,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_134
);
HV_reg_3_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in27_7,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_135
);
HV_reg_3_7_i_1 : CARRY4
 port map (
   CI => HV_reg_3_2_i_1_n_0,
   CYINIT => '0',
   DI(0) => d_4,
   DI(1) => d_5,
   DI(2) => d_6,
   DI(3) => d_7,
   S(0) => HV_3_7_i_5_n_0,
   S(1) => HV_3_7_i_4_n_0,
   S(2) => HV_3_7_i_3_n_0,
   S(3) => HV_3_7_i_2_n_0,
   CO(0) => HV_reg_3_7_i_1_n_3,
   CO(1) => HV_reg_3_7_i_1_n_2,
   CO(2) => HV_reg_3_7_i_1_n_1,
   CO(3) => HV_reg_3_7_i_1_n_0,
   O(0) => in27_4,
   O(1) => in27_5,
   O(2) => in27_6,
   O(3) => in27_7
);
HV_reg_3_8 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_3_8_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_136
);
HV_reg_3_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in27_9,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_137
);
HV_reg_4_0 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_4_0_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_96
);
HV_reg_4_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in28_10,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_106
);
HV_reg_4_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in28_11,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_107
);
HV_reg_4_11_i_1 : CARRY4
 port map (
   CI => HV_reg_4_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => ROTR11_out_3,
   DI(1) => ROTR11_out_2,
   DI(2) => ROTR11_out_1,
   DI(3) => ROTR11_out_32,
   S(0) => HV_4_11_i_5_n_0,
   S(1) => HV_4_11_i_4_n_0,
   S(2) => HV_4_11_i_3_n_0,
   S(3) => HV_4_11_i_2_n_0,
   CO(0) => HV_reg_4_11_i_1_n_3,
   CO(1) => HV_reg_4_11_i_1_n_2,
   CO(2) => HV_reg_4_11_i_1_n_1,
   CO(3) => HV_reg_4_11_i_1_n_0,
   O(0) => in28_8,
   O(1) => in28_9,
   O(2) => in28_10,
   O(3) => in28_11
);
HV_reg_4_12 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_4_12_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_108
);
HV_reg_4_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in28_13,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_109
);
HV_reg_4_14 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_4_14_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_110
);
HV_reg_4_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in28_15,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_111
);
HV_reg_4_15_i_1 : CARRY4
 port map (
   CI => HV_reg_4_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => ROTR11_out_31,
   DI(1) => ROTR11_out_30,
   DI(2) => ROTR11_out_29,
   DI(3) => ROTR11_out_28,
   S(0) => HV_4_15_i_5_n_0,
   S(1) => HV_4_15_i_4_n_0,
   S(2) => HV_4_15_i_3_n_0,
   S(3) => HV_4_15_i_2_n_0,
   CO(0) => HV_reg_4_15_i_1_n_3,
   CO(1) => HV_reg_4_15_i_1_n_2,
   CO(2) => HV_reg_4_15_i_1_n_1,
   CO(3) => HV_reg_4_15_i_1_n_0,
   O(0) => in28_12,
   O(1) => in28_13,
   O(2) => in28_14,
   O(3) => in28_15
);
HV_reg_4_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in28_16,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_112
);
HV_reg_4_16_i_1 : CARRY4
 port map (
   CI => HV_reg_4_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => ROTR11_out_27,
   DI(1) => ROTR11_out_26,
   DI(2) => ROTR11_out_25,
   DI(3) => ROTR11_out_24,
   S(0) => HV_4_16_i_5_n_0,
   S(1) => HV_4_16_i_4_n_0,
   S(2) => HV_4_16_i_3_n_0,
   S(3) => HV_4_16_i_2_n_0,
   CO(0) => HV_reg_4_16_i_1_n_3,
   CO(1) => HV_reg_4_16_i_1_n_2,
   CO(2) => HV_reg_4_16_i_1_n_1,
   CO(3) => HV_reg_4_16_i_1_n_0,
   O(0) => in28_16,
   O(1) => in28_17,
   O(2) => in28_18,
   O(3) => in28_19
);
HV_reg_4_17 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_4_17_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_113
);
HV_reg_4_18 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_4_18_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_114
);
HV_reg_4_19 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_4_19_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_115
);
HV_reg_4_1 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_4_1_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_97
);
HV_reg_4_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in28_20,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_116
);
HV_reg_4_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in28_21,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_117
);
HV_reg_4_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in28_22,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_118
);
HV_reg_4_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in28_23,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_119
);
HV_reg_4_23_i_1 : CARRY4
 port map (
   CI => HV_reg_4_16_i_1_n_0,
   CYINIT => '0',
   DI(0) => ROTR11_out_23,
   DI(1) => ROTR11_out_22,
   DI(2) => ROTR11_out_21,
   DI(3) => ROTR11_out_20,
   S(0) => HV_4_23_i_5_n_0,
   S(1) => HV_4_23_i_4_n_0,
   S(2) => HV_4_23_i_3_n_0,
   S(3) => HV_4_23_i_2_n_0,
   CO(0) => HV_reg_4_23_i_1_n_3,
   CO(1) => HV_reg_4_23_i_1_n_2,
   CO(2) => HV_reg_4_23_i_1_n_1,
   CO(3) => HV_reg_4_23_i_1_n_0,
   O(0) => in28_20,
   O(1) => in28_21,
   O(2) => in28_22,
   O(3) => in28_23
);
HV_reg_4_24 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_4_24_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_120
);
HV_reg_4_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in28_25,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_121
);
HV_reg_4_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in28_26,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_122
);
HV_reg_4_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in28_27,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_123
);
HV_reg_4_27_i_1 : CARRY4
 port map (
   CI => HV_reg_4_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => ROTR11_out_19,
   DI(1) => ROTR11_out_18,
   DI(2) => ROTR11_out_17,
   DI(3) => ROTR11_out_16,
   S(0) => HV_4_27_i_5_n_0,
   S(1) => HV_4_27_i_4_n_0,
   S(2) => HV_4_27_i_3_n_0,
   S(3) => HV_4_27_i_2_n_0,
   CO(0) => HV_reg_4_27_i_1_n_3,
   CO(1) => HV_reg_4_27_i_1_n_2,
   CO(2) => HV_reg_4_27_i_1_n_1,
   CO(3) => HV_reg_4_27_i_1_n_0,
   O(0) => in28_24,
   O(1) => in28_25,
   O(2) => in28_26,
   O(3) => in28_27
);
HV_reg_4_28 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_4_28_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_124
);
HV_reg_4_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in28_29,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_125
);
HV_reg_4_2 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_4_2_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_98
);
HV_reg_4_30 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_4_30_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_126
);
HV_reg_4_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in28_31,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_127
);
HV_reg_4_31_i_1 : CARRY4
 port map (
   CI => HV_reg_4_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => ROTR11_out_15,
   DI(1) => ROTR11_out_14,
   DI(2) => ROTR11_out_13,
   DI(3) => '0',
   S(0) => HV_4_31_i_5_n_0,
   S(1) => HV_4_31_i_4_n_0,
   S(2) => HV_4_31_i_3_n_0,
   S(3) => HV_4_31_i_2_n_0,
   CO(0) => HV_reg_4_31_i_1_n_3,
   CO(1) => HV_reg_4_31_i_1_n_2,
   CO(2) => HV_reg_4_31_i_1_n_1,
   CO(3) => NLW_HV_reg_4_31_i_1_CO_UNCONNECTED_3,
   O(0) => in28_28,
   O(1) => in28_29,
   O(2) => in28_30,
   O(3) => in28_31
);
HV_reg_4_3 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_4_3_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_99
);
HV_reg_4_4 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_4_4_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_100
);
HV_reg_4_5 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_4_5_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_101
);
HV_reg_4_6 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_4_6_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_102
);
HV_reg_4_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in28_7,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_103
);
HV_reg_4_7_i_1 : CARRY4
 port map (
   CI => HV_reg_4_7_i_2_n_0,
   CYINIT => '0',
   DI(0) => ROTR11_out_7,
   DI(1) => ROTR11_out_6,
   DI(2) => ROTR11_out_5,
   DI(3) => ROTR11_out_4,
   S(0) => HV_4_7_i_6_n_0,
   S(1) => HV_4_7_i_5_n_0,
   S(2) => HV_4_7_i_4_n_0,
   S(3) => HV_4_7_i_3_n_0,
   CO(0) => HV_reg_4_7_i_1_n_3,
   CO(1) => HV_reg_4_7_i_1_n_2,
   CO(2) => HV_reg_4_7_i_1_n_1,
   CO(3) => HV_reg_4_7_i_1_n_0,
   O(0) => in28_4,
   O(1) => in28_5,
   O(2) => in28_6,
   O(3) => in28_7
);
HV_reg_4_7_i_2 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => ROTR11_out_11,
   DI(1) => ROTR11_out_10,
   DI(2) => ROTR11_out_9,
   DI(3) => ROTR11_out_8,
   S(0) => HV_4_7_i_10_n_0,
   S(1) => HV_4_7_i_9_n_0,
   S(2) => HV_4_7_i_8_n_0,
   S(3) => HV_4_7_i_7_n_0,
   CO(0) => HV_reg_4_7_i_2_n_3,
   CO(1) => HV_reg_4_7_i_2_n_2,
   CO(2) => HV_reg_4_7_i_2_n_1,
   CO(3) => HV_reg_4_7_i_2_n_0,
   O(0) => in28_0,
   O(1) => in28_1,
   O(2) => in28_2,
   O(3) => in28_3
);
HV_reg_4_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in28_8,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_104
);
HV_reg_4_9 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_4_9_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_105
);
HV_reg_5_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in29_0,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_64
);
HV_reg_5_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in29_10,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_74
);
HV_reg_5_10_i_1 : CARRY4
 port map (
   CI => HV_reg_5_6_i_1_n_0,
   CYINIT => '0',
   DI(0) => f_reg_n_0_8,
   DI(1) => f_reg_n_0_9,
   DI(2) => f_reg_n_0_10,
   DI(3) => f_reg_n_0_11,
   S(0) => HV_5_10_i_5_n_0,
   S(1) => HV_5_10_i_4_n_0,
   S(2) => HV_5_10_i_3_n_0,
   S(3) => HV_5_10_i_2_n_0,
   CO(0) => HV_reg_5_10_i_1_n_3,
   CO(1) => HV_reg_5_10_i_1_n_2,
   CO(2) => HV_reg_5_10_i_1_n_1,
   CO(3) => HV_reg_5_10_i_1_n_0,
   O(0) => in29_8,
   O(1) => in29_9,
   O(2) => in29_10,
   O(3) => in29_11
);
HV_reg_5_11 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_5_11_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_75
);
HV_reg_5_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in29_12,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_76
);
HV_reg_5_13 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_5_13_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_77
);
HV_reg_5_14 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_5_14_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_78
);
HV_reg_5_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in29_15,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_79
);
HV_reg_5_15_i_1 : CARRY4
 port map (
   CI => HV_reg_5_10_i_1_n_0,
   CYINIT => '0',
   DI(0) => f_reg_n_0_12,
   DI(1) => f_reg_n_0_13,
   DI(2) => f_reg_n_0_14,
   DI(3) => f_reg_n_0_15,
   S(0) => HV_5_15_i_5_n_0,
   S(1) => HV_5_15_i_4_n_0,
   S(2) => HV_5_15_i_3_n_0,
   S(3) => HV_5_15_i_2_n_0,
   CO(0) => HV_reg_5_15_i_1_n_3,
   CO(1) => HV_reg_5_15_i_1_n_2,
   CO(2) => HV_reg_5_15_i_1_n_1,
   CO(3) => HV_reg_5_15_i_1_n_0,
   O(0) => in29_12,
   O(1) => in29_13,
   O(2) => in29_14,
   O(3) => in29_15
);
HV_reg_5_16 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_5_16_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_80
);
HV_reg_5_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in29_17,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_81
);
HV_reg_5_18 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_5_18_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_82
);
HV_reg_5_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in29_19,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_83
);
HV_reg_5_19_i_1 : CARRY4
 port map (
   CI => HV_reg_5_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => f_reg_n_0_16,
   DI(1) => f_reg_n_0_17,
   DI(2) => f_reg_n_0_18,
   DI(3) => f_reg_n_0_19,
   S(0) => HV_5_19_i_5_n_0,
   S(1) => HV_5_19_i_4_n_0,
   S(2) => HV_5_19_i_3_n_0,
   S(3) => HV_5_19_i_2_n_0,
   CO(0) => HV_reg_5_19_i_1_n_3,
   CO(1) => HV_reg_5_19_i_1_n_2,
   CO(2) => HV_reg_5_19_i_1_n_1,
   CO(3) => HV_reg_5_19_i_1_n_0,
   O(0) => in29_16,
   O(1) => in29_17,
   O(2) => in29_18,
   O(3) => in29_19
);
HV_reg_5_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in29_1,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_65
);
HV_reg_5_1_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => f_reg_n_0_0,
   DI(1) => f_reg_n_0_1,
   DI(2) => f_reg_n_0_2,
   DI(3) => f_reg_n_0_3,
   S(0) => HV_5_1_i_5_n_0,
   S(1) => HV_5_1_i_4_n_0,
   S(2) => HV_5_1_i_3_n_0,
   S(3) => HV_5_1_i_2_n_0,
   CO(0) => HV_reg_5_1_i_1_n_3,
   CO(1) => HV_reg_5_1_i_1_n_2,
   CO(2) => HV_reg_5_1_i_1_n_1,
   CO(3) => HV_reg_5_1_i_1_n_0,
   O(0) => in29_0,
   O(1) => in29_1,
   O(2) => in29_2,
   O(3) => in29_3
);
HV_reg_5_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in29_20,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_84
);
HV_reg_5_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in29_21,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_85
);
HV_reg_5_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in29_22,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_86
);
HV_reg_5_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in29_23,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_87
);
HV_reg_5_23_i_1 : CARRY4
 port map (
   CI => HV_reg_5_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => f_reg_n_0_20,
   DI(1) => f_reg_n_0_21,
   DI(2) => f_reg_n_0_22,
   DI(3) => f_reg_n_0_23,
   S(0) => HV_5_23_i_5_n_0,
   S(1) => HV_5_23_i_4_n_0,
   S(2) => HV_5_23_i_3_n_0,
   S(3) => HV_5_23_i_2_n_0,
   CO(0) => HV_reg_5_23_i_1_n_3,
   CO(1) => HV_reg_5_23_i_1_n_2,
   CO(2) => HV_reg_5_23_i_1_n_1,
   CO(3) => HV_reg_5_23_i_1_n_0,
   O(0) => in29_20,
   O(1) => in29_21,
   O(2) => in29_22,
   O(3) => in29_23
);
HV_reg_5_24 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_5_24_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_88
);
HV_reg_5_25 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_5_25_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_89
);
HV_reg_5_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in29_26,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_90
);
HV_reg_5_26_i_1 : CARRY4
 port map (
   CI => HV_reg_5_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => f_reg_n_0_24,
   DI(1) => f_reg_n_0_25,
   DI(2) => f_reg_n_0_26,
   DI(3) => f_reg_n_0_27,
   S(0) => HV_5_26_i_5_n_0,
   S(1) => HV_5_26_i_4_n_0,
   S(2) => HV_5_26_i_3_n_0,
   S(3) => HV_5_26_i_2_n_0,
   CO(0) => HV_reg_5_26_i_1_n_3,
   CO(1) => HV_reg_5_26_i_1_n_2,
   CO(2) => HV_reg_5_26_i_1_n_1,
   CO(3) => HV_reg_5_26_i_1_n_0,
   O(0) => in29_24,
   O(1) => in29_25,
   O(2) => in29_26,
   O(3) => in29_27
);
HV_reg_5_27 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_5_27_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_91
);
HV_reg_5_28 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_5_28_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_92
);
HV_reg_5_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in29_29,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_93
);
HV_reg_5_2 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_5_2_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_66
);
HV_reg_5_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in29_30,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_94
);
HV_reg_5_30_i_1 : CARRY4
 port map (
   CI => HV_reg_5_26_i_1_n_0,
   CYINIT => '0',
   DI(0) => f_reg_n_0_28,
   DI(1) => f_reg_n_0_29,
   DI(2) => f_reg_n_0_30,
   DI(3) => '0',
   S(0) => HV_5_30_i_5_n_0,
   S(1) => HV_5_30_i_4_n_0,
   S(2) => HV_5_30_i_3_n_0,
   S(3) => HV_5_30_i_2_n_0,
   CO(0) => HV_reg_5_30_i_1_n_3,
   CO(1) => HV_reg_5_30_i_1_n_2,
   CO(2) => HV_reg_5_30_i_1_n_1,
   CO(3) => NLW_HV_reg_5_30_i_1_CO_UNCONNECTED_3,
   O(0) => in29_28,
   O(1) => in29_29,
   O(2) => in29_30,
   O(3) => in29_31
);
HV_reg_5_31 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_5_31_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_95
);
HV_reg_5_3 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_5_3_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_67
);
HV_reg_5_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in29_4,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_68
);
HV_reg_5_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in29_5,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_69
);
HV_reg_5_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in29_6,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_70
);
HV_reg_5_6_i_1 : CARRY4
 port map (
   CI => HV_reg_5_1_i_1_n_0,
   CYINIT => '0',
   DI(0) => f_reg_n_0_4,
   DI(1) => f_reg_n_0_5,
   DI(2) => f_reg_n_0_6,
   DI(3) => f_reg_n_0_7,
   S(0) => HV_5_6_i_5_n_0,
   S(1) => HV_5_6_i_4_n_0,
   S(2) => HV_5_6_i_3_n_0,
   S(3) => HV_5_6_i_2_n_0,
   CO(0) => HV_reg_5_6_i_1_n_3,
   CO(1) => HV_reg_5_6_i_1_n_2,
   CO(2) => HV_reg_5_6_i_1_n_1,
   CO(3) => HV_reg_5_6_i_1_n_0,
   O(0) => in29_4,
   O(1) => in29_5,
   O(2) => in29_6,
   O(3) => in29_7
);
HV_reg_5_7 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_5_7_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_71
);
HV_reg_5_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in29_8,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_72
);
HV_reg_5_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in29_9,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_73
);
HV_reg_6_0 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_6_0_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_32
);
HV_reg_6_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in30_10,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_42
);
HV_reg_6_10_i_1 : CARRY4
 port map (
   CI => HV_reg_6_6_i_1_n_0,
   CYINIT => '0',
   DI(0) => g_reg_n_0_8,
   DI(1) => g_reg_n_0_9,
   DI(2) => g_reg_n_0_10,
   DI(3) => g_reg_n_0_11,
   S(0) => HV_6_10_i_5_n_0,
   S(1) => HV_6_10_i_4_n_0,
   S(2) => HV_6_10_i_3_n_0,
   S(3) => HV_6_10_i_2_n_0,
   CO(0) => HV_reg_6_10_i_1_n_3,
   CO(1) => HV_reg_6_10_i_1_n_2,
   CO(2) => HV_reg_6_10_i_1_n_1,
   CO(3) => HV_reg_6_10_i_1_n_0,
   O(0) => in30_8,
   O(1) => in30_9,
   O(2) => in30_10,
   O(3) => in30_11
);
HV_reg_6_11 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_6_11_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_43
);
HV_reg_6_12 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_6_12_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_44
);
HV_reg_6_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in30_13,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_45
);
HV_reg_6_13_i_1 : CARRY4
 port map (
   CI => HV_reg_6_10_i_1_n_0,
   CYINIT => '0',
   DI(0) => g_reg_n_0_12,
   DI(1) => g_reg_n_0_13,
   DI(2) => g_reg_n_0_14,
   DI(3) => g_reg_n_0_15,
   S(0) => HV_6_13_i_5_n_0,
   S(1) => HV_6_13_i_4_n_0,
   S(2) => HV_6_13_i_3_n_0,
   S(3) => HV_6_13_i_2_n_0,
   CO(0) => HV_reg_6_13_i_1_n_3,
   CO(1) => HV_reg_6_13_i_1_n_2,
   CO(2) => HV_reg_6_13_i_1_n_1,
   CO(3) => HV_reg_6_13_i_1_n_0,
   O(0) => in30_12,
   O(1) => in30_13,
   O(2) => in30_14,
   O(3) => in30_15
);
HV_reg_6_14 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_6_14_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_46
);
HV_reg_6_15 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_6_15_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_47
);
HV_reg_6_16 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_6_16_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_48
);
HV_reg_6_17 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_6_17_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_49
);
HV_reg_6_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in30_18,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_50
);
HV_reg_6_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in30_19,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_51
);
HV_reg_6_19_i_1 : CARRY4
 port map (
   CI => HV_reg_6_13_i_1_n_0,
   CYINIT => '0',
   DI(0) => g_reg_n_0_16,
   DI(1) => g_reg_n_0_17,
   DI(2) => g_reg_n_0_18,
   DI(3) => g_reg_n_0_19,
   S(0) => HV_6_19_i_5_n_0,
   S(1) => HV_6_19_i_4_n_0,
   S(2) => HV_6_19_i_3_n_0,
   S(3) => HV_6_19_i_2_n_0,
   CO(0) => HV_reg_6_19_i_1_n_3,
   CO(1) => HV_reg_6_19_i_1_n_2,
   CO(2) => HV_reg_6_19_i_1_n_1,
   CO(3) => HV_reg_6_19_i_1_n_0,
   O(0) => in30_16,
   O(1) => in30_17,
   O(2) => in30_18,
   O(3) => in30_19
);
HV_reg_6_1 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_6_1_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_33
);
HV_reg_6_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in30_20,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_52
);
HV_reg_6_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in30_21,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_53
);
HV_reg_6_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in30_22,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_54
);
HV_reg_6_22_i_1 : CARRY4
 port map (
   CI => HV_reg_6_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => g_reg_n_0_20,
   DI(1) => g_reg_n_0_21,
   DI(2) => g_reg_n_0_22,
   DI(3) => g_reg_n_0_23,
   S(0) => HV_6_22_i_5_n_0,
   S(1) => HV_6_22_i_4_n_0,
   S(2) => HV_6_22_i_3_n_0,
   S(3) => HV_6_22_i_2_n_0,
   CO(0) => HV_reg_6_22_i_1_n_3,
   CO(1) => HV_reg_6_22_i_1_n_2,
   CO(2) => HV_reg_6_22_i_1_n_1,
   CO(3) => HV_reg_6_22_i_1_n_0,
   O(0) => in30_20,
   O(1) => in30_21,
   O(2) => in30_22,
   O(3) => in30_23
);
HV_reg_6_23 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_6_23_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_55
);
HV_reg_6_24 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_6_24_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_56
);
HV_reg_6_25 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_6_25_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_57
);
HV_reg_6_26 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_6_26_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_58
);
HV_reg_6_27 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_6_27_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_59
);
HV_reg_6_28 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_6_28_i_2_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_60
);
HV_reg_6_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in30_29,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_61
);
HV_reg_6_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in30_2,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_34
);
HV_reg_6_2_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => g_reg_n_0_0,
   DI(1) => g_reg_n_0_1,
   DI(2) => g_reg_n_0_2,
   DI(3) => g_reg_n_0_3,
   S(0) => HV_6_2_i_5_n_0,
   S(1) => HV_6_2_i_4_n_0,
   S(2) => HV_6_2_i_3_n_0,
   S(3) => HV_6_2_i_2_n_0,
   CO(0) => HV_reg_6_2_i_1_n_3,
   CO(1) => HV_reg_6_2_i_1_n_2,
   CO(2) => HV_reg_6_2_i_1_n_1,
   CO(3) => HV_reg_6_2_i_1_n_0,
   O(0) => in30_0,
   O(1) => in30_1,
   O(2) => in30_2,
   O(3) => in30_3
);
HV_reg_6_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in30_30,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_62
);
HV_reg_6_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in30_31,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_63
);
HV_reg_6_31_i_3 : CARRY4
 port map (
   CI => HV_reg_6_31_i_4_n_0,
   CYINIT => '0',
   DI(0) => g_reg_n_0_28,
   DI(1) => g_reg_n_0_29,
   DI(2) => g_reg_n_0_30,
   DI(3) => '0',
   S(0) => HV_6_31_i_8_n_0,
   S(1) => HV_6_31_i_7_n_0,
   S(2) => HV_6_31_i_6_n_0,
   S(3) => HV_6_31_i_5_n_0,
   CO(0) => HV_reg_6_31_i_3_n_3,
   CO(1) => HV_reg_6_31_i_3_n_2,
   CO(2) => HV_reg_6_31_i_3_n_1,
   CO(3) => NLW_HV_reg_6_31_i_3_CO_UNCONNECTED_3,
   O(0) => in30_28,
   O(1) => in30_29,
   O(2) => in30_30,
   O(3) => in30_31
);
HV_reg_6_31_i_4 : CARRY4
 port map (
   CI => HV_reg_6_22_i_1_n_0,
   CYINIT => '0',
   DI(0) => g_reg_n_0_24,
   DI(1) => g_reg_n_0_25,
   DI(2) => g_reg_n_0_26,
   DI(3) => g_reg_n_0_27,
   S(0) => HV_6_31_i_12_n_0,
   S(1) => HV_6_31_i_11_n_0,
   S(2) => HV_6_31_i_10_n_0,
   S(3) => HV_6_31_i_9_n_0,
   CO(0) => HV_reg_6_31_i_4_n_3,
   CO(1) => HV_reg_6_31_i_4_n_2,
   CO(2) => HV_reg_6_31_i_4_n_1,
   CO(3) => HV_reg_6_31_i_4_n_0,
   O(0) => in30_24,
   O(1) => in30_25,
   O(2) => in30_26,
   O(3) => in30_27
);
HV_reg_6_3 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_6_3_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_35
);
HV_reg_6_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in30_4,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_36
);
HV_reg_6_5 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_6_5_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_37
);
HV_reg_6_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in30_6,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_38
);
HV_reg_6_6_i_1 : CARRY4
 port map (
   CI => HV_reg_6_2_i_1_n_0,
   CYINIT => '0',
   DI(0) => g_reg_n_0_4,
   DI(1) => g_reg_n_0_5,
   DI(2) => g_reg_n_0_6,
   DI(3) => g_reg_n_0_7,
   S(0) => HV_6_6_i_5_n_0,
   S(1) => HV_6_6_i_4_n_0,
   S(2) => HV_6_6_i_3_n_0,
   S(3) => HV_6_6_i_2_n_0,
   CO(0) => HV_reg_6_6_i_1_n_3,
   CO(1) => HV_reg_6_6_i_1_n_2,
   CO(2) => HV_reg_6_6_i_1_n_1,
   CO(3) => HV_reg_6_6_i_1_n_0,
   O(0) => in30_4,
   O(1) => in30_5,
   O(2) => in30_6,
   O(3) => in30_7
);
HV_reg_6_7 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_6_7_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_39
);
HV_reg_6_8 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_6_8_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_40
);
HV_reg_6_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in30_9,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_41
);
HV_reg_7_0 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_7_0_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_0
);
HV_reg_7_10 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_7_10_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_10
);
HV_reg_7_11 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_7_11_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_11
);
HV_reg_7_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in31_12,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_12
);
HV_reg_7_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in31_13,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_13
);
HV_reg_7_13_i_1 : CARRY4
 port map (
   CI => HV_reg_7_9_i_1_n_0,
   CYINIT => '0',
   DI(0) => h_12,
   DI(1) => h_13,
   DI(2) => h_14,
   DI(3) => h_15,
   S(0) => HV_7_13_i_5_n_0,
   S(1) => HV_7_13_i_4_n_0,
   S(2) => HV_7_13_i_3_n_0,
   S(3) => HV_7_13_i_2_n_0,
   CO(0) => HV_reg_7_13_i_1_n_3,
   CO(1) => HV_reg_7_13_i_1_n_2,
   CO(2) => HV_reg_7_13_i_1_n_1,
   CO(3) => HV_reg_7_13_i_1_n_0,
   O(0) => in31_12,
   O(1) => in31_13,
   O(2) => in31_14,
   O(3) => in31_15
);
HV_reg_7_14 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_7_14_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_14
);
HV_reg_7_15 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_7_15_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_15
);
HV_reg_7_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in31_16,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_16
);
HV_reg_7_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in31_17,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_17
);
HV_reg_7_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in31_18,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_18
);
HV_reg_7_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in31_19,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_19
);
HV_reg_7_19_i_1 : CARRY4
 port map (
   CI => HV_reg_7_13_i_1_n_0,
   CYINIT => '0',
   DI(0) => h_16,
   DI(1) => h_17,
   DI(2) => h_18,
   DI(3) => h_19,
   S(0) => HV_7_19_i_5_n_0,
   S(1) => HV_7_19_i_4_n_0,
   S(2) => HV_7_19_i_3_n_0,
   S(3) => HV_7_19_i_2_n_0,
   CO(0) => HV_reg_7_19_i_1_n_3,
   CO(1) => HV_reg_7_19_i_1_n_2,
   CO(2) => HV_reg_7_19_i_1_n_1,
   CO(3) => HV_reg_7_19_i_1_n_0,
   O(0) => in31_16,
   O(1) => in31_17,
   O(2) => in31_18,
   O(3) => in31_19
);
HV_reg_7_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in31_1,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_1
);
HV_reg_7_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in31_20,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_20
);
HV_reg_7_20_i_1 : CARRY4
 port map (
   CI => HV_reg_7_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => h_20,
   DI(1) => h_21,
   DI(2) => h_22,
   DI(3) => h_23,
   S(0) => HV_7_20_i_5_n_0,
   S(1) => HV_7_20_i_4_n_0,
   S(2) => HV_7_20_i_3_n_0,
   S(3) => HV_7_20_i_2_n_0,
   CO(0) => HV_reg_7_20_i_1_n_3,
   CO(1) => HV_reg_7_20_i_1_n_2,
   CO(2) => HV_reg_7_20_i_1_n_1,
   CO(3) => HV_reg_7_20_i_1_n_0,
   O(0) => in31_20,
   O(1) => in31_21,
   O(2) => in31_22,
   O(3) => in31_23
);
HV_reg_7_21 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_7_21_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_21
);
HV_reg_7_22 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_7_22_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_22
);
HV_reg_7_23 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_7_23_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_23
);
HV_reg_7_24 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_7_24_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_24
);
HV_reg_7_25 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_7_25_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_25
);
HV_reg_7_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in31_26,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_26
);
HV_reg_7_26_i_1 : CARRY4
 port map (
   CI => HV_reg_7_20_i_1_n_0,
   CYINIT => '0',
   DI(0) => h_24,
   DI(1) => h_25,
   DI(2) => h_26,
   DI(3) => h_27,
   S(0) => HV_7_26_i_5_n_0,
   S(1) => HV_7_26_i_4_n_0,
   S(2) => HV_7_26_i_3_n_0,
   S(3) => HV_7_26_i_2_n_0,
   CO(0) => HV_reg_7_26_i_1_n_3,
   CO(1) => HV_reg_7_26_i_1_n_2,
   CO(2) => HV_reg_7_26_i_1_n_1,
   CO(3) => HV_reg_7_26_i_1_n_0,
   O(0) => in31_24,
   O(1) => in31_25,
   O(2) => in31_26,
   O(3) => in31_27
);
HV_reg_7_27 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_7_27_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_27
);
HV_reg_7_28 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_7_28_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_28
);
HV_reg_7_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in31_29,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_29
);
HV_reg_7_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in31_2,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_2
);
HV_reg_7_2_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => h_0,
   DI(1) => h_1,
   DI(2) => h_2,
   DI(3) => h_3,
   S(0) => HV_7_2_i_5_n_0,
   S(1) => HV_7_2_i_4_n_0,
   S(2) => HV_7_2_i_3_n_0,
   S(3) => HV_7_2_i_2_n_0,
   CO(0) => HV_reg_7_2_i_1_n_3,
   CO(1) => HV_reg_7_2_i_1_n_2,
   CO(2) => HV_reg_7_2_i_1_n_1,
   CO(3) => HV_reg_7_2_i_1_n_0,
   O(0) => in31_0,
   O(1) => in31_1,
   O(2) => in31_2,
   O(3) => in31_3
);
HV_reg_7_30 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_7_30_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_30
);
HV_reg_7_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in31_31,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_31
);
HV_reg_7_31_i_1 : CARRY4
 port map (
   CI => HV_reg_7_26_i_1_n_0,
   CYINIT => '0',
   DI(0) => h_28,
   DI(1) => h_29,
   DI(2) => h_30,
   DI(3) => '0',
   S(0) => HV_7_31_i_5_n_0,
   S(1) => HV_7_31_i_4_n_0,
   S(2) => HV_7_31_i_3_n_0,
   S(3) => HV_7_31_i_2_n_0,
   CO(0) => HV_reg_7_31_i_1_n_3,
   CO(1) => HV_reg_7_31_i_1_n_2,
   CO(2) => HV_reg_7_31_i_1_n_1,
   CO(3) => NLW_HV_reg_7_31_i_1_CO_UNCONNECTED_3,
   O(0) => in31_28,
   O(1) => in31_29,
   O(2) => in31_30,
   O(3) => in31_31
);
HV_reg_7_3 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_7_3_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_3
);
HV_reg_7_4 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_7_4_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_4
);
HV_reg_7_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in31_5,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_5
);
HV_reg_7_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in31_6,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_6
);
HV_reg_7_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in31_7,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_7
);
HV_reg_7_7_i_1 : CARRY4
 port map (
   CI => HV_reg_7_2_i_1_n_0,
   CYINIT => '0',
   DI(0) => h_4,
   DI(1) => h_5,
   DI(2) => h_6,
   DI(3) => h_7,
   S(0) => HV_7_7_i_5_n_0,
   S(1) => HV_7_7_i_4_n_0,
   S(2) => HV_7_7_i_3_n_0,
   S(3) => HV_7_7_i_2_n_0,
   CO(0) => HV_reg_7_7_i_1_n_3,
   CO(1) => HV_reg_7_7_i_1_n_2,
   CO(2) => HV_reg_7_7_i_1_n_1,
   CO(3) => HV_reg_7_7_i_1_n_0,
   O(0) => in31_4,
   O(1) => in31_5,
   O(2) => in31_6,
   O(3) => in31_7
);
HV_reg_7_8 : FDSE
  generic map(
   INIT => '1'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => HV_7_8_i_1_n_0,
   S => HV_6_28_i_1_n_0,
   Q => data_out_OBUF_8
);
HV_reg_7_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => HV_reg_0_0,
   D => in31_9,
   R => HV_6_31_i_1_n_0,
   Q => data_out_OBUF_9
);
HV_reg_7_9_i_1 : CARRY4
 port map (
   CI => HV_reg_7_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => h_8,
   DI(1) => h_9,
   DI(2) => h_10,
   DI(3) => h_11,
   S(0) => HV_7_9_i_5_n_0,
   S(1) => HV_7_9_i_4_n_0,
   S(2) => HV_7_9_i_3_n_0,
   S(3) => HV_7_9_i_2_n_0,
   CO(0) => HV_reg_7_9_i_1_n_3,
   CO(1) => HV_reg_7_9_i_1_n_2,
   CO(2) => HV_reg_7_9_i_1_n_1,
   CO(3) => HV_reg_7_9_i_1_n_0,
   O(0) => in31_8,
   O(1) => in31_9,
   O(2) => in31_10,
   O(3) => in31_11
);
h_0_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => g_reg_n_0_0,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_0,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => h_0_i_1_n_0
);
h_10_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => g_reg_n_0_10,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_10,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => h_10_i_1_n_0
);
h_11_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => g_reg_n_0_11,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_11,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => h_11_i_1_n_0
);
h_12_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => g_reg_n_0_12,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_12,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => h_12_i_1_n_0
);
h_13_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => g_reg_n_0_13,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_13,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => h_13_i_1_n_0
);
h_14_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => g_reg_n_0_14,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_14,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => h_14_i_1_n_0
);
h_15_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => g_reg_n_0_15,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_15,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => h_15_i_1_n_0
);
h_16_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => g_reg_n_0_16,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_16,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => h_16_i_1_n_0
);
h_17_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => g_reg_n_0_17,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_17,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => h_17_i_1_n_0
);
h_18_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => g_reg_n_0_18,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_18,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => h_18_i_1_n_0
);
h_19_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => g_reg_n_0_19,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_19,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => h_19_i_1_n_0
);
h_1_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => g_reg_n_0_1,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_1,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => h_1_i_1_n_0
);
h_20_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => g_reg_n_0_20,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_20,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => h_20_i_1_n_0
);
h_21_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => g_reg_n_0_21,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_21,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => h_21_i_1_n_0
);
h_22_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => g_reg_n_0_22,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_22,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => h_22_i_1_n_0
);
h_23_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => g_reg_n_0_23,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_23,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => h_23_i_1_n_0
);
h_24_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => g_reg_n_0_24,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_24,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => h_24_i_1_n_0
);
h_25_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => g_reg_n_0_25,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_25,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => h_25_i_1_n_0
);
h_26_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => g_reg_n_0_26,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_26,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => h_26_i_1_n_0
);
h_27_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => g_reg_n_0_27,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_27,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => h_27_i_1_n_0
);
h_28_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => g_reg_n_0_28,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_28,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => h_28_i_1_n_0
);
h_29_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => g_reg_n_0_29,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_29,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => h_29_i_1_n_0
);
h_2_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => g_reg_n_0_2,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_2,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => h_2_i_1_n_0
);
h_30_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => g_reg_n_0_30,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_30,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => h_30_i_1_n_0
);
h_31_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => g_reg_n_0_31,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_31,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => h_31_i_1_n_0
);
h_3_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => g_reg_n_0_3,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_3,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => h_3_i_1_n_0
);
h_4_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => g_reg_n_0_4,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_4,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => h_4_i_1_n_0
);
h_5_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => g_reg_n_0_5,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_5,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => h_5_i_1_n_0
);
h_6_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => g_reg_n_0_6,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_6,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => h_6_i_1_n_0
);
h_7_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => g_reg_n_0_7,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_7,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => h_7_i_1_n_0
);
h_8_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => g_reg_n_0_8,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_8,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => h_8_i_1_n_0
);
h_9_i_1 : LUT4
  generic map(
   INIT => X"f888"
  )
 port map (
   I0 => g_reg_n_0_9,
   I1 => FSM_onehot_CURRENT_STATE_reg_n_0_11,
   I2 => data_out_OBUF_9,
   I3 => FSM_onehot_CURRENT_STATE_reg_n_0_7,
   O => h_9_i_1_n_0
);
h_reg_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => h_0_i_1_n_0,
   R => '0',
   Q => h_0
);
h_reg_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => h_10_i_1_n_0,
   R => '0',
   Q => h_10
);
h_reg_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => h_11_i_1_n_0,
   R => '0',
   Q => h_11
);
h_reg_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => h_12_i_1_n_0,
   R => '0',
   Q => h_12
);
h_reg_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => h_13_i_1_n_0,
   R => '0',
   Q => h_13
);
h_reg_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => h_14_i_1_n_0,
   R => '0',
   Q => h_14
);
h_reg_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => h_15_i_1_n_0,
   R => '0',
   Q => h_15
);
h_reg_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => h_16_i_1_n_0,
   R => '0',
   Q => h_16
);
h_reg_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => h_17_i_1_n_0,
   R => '0',
   Q => h_17
);
h_reg_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => h_18_i_1_n_0,
   R => '0',
   Q => h_18
);
h_reg_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => h_19_i_1_n_0,
   R => '0',
   Q => h_19
);
h_reg_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => h_1_i_1_n_0,
   R => '0',
   Q => h_1
);
h_reg_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => h_20_i_1_n_0,
   R => '0',
   Q => h_20
);
h_reg_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => h_21_i_1_n_0,
   R => '0',
   Q => h_21
);
h_reg_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => h_22_i_1_n_0,
   R => '0',
   Q => h_22
);
h_reg_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => h_23_i_1_n_0,
   R => '0',
   Q => h_23
);
h_reg_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => h_24_i_1_n_0,
   R => '0',
   Q => h_24
);
h_reg_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => h_25_i_1_n_0,
   R => '0',
   Q => h_25
);
h_reg_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => h_26_i_1_n_0,
   R => '0',
   Q => h_26
);
h_reg_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => h_27_i_1_n_0,
   R => '0',
   Q => h_27
);
h_reg_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => h_28_i_1_n_0,
   R => '0',
   Q => h_28
);
h_reg_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => h_29_i_1_n_0,
   R => '0',
   Q => h_29
);
h_reg_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => h_2_i_1_n_0,
   R => '0',
   Q => h_2
);
h_reg_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => h_30_i_1_n_0,
   R => '0',
   Q => h_30
);
h_reg_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => h_31_i_1_n_0,
   R => '0',
   Q => h_31
);
h_reg_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => h_3_i_1_n_0,
   R => '0',
   Q => h_3
);
h_reg_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => h_4_i_1_n_0,
   R => '0',
   Q => h_4
);
h_reg_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => h_5_i_1_n_0,
   R => '0',
   Q => h_5
);
h_reg_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => h_6_i_1_n_0,
   R => '0',
   Q => h_6
);
h_reg_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => h_7_i_1_n_0,
   R => '0',
   Q => h_7
);
h_reg_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => h_8_i_1_n_0,
   R => '0',
   Q => h_8
);
h_reg_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => a_31_i_1_n_0,
   D => h_9_i_1_n_0,
   R => '0',
   Q => h_9
);
msg_block_in_IBUF_0_inst : IBUF
 port map (
   I => msg_block_in_0,
   O => msg_block_in_IBUF_0
);
msg_block_in_IBUF_100_inst : IBUF
 port map (
   I => msg_block_in_100,
   O => msg_block_in_IBUF_100
);
msg_block_in_IBUF_101_inst : IBUF
 port map (
   I => msg_block_in_101,
   O => msg_block_in_IBUF_101
);
msg_block_in_IBUF_102_inst : IBUF
 port map (
   I => msg_block_in_102,
   O => msg_block_in_IBUF_102
);
msg_block_in_IBUF_103_inst : IBUF
 port map (
   I => msg_block_in_103,
   O => msg_block_in_IBUF_103
);
msg_block_in_IBUF_104_inst : IBUF
 port map (
   I => msg_block_in_104,
   O => msg_block_in_IBUF_104
);
msg_block_in_IBUF_105_inst : IBUF
 port map (
   I => msg_block_in_105,
   O => msg_block_in_IBUF_105
);
msg_block_in_IBUF_106_inst : IBUF
 port map (
   I => msg_block_in_106,
   O => msg_block_in_IBUF_106
);
msg_block_in_IBUF_107_inst : IBUF
 port map (
   I => msg_block_in_107,
   O => msg_block_in_IBUF_107
);
msg_block_in_IBUF_108_inst : IBUF
 port map (
   I => msg_block_in_108,
   O => msg_block_in_IBUF_108
);
msg_block_in_IBUF_109_inst : IBUF
 port map (
   I => msg_block_in_109,
   O => msg_block_in_IBUF_109
);
msg_block_in_IBUF_10_inst : IBUF
 port map (
   I => msg_block_in_10,
   O => msg_block_in_IBUF_10
);
msg_block_in_IBUF_110_inst : IBUF
 port map (
   I => msg_block_in_110,
   O => msg_block_in_IBUF_110
);
msg_block_in_IBUF_111_inst : IBUF
 port map (
   I => msg_block_in_111,
   O => msg_block_in_IBUF_111
);
msg_block_in_IBUF_112_inst : IBUF
 port map (
   I => msg_block_in_112,
   O => msg_block_in_IBUF_112
);
msg_block_in_IBUF_113_inst : IBUF
 port map (
   I => msg_block_in_113,
   O => msg_block_in_IBUF_113
);
msg_block_in_IBUF_114_inst : IBUF
 port map (
   I => msg_block_in_114,
   O => msg_block_in_IBUF_114
);
msg_block_in_IBUF_115_inst : IBUF
 port map (
   I => msg_block_in_115,
   O => msg_block_in_IBUF_115
);
msg_block_in_IBUF_116_inst : IBUF
 port map (
   I => msg_block_in_116,
   O => msg_block_in_IBUF_116
);
msg_block_in_IBUF_117_inst : IBUF
 port map (
   I => msg_block_in_117,
   O => msg_block_in_IBUF_117
);
msg_block_in_IBUF_118_inst : IBUF
 port map (
   I => msg_block_in_118,
   O => msg_block_in_IBUF_118
);
msg_block_in_IBUF_119_inst : IBUF
 port map (
   I => msg_block_in_119,
   O => msg_block_in_IBUF_119
);
msg_block_in_IBUF_11_inst : IBUF
 port map (
   I => msg_block_in_11,
   O => msg_block_in_IBUF_11
);
msg_block_in_IBUF_120_inst : IBUF
 port map (
   I => msg_block_in_120,
   O => msg_block_in_IBUF_120
);
msg_block_in_IBUF_121_inst : IBUF
 port map (
   I => msg_block_in_121,
   O => msg_block_in_IBUF_121
);
msg_block_in_IBUF_122_inst : IBUF
 port map (
   I => msg_block_in_122,
   O => msg_block_in_IBUF_122
);
msg_block_in_IBUF_123_inst : IBUF
 port map (
   I => msg_block_in_123,
   O => msg_block_in_IBUF_123
);
msg_block_in_IBUF_124_inst : IBUF
 port map (
   I => msg_block_in_124,
   O => msg_block_in_IBUF_124
);
msg_block_in_IBUF_125_inst : IBUF
 port map (
   I => msg_block_in_125,
   O => msg_block_in_IBUF_125
);
msg_block_in_IBUF_126_inst : IBUF
 port map (
   I => msg_block_in_126,
   O => msg_block_in_IBUF_126
);
msg_block_in_IBUF_127_inst : IBUF
 port map (
   I => msg_block_in_127,
   O => msg_block_in_IBUF_127
);
msg_block_in_IBUF_128_inst : IBUF
 port map (
   I => msg_block_in_128,
   O => msg_block_in_IBUF_128
);
msg_block_in_IBUF_129_inst : IBUF
 port map (
   I => msg_block_in_129,
   O => msg_block_in_IBUF_129
);
msg_block_in_IBUF_12_inst : IBUF
 port map (
   I => msg_block_in_12,
   O => msg_block_in_IBUF_12
);
msg_block_in_IBUF_130_inst : IBUF
 port map (
   I => msg_block_in_130,
   O => msg_block_in_IBUF_130
);
msg_block_in_IBUF_131_inst : IBUF
 port map (
   I => msg_block_in_131,
   O => msg_block_in_IBUF_131
);
msg_block_in_IBUF_132_inst : IBUF
 port map (
   I => msg_block_in_132,
   O => msg_block_in_IBUF_132
);
msg_block_in_IBUF_133_inst : IBUF
 port map (
   I => msg_block_in_133,
   O => msg_block_in_IBUF_133
);
msg_block_in_IBUF_134_inst : IBUF
 port map (
   I => msg_block_in_134,
   O => msg_block_in_IBUF_134
);
msg_block_in_IBUF_135_inst : IBUF
 port map (
   I => msg_block_in_135,
   O => msg_block_in_IBUF_135
);
msg_block_in_IBUF_136_inst : IBUF
 port map (
   I => msg_block_in_136,
   O => msg_block_in_IBUF_136
);
msg_block_in_IBUF_137_inst : IBUF
 port map (
   I => msg_block_in_137,
   O => msg_block_in_IBUF_137
);
msg_block_in_IBUF_138_inst : IBUF
 port map (
   I => msg_block_in_138,
   O => msg_block_in_IBUF_138
);
msg_block_in_IBUF_139_inst : IBUF
 port map (
   I => msg_block_in_139,
   O => msg_block_in_IBUF_139
);
msg_block_in_IBUF_13_inst : IBUF
 port map (
   I => msg_block_in_13,
   O => msg_block_in_IBUF_13
);
msg_block_in_IBUF_140_inst : IBUF
 port map (
   I => msg_block_in_140,
   O => msg_block_in_IBUF_140
);
msg_block_in_IBUF_141_inst : IBUF
 port map (
   I => msg_block_in_141,
   O => msg_block_in_IBUF_141
);
msg_block_in_IBUF_142_inst : IBUF
 port map (
   I => msg_block_in_142,
   O => msg_block_in_IBUF_142
);
msg_block_in_IBUF_143_inst : IBUF
 port map (
   I => msg_block_in_143,
   O => msg_block_in_IBUF_143
);
msg_block_in_IBUF_144_inst : IBUF
 port map (
   I => msg_block_in_144,
   O => msg_block_in_IBUF_144
);
msg_block_in_IBUF_145_inst : IBUF
 port map (
   I => msg_block_in_145,
   O => msg_block_in_IBUF_145
);
msg_block_in_IBUF_146_inst : IBUF
 port map (
   I => msg_block_in_146,
   O => msg_block_in_IBUF_146
);
msg_block_in_IBUF_147_inst : IBUF
 port map (
   I => msg_block_in_147,
   O => msg_block_in_IBUF_147
);
msg_block_in_IBUF_148_inst : IBUF
 port map (
   I => msg_block_in_148,
   O => msg_block_in_IBUF_148
);
msg_block_in_IBUF_149_inst : IBUF
 port map (
   I => msg_block_in_149,
   O => msg_block_in_IBUF_149
);
msg_block_in_IBUF_14_inst : IBUF
 port map (
   I => msg_block_in_14,
   O => msg_block_in_IBUF_14
);
msg_block_in_IBUF_150_inst : IBUF
 port map (
   I => msg_block_in_150,
   O => msg_block_in_IBUF_150
);
msg_block_in_IBUF_151_inst : IBUF
 port map (
   I => msg_block_in_151,
   O => msg_block_in_IBUF_151
);
msg_block_in_IBUF_152_inst : IBUF
 port map (
   I => msg_block_in_152,
   O => msg_block_in_IBUF_152
);
msg_block_in_IBUF_153_inst : IBUF
 port map (
   I => msg_block_in_153,
   O => msg_block_in_IBUF_153
);
msg_block_in_IBUF_154_inst : IBUF
 port map (
   I => msg_block_in_154,
   O => msg_block_in_IBUF_154
);
msg_block_in_IBUF_155_inst : IBUF
 port map (
   I => msg_block_in_155,
   O => msg_block_in_IBUF_155
);
msg_block_in_IBUF_156_inst : IBUF
 port map (
   I => msg_block_in_156,
   O => msg_block_in_IBUF_156
);
msg_block_in_IBUF_157_inst : IBUF
 port map (
   I => msg_block_in_157,
   O => msg_block_in_IBUF_157
);
msg_block_in_IBUF_158_inst : IBUF
 port map (
   I => msg_block_in_158,
   O => msg_block_in_IBUF_158
);
msg_block_in_IBUF_159_inst : IBUF
 port map (
   I => msg_block_in_159,
   O => msg_block_in_IBUF_159
);
msg_block_in_IBUF_15_inst : IBUF
 port map (
   I => msg_block_in_15,
   O => msg_block_in_IBUF_15
);
msg_block_in_IBUF_160_inst : IBUF
 port map (
   I => msg_block_in_160,
   O => msg_block_in_IBUF_160
);
msg_block_in_IBUF_161_inst : IBUF
 port map (
   I => msg_block_in_161,
   O => msg_block_in_IBUF_161
);
msg_block_in_IBUF_162_inst : IBUF
 port map (
   I => msg_block_in_162,
   O => msg_block_in_IBUF_162
);
msg_block_in_IBUF_163_inst : IBUF
 port map (
   I => msg_block_in_163,
   O => msg_block_in_IBUF_163
);
msg_block_in_IBUF_164_inst : IBUF
 port map (
   I => msg_block_in_164,
   O => msg_block_in_IBUF_164
);
msg_block_in_IBUF_165_inst : IBUF
 port map (
   I => msg_block_in_165,
   O => msg_block_in_IBUF_165
);
msg_block_in_IBUF_166_inst : IBUF
 port map (
   I => msg_block_in_166,
   O => msg_block_in_IBUF_166
);
msg_block_in_IBUF_167_inst : IBUF
 port map (
   I => msg_block_in_167,
   O => msg_block_in_IBUF_167
);
msg_block_in_IBUF_168_inst : IBUF
 port map (
   I => msg_block_in_168,
   O => msg_block_in_IBUF_168
);
msg_block_in_IBUF_169_inst : IBUF
 port map (
   I => msg_block_in_169,
   O => msg_block_in_IBUF_169
);
msg_block_in_IBUF_16_inst : IBUF
 port map (
   I => msg_block_in_16,
   O => msg_block_in_IBUF_16
);
msg_block_in_IBUF_170_inst : IBUF
 port map (
   I => msg_block_in_170,
   O => msg_block_in_IBUF_170
);
msg_block_in_IBUF_171_inst : IBUF
 port map (
   I => msg_block_in_171,
   O => msg_block_in_IBUF_171
);
msg_block_in_IBUF_172_inst : IBUF
 port map (
   I => msg_block_in_172,
   O => msg_block_in_IBUF_172
);
msg_block_in_IBUF_173_inst : IBUF
 port map (
   I => msg_block_in_173,
   O => msg_block_in_IBUF_173
);
msg_block_in_IBUF_174_inst : IBUF
 port map (
   I => msg_block_in_174,
   O => msg_block_in_IBUF_174
);
msg_block_in_IBUF_175_inst : IBUF
 port map (
   I => msg_block_in_175,
   O => msg_block_in_IBUF_175
);
msg_block_in_IBUF_176_inst : IBUF
 port map (
   I => msg_block_in_176,
   O => msg_block_in_IBUF_176
);
msg_block_in_IBUF_177_inst : IBUF
 port map (
   I => msg_block_in_177,
   O => msg_block_in_IBUF_177
);
msg_block_in_IBUF_178_inst : IBUF
 port map (
   I => msg_block_in_178,
   O => msg_block_in_IBUF_178
);
msg_block_in_IBUF_179_inst : IBUF
 port map (
   I => msg_block_in_179,
   O => msg_block_in_IBUF_179
);
msg_block_in_IBUF_17_inst : IBUF
 port map (
   I => msg_block_in_17,
   O => msg_block_in_IBUF_17
);
msg_block_in_IBUF_180_inst : IBUF
 port map (
   I => msg_block_in_180,
   O => msg_block_in_IBUF_180
);
msg_block_in_IBUF_181_inst : IBUF
 port map (
   I => msg_block_in_181,
   O => msg_block_in_IBUF_181
);
msg_block_in_IBUF_182_inst : IBUF
 port map (
   I => msg_block_in_182,
   O => msg_block_in_IBUF_182
);
msg_block_in_IBUF_183_inst : IBUF
 port map (
   I => msg_block_in_183,
   O => msg_block_in_IBUF_183
);
msg_block_in_IBUF_184_inst : IBUF
 port map (
   I => msg_block_in_184,
   O => msg_block_in_IBUF_184
);
msg_block_in_IBUF_185_inst : IBUF
 port map (
   I => msg_block_in_185,
   O => msg_block_in_IBUF_185
);
msg_block_in_IBUF_186_inst : IBUF
 port map (
   I => msg_block_in_186,
   O => msg_block_in_IBUF_186
);
msg_block_in_IBUF_187_inst : IBUF
 port map (
   I => msg_block_in_187,
   O => msg_block_in_IBUF_187
);
msg_block_in_IBUF_188_inst : IBUF
 port map (
   I => msg_block_in_188,
   O => msg_block_in_IBUF_188
);
msg_block_in_IBUF_189_inst : IBUF
 port map (
   I => msg_block_in_189,
   O => msg_block_in_IBUF_189
);
msg_block_in_IBUF_18_inst : IBUF
 port map (
   I => msg_block_in_18,
   O => msg_block_in_IBUF_18
);
msg_block_in_IBUF_190_inst : IBUF
 port map (
   I => msg_block_in_190,
   O => msg_block_in_IBUF_190
);
msg_block_in_IBUF_191_inst : IBUF
 port map (
   I => msg_block_in_191,
   O => msg_block_in_IBUF_191
);
msg_block_in_IBUF_192_inst : IBUF
 port map (
   I => msg_block_in_192,
   O => msg_block_in_IBUF_192
);
msg_block_in_IBUF_193_inst : IBUF
 port map (
   I => msg_block_in_193,
   O => msg_block_in_IBUF_193
);
msg_block_in_IBUF_194_inst : IBUF
 port map (
   I => msg_block_in_194,
   O => msg_block_in_IBUF_194
);
msg_block_in_IBUF_195_inst : IBUF
 port map (
   I => msg_block_in_195,
   O => msg_block_in_IBUF_195
);
msg_block_in_IBUF_196_inst : IBUF
 port map (
   I => msg_block_in_196,
   O => msg_block_in_IBUF_196
);
msg_block_in_IBUF_197_inst : IBUF
 port map (
   I => msg_block_in_197,
   O => msg_block_in_IBUF_197
);
msg_block_in_IBUF_198_inst : IBUF
 port map (
   I => msg_block_in_198,
   O => msg_block_in_IBUF_198
);
msg_block_in_IBUF_199_inst : IBUF
 port map (
   I => msg_block_in_199,
   O => msg_block_in_IBUF_199
);
msg_block_in_IBUF_19_inst : IBUF
 port map (
   I => msg_block_in_19,
   O => msg_block_in_IBUF_19
);
msg_block_in_IBUF_1_inst : IBUF
 port map (
   I => msg_block_in_1,
   O => msg_block_in_IBUF_1
);
msg_block_in_IBUF_200_inst : IBUF
 port map (
   I => msg_block_in_200,
   O => msg_block_in_IBUF_200
);
msg_block_in_IBUF_201_inst : IBUF
 port map (
   I => msg_block_in_201,
   O => msg_block_in_IBUF_201
);
msg_block_in_IBUF_202_inst : IBUF
 port map (
   I => msg_block_in_202,
   O => msg_block_in_IBUF_202
);
msg_block_in_IBUF_203_inst : IBUF
 port map (
   I => msg_block_in_203,
   O => msg_block_in_IBUF_203
);
msg_block_in_IBUF_204_inst : IBUF
 port map (
   I => msg_block_in_204,
   O => msg_block_in_IBUF_204
);
msg_block_in_IBUF_205_inst : IBUF
 port map (
   I => msg_block_in_205,
   O => msg_block_in_IBUF_205
);
msg_block_in_IBUF_206_inst : IBUF
 port map (
   I => msg_block_in_206,
   O => msg_block_in_IBUF_206
);
msg_block_in_IBUF_207_inst : IBUF
 port map (
   I => msg_block_in_207,
   O => msg_block_in_IBUF_207
);
msg_block_in_IBUF_208_inst : IBUF
 port map (
   I => msg_block_in_208,
   O => msg_block_in_IBUF_208
);
msg_block_in_IBUF_209_inst : IBUF
 port map (
   I => msg_block_in_209,
   O => msg_block_in_IBUF_209
);
msg_block_in_IBUF_20_inst : IBUF
 port map (
   I => msg_block_in_20,
   O => msg_block_in_IBUF_20
);
msg_block_in_IBUF_210_inst : IBUF
 port map (
   I => msg_block_in_210,
   O => msg_block_in_IBUF_210
);
msg_block_in_IBUF_211_inst : IBUF
 port map (
   I => msg_block_in_211,
   O => msg_block_in_IBUF_211
);
msg_block_in_IBUF_212_inst : IBUF
 port map (
   I => msg_block_in_212,
   O => msg_block_in_IBUF_212
);
msg_block_in_IBUF_213_inst : IBUF
 port map (
   I => msg_block_in_213,
   O => msg_block_in_IBUF_213
);
msg_block_in_IBUF_214_inst : IBUF
 port map (
   I => msg_block_in_214,
   O => msg_block_in_IBUF_214
);
msg_block_in_IBUF_215_inst : IBUF
 port map (
   I => msg_block_in_215,
   O => msg_block_in_IBUF_215
);
msg_block_in_IBUF_216_inst : IBUF
 port map (
   I => msg_block_in_216,
   O => msg_block_in_IBUF_216
);
msg_block_in_IBUF_217_inst : IBUF
 port map (
   I => msg_block_in_217,
   O => msg_block_in_IBUF_217
);
msg_block_in_IBUF_218_inst : IBUF
 port map (
   I => msg_block_in_218,
   O => msg_block_in_IBUF_218
);
msg_block_in_IBUF_219_inst : IBUF
 port map (
   I => msg_block_in_219,
   O => msg_block_in_IBUF_219
);
msg_block_in_IBUF_21_inst : IBUF
 port map (
   I => msg_block_in_21,
   O => msg_block_in_IBUF_21
);
msg_block_in_IBUF_220_inst : IBUF
 port map (
   I => msg_block_in_220,
   O => msg_block_in_IBUF_220
);
msg_block_in_IBUF_221_inst : IBUF
 port map (
   I => msg_block_in_221,
   O => msg_block_in_IBUF_221
);
msg_block_in_IBUF_222_inst : IBUF
 port map (
   I => msg_block_in_222,
   O => msg_block_in_IBUF_222
);
msg_block_in_IBUF_223_inst : IBUF
 port map (
   I => msg_block_in_223,
   O => msg_block_in_IBUF_223
);
msg_block_in_IBUF_224_inst : IBUF
 port map (
   I => msg_block_in_224,
   O => msg_block_in_IBUF_224
);
msg_block_in_IBUF_225_inst : IBUF
 port map (
   I => msg_block_in_225,
   O => msg_block_in_IBUF_225
);
msg_block_in_IBUF_226_inst : IBUF
 port map (
   I => msg_block_in_226,
   O => msg_block_in_IBUF_226
);
msg_block_in_IBUF_227_inst : IBUF
 port map (
   I => msg_block_in_227,
   O => msg_block_in_IBUF_227
);
msg_block_in_IBUF_228_inst : IBUF
 port map (
   I => msg_block_in_228,
   O => msg_block_in_IBUF_228
);
msg_block_in_IBUF_229_inst : IBUF
 port map (
   I => msg_block_in_229,
   O => msg_block_in_IBUF_229
);
msg_block_in_IBUF_22_inst : IBUF
 port map (
   I => msg_block_in_22,
   O => msg_block_in_IBUF_22
);
msg_block_in_IBUF_230_inst : IBUF
 port map (
   I => msg_block_in_230,
   O => msg_block_in_IBUF_230
);
msg_block_in_IBUF_231_inst : IBUF
 port map (
   I => msg_block_in_231,
   O => msg_block_in_IBUF_231
);
msg_block_in_IBUF_232_inst : IBUF
 port map (
   I => msg_block_in_232,
   O => msg_block_in_IBUF_232
);
msg_block_in_IBUF_233_inst : IBUF
 port map (
   I => msg_block_in_233,
   O => msg_block_in_IBUF_233
);
msg_block_in_IBUF_234_inst : IBUF
 port map (
   I => msg_block_in_234,
   O => msg_block_in_IBUF_234
);
msg_block_in_IBUF_235_inst : IBUF
 port map (
   I => msg_block_in_235,
   O => msg_block_in_IBUF_235
);
msg_block_in_IBUF_236_inst : IBUF
 port map (
   I => msg_block_in_236,
   O => msg_block_in_IBUF_236
);
msg_block_in_IBUF_237_inst : IBUF
 port map (
   I => msg_block_in_237,
   O => msg_block_in_IBUF_237
);
msg_block_in_IBUF_238_inst : IBUF
 port map (
   I => msg_block_in_238,
   O => msg_block_in_IBUF_238
);
msg_block_in_IBUF_239_inst : IBUF
 port map (
   I => msg_block_in_239,
   O => msg_block_in_IBUF_239
);
msg_block_in_IBUF_23_inst : IBUF
 port map (
   I => msg_block_in_23,
   O => msg_block_in_IBUF_23
);
msg_block_in_IBUF_240_inst : IBUF
 port map (
   I => msg_block_in_240,
   O => msg_block_in_IBUF_240
);
msg_block_in_IBUF_241_inst : IBUF
 port map (
   I => msg_block_in_241,
   O => msg_block_in_IBUF_241
);
msg_block_in_IBUF_242_inst : IBUF
 port map (
   I => msg_block_in_242,
   O => msg_block_in_IBUF_242
);
msg_block_in_IBUF_243_inst : IBUF
 port map (
   I => msg_block_in_243,
   O => msg_block_in_IBUF_243
);
msg_block_in_IBUF_244_inst : IBUF
 port map (
   I => msg_block_in_244,
   O => msg_block_in_IBUF_244
);
msg_block_in_IBUF_245_inst : IBUF
 port map (
   I => msg_block_in_245,
   O => msg_block_in_IBUF_245
);
msg_block_in_IBUF_246_inst : IBUF
 port map (
   I => msg_block_in_246,
   O => msg_block_in_IBUF_246
);
msg_block_in_IBUF_247_inst : IBUF
 port map (
   I => msg_block_in_247,
   O => msg_block_in_IBUF_247
);
msg_block_in_IBUF_248_inst : IBUF
 port map (
   I => msg_block_in_248,
   O => msg_block_in_IBUF_248
);
msg_block_in_IBUF_249_inst : IBUF
 port map (
   I => msg_block_in_249,
   O => msg_block_in_IBUF_249
);
msg_block_in_IBUF_24_inst : IBUF
 port map (
   I => msg_block_in_24,
   O => msg_block_in_IBUF_24
);
msg_block_in_IBUF_250_inst : IBUF
 port map (
   I => msg_block_in_250,
   O => msg_block_in_IBUF_250
);
msg_block_in_IBUF_251_inst : IBUF
 port map (
   I => msg_block_in_251,
   O => msg_block_in_IBUF_251
);
msg_block_in_IBUF_252_inst : IBUF
 port map (
   I => msg_block_in_252,
   O => msg_block_in_IBUF_252
);
msg_block_in_IBUF_253_inst : IBUF
 port map (
   I => msg_block_in_253,
   O => msg_block_in_IBUF_253
);
msg_block_in_IBUF_254_inst : IBUF
 port map (
   I => msg_block_in_254,
   O => msg_block_in_IBUF_254
);
msg_block_in_IBUF_255_inst : IBUF
 port map (
   I => msg_block_in_255,
   O => msg_block_in_IBUF_255
);
msg_block_in_IBUF_256_inst : IBUF
 port map (
   I => msg_block_in_256,
   O => msg_block_in_IBUF_256
);
msg_block_in_IBUF_257_inst : IBUF
 port map (
   I => msg_block_in_257,
   O => msg_block_in_IBUF_257
);
msg_block_in_IBUF_258_inst : IBUF
 port map (
   I => msg_block_in_258,
   O => msg_block_in_IBUF_258
);
msg_block_in_IBUF_259_inst : IBUF
 port map (
   I => msg_block_in_259,
   O => msg_block_in_IBUF_259
);
msg_block_in_IBUF_25_inst : IBUF
 port map (
   I => msg_block_in_25,
   O => msg_block_in_IBUF_25
);
msg_block_in_IBUF_260_inst : IBUF
 port map (
   I => msg_block_in_260,
   O => msg_block_in_IBUF_260
);
msg_block_in_IBUF_261_inst : IBUF
 port map (
   I => msg_block_in_261,
   O => msg_block_in_IBUF_261
);
msg_block_in_IBUF_262_inst : IBUF
 port map (
   I => msg_block_in_262,
   O => msg_block_in_IBUF_262
);
msg_block_in_IBUF_263_inst : IBUF
 port map (
   I => msg_block_in_263,
   O => msg_block_in_IBUF_263
);
msg_block_in_IBUF_264_inst : IBUF
 port map (
   I => msg_block_in_264,
   O => msg_block_in_IBUF_264
);
msg_block_in_IBUF_265_inst : IBUF
 port map (
   I => msg_block_in_265,
   O => msg_block_in_IBUF_265
);
msg_block_in_IBUF_266_inst : IBUF
 port map (
   I => msg_block_in_266,
   O => msg_block_in_IBUF_266
);
msg_block_in_IBUF_267_inst : IBUF
 port map (
   I => msg_block_in_267,
   O => msg_block_in_IBUF_267
);
msg_block_in_IBUF_268_inst : IBUF
 port map (
   I => msg_block_in_268,
   O => msg_block_in_IBUF_268
);
msg_block_in_IBUF_269_inst : IBUF
 port map (
   I => msg_block_in_269,
   O => msg_block_in_IBUF_269
);
msg_block_in_IBUF_26_inst : IBUF
 port map (
   I => msg_block_in_26,
   O => msg_block_in_IBUF_26
);
msg_block_in_IBUF_270_inst : IBUF
 port map (
   I => msg_block_in_270,
   O => msg_block_in_IBUF_270
);
msg_block_in_IBUF_271_inst : IBUF
 port map (
   I => msg_block_in_271,
   O => msg_block_in_IBUF_271
);
msg_block_in_IBUF_272_inst : IBUF
 port map (
   I => msg_block_in_272,
   O => msg_block_in_IBUF_272
);
msg_block_in_IBUF_273_inst : IBUF
 port map (
   I => msg_block_in_273,
   O => msg_block_in_IBUF_273
);
msg_block_in_IBUF_274_inst : IBUF
 port map (
   I => msg_block_in_274,
   O => msg_block_in_IBUF_274
);
msg_block_in_IBUF_275_inst : IBUF
 port map (
   I => msg_block_in_275,
   O => msg_block_in_IBUF_275
);
msg_block_in_IBUF_276_inst : IBUF
 port map (
   I => msg_block_in_276,
   O => msg_block_in_IBUF_276
);
msg_block_in_IBUF_277_inst : IBUF
 port map (
   I => msg_block_in_277,
   O => msg_block_in_IBUF_277
);
msg_block_in_IBUF_278_inst : IBUF
 port map (
   I => msg_block_in_278,
   O => msg_block_in_IBUF_278
);
msg_block_in_IBUF_279_inst : IBUF
 port map (
   I => msg_block_in_279,
   O => msg_block_in_IBUF_279
);
msg_block_in_IBUF_27_inst : IBUF
 port map (
   I => msg_block_in_27,
   O => msg_block_in_IBUF_27
);
msg_block_in_IBUF_280_inst : IBUF
 port map (
   I => msg_block_in_280,
   O => msg_block_in_IBUF_280
);
msg_block_in_IBUF_281_inst : IBUF
 port map (
   I => msg_block_in_281,
   O => msg_block_in_IBUF_281
);
msg_block_in_IBUF_282_inst : IBUF
 port map (
   I => msg_block_in_282,
   O => msg_block_in_IBUF_282
);
msg_block_in_IBUF_283_inst : IBUF
 port map (
   I => msg_block_in_283,
   O => msg_block_in_IBUF_283
);
msg_block_in_IBUF_284_inst : IBUF
 port map (
   I => msg_block_in_284,
   O => msg_block_in_IBUF_284
);
msg_block_in_IBUF_285_inst : IBUF
 port map (
   I => msg_block_in_285,
   O => msg_block_in_IBUF_285
);
msg_block_in_IBUF_286_inst : IBUF
 port map (
   I => msg_block_in_286,
   O => msg_block_in_IBUF_286
);
msg_block_in_IBUF_287_inst : IBUF
 port map (
   I => msg_block_in_287,
   O => msg_block_in_IBUF_287
);
msg_block_in_IBUF_288_inst : IBUF
 port map (
   I => msg_block_in_288,
   O => msg_block_in_IBUF_288
);
msg_block_in_IBUF_289_inst : IBUF
 port map (
   I => msg_block_in_289,
   O => msg_block_in_IBUF_289
);
msg_block_in_IBUF_28_inst : IBUF
 port map (
   I => msg_block_in_28,
   O => msg_block_in_IBUF_28
);
msg_block_in_IBUF_290_inst : IBUF
 port map (
   I => msg_block_in_290,
   O => msg_block_in_IBUF_290
);
msg_block_in_IBUF_291_inst : IBUF
 port map (
   I => msg_block_in_291,
   O => msg_block_in_IBUF_291
);
msg_block_in_IBUF_292_inst : IBUF
 port map (
   I => msg_block_in_292,
   O => msg_block_in_IBUF_292
);
msg_block_in_IBUF_293_inst : IBUF
 port map (
   I => msg_block_in_293,
   O => msg_block_in_IBUF_293
);
msg_block_in_IBUF_294_inst : IBUF
 port map (
   I => msg_block_in_294,
   O => msg_block_in_IBUF_294
);
msg_block_in_IBUF_295_inst : IBUF
 port map (
   I => msg_block_in_295,
   O => msg_block_in_IBUF_295
);
msg_block_in_IBUF_296_inst : IBUF
 port map (
   I => msg_block_in_296,
   O => msg_block_in_IBUF_296
);
msg_block_in_IBUF_297_inst : IBUF
 port map (
   I => msg_block_in_297,
   O => msg_block_in_IBUF_297
);
msg_block_in_IBUF_298_inst : IBUF
 port map (
   I => msg_block_in_298,
   O => msg_block_in_IBUF_298
);
msg_block_in_IBUF_299_inst : IBUF
 port map (
   I => msg_block_in_299,
   O => msg_block_in_IBUF_299
);
msg_block_in_IBUF_29_inst : IBUF
 port map (
   I => msg_block_in_29,
   O => msg_block_in_IBUF_29
);
msg_block_in_IBUF_2_inst : IBUF
 port map (
   I => msg_block_in_2,
   O => msg_block_in_IBUF_2
);
msg_block_in_IBUF_300_inst : IBUF
 port map (
   I => msg_block_in_300,
   O => msg_block_in_IBUF_300
);
msg_block_in_IBUF_301_inst : IBUF
 port map (
   I => msg_block_in_301,
   O => msg_block_in_IBUF_301
);
msg_block_in_IBUF_302_inst : IBUF
 port map (
   I => msg_block_in_302,
   O => msg_block_in_IBUF_302
);
msg_block_in_IBUF_303_inst : IBUF
 port map (
   I => msg_block_in_303,
   O => msg_block_in_IBUF_303
);
msg_block_in_IBUF_304_inst : IBUF
 port map (
   I => msg_block_in_304,
   O => msg_block_in_IBUF_304
);
msg_block_in_IBUF_305_inst : IBUF
 port map (
   I => msg_block_in_305,
   O => msg_block_in_IBUF_305
);
msg_block_in_IBUF_306_inst : IBUF
 port map (
   I => msg_block_in_306,
   O => msg_block_in_IBUF_306
);
msg_block_in_IBUF_307_inst : IBUF
 port map (
   I => msg_block_in_307,
   O => msg_block_in_IBUF_307
);
msg_block_in_IBUF_308_inst : IBUF
 port map (
   I => msg_block_in_308,
   O => msg_block_in_IBUF_308
);
msg_block_in_IBUF_309_inst : IBUF
 port map (
   I => msg_block_in_309,
   O => msg_block_in_IBUF_309
);
msg_block_in_IBUF_30_inst : IBUF
 port map (
   I => msg_block_in_30,
   O => msg_block_in_IBUF_30
);
msg_block_in_IBUF_310_inst : IBUF
 port map (
   I => msg_block_in_310,
   O => msg_block_in_IBUF_310
);
msg_block_in_IBUF_311_inst : IBUF
 port map (
   I => msg_block_in_311,
   O => msg_block_in_IBUF_311
);
msg_block_in_IBUF_312_inst : IBUF
 port map (
   I => msg_block_in_312,
   O => msg_block_in_IBUF_312
);
msg_block_in_IBUF_313_inst : IBUF
 port map (
   I => msg_block_in_313,
   O => msg_block_in_IBUF_313
);
msg_block_in_IBUF_314_inst : IBUF
 port map (
   I => msg_block_in_314,
   O => msg_block_in_IBUF_314
);
msg_block_in_IBUF_315_inst : IBUF
 port map (
   I => msg_block_in_315,
   O => msg_block_in_IBUF_315
);
msg_block_in_IBUF_316_inst : IBUF
 port map (
   I => msg_block_in_316,
   O => msg_block_in_IBUF_316
);
msg_block_in_IBUF_317_inst : IBUF
 port map (
   I => msg_block_in_317,
   O => msg_block_in_IBUF_317
);
msg_block_in_IBUF_318_inst : IBUF
 port map (
   I => msg_block_in_318,
   O => msg_block_in_IBUF_318
);
msg_block_in_IBUF_319_inst : IBUF
 port map (
   I => msg_block_in_319,
   O => msg_block_in_IBUF_319
);
msg_block_in_IBUF_31_inst : IBUF
 port map (
   I => msg_block_in_31,
   O => msg_block_in_IBUF_31
);
msg_block_in_IBUF_320_inst : IBUF
 port map (
   I => msg_block_in_320,
   O => msg_block_in_IBUF_320
);
msg_block_in_IBUF_321_inst : IBUF
 port map (
   I => msg_block_in_321,
   O => msg_block_in_IBUF_321
);
msg_block_in_IBUF_322_inst : IBUF
 port map (
   I => msg_block_in_322,
   O => msg_block_in_IBUF_322
);
msg_block_in_IBUF_323_inst : IBUF
 port map (
   I => msg_block_in_323,
   O => msg_block_in_IBUF_323
);
msg_block_in_IBUF_324_inst : IBUF
 port map (
   I => msg_block_in_324,
   O => msg_block_in_IBUF_324
);
msg_block_in_IBUF_325_inst : IBUF
 port map (
   I => msg_block_in_325,
   O => msg_block_in_IBUF_325
);
msg_block_in_IBUF_326_inst : IBUF
 port map (
   I => msg_block_in_326,
   O => msg_block_in_IBUF_326
);
msg_block_in_IBUF_327_inst : IBUF
 port map (
   I => msg_block_in_327,
   O => msg_block_in_IBUF_327
);
msg_block_in_IBUF_328_inst : IBUF
 port map (
   I => msg_block_in_328,
   O => msg_block_in_IBUF_328
);
msg_block_in_IBUF_329_inst : IBUF
 port map (
   I => msg_block_in_329,
   O => msg_block_in_IBUF_329
);
msg_block_in_IBUF_32_inst : IBUF
 port map (
   I => msg_block_in_32,
   O => msg_block_in_IBUF_32
);
msg_block_in_IBUF_330_inst : IBUF
 port map (
   I => msg_block_in_330,
   O => msg_block_in_IBUF_330
);
msg_block_in_IBUF_331_inst : IBUF
 port map (
   I => msg_block_in_331,
   O => msg_block_in_IBUF_331
);
msg_block_in_IBUF_332_inst : IBUF
 port map (
   I => msg_block_in_332,
   O => msg_block_in_IBUF_332
);
msg_block_in_IBUF_333_inst : IBUF
 port map (
   I => msg_block_in_333,
   O => msg_block_in_IBUF_333
);
msg_block_in_IBUF_334_inst : IBUF
 port map (
   I => msg_block_in_334,
   O => msg_block_in_IBUF_334
);
msg_block_in_IBUF_335_inst : IBUF
 port map (
   I => msg_block_in_335,
   O => msg_block_in_IBUF_335
);
msg_block_in_IBUF_336_inst : IBUF
 port map (
   I => msg_block_in_336,
   O => msg_block_in_IBUF_336
);
msg_block_in_IBUF_337_inst : IBUF
 port map (
   I => msg_block_in_337,
   O => msg_block_in_IBUF_337
);
msg_block_in_IBUF_338_inst : IBUF
 port map (
   I => msg_block_in_338,
   O => msg_block_in_IBUF_338
);
msg_block_in_IBUF_339_inst : IBUF
 port map (
   I => msg_block_in_339,
   O => msg_block_in_IBUF_339
);
msg_block_in_IBUF_33_inst : IBUF
 port map (
   I => msg_block_in_33,
   O => msg_block_in_IBUF_33
);
msg_block_in_IBUF_340_inst : IBUF
 port map (
   I => msg_block_in_340,
   O => msg_block_in_IBUF_340
);
msg_block_in_IBUF_341_inst : IBUF
 port map (
   I => msg_block_in_341,
   O => msg_block_in_IBUF_341
);
msg_block_in_IBUF_342_inst : IBUF
 port map (
   I => msg_block_in_342,
   O => msg_block_in_IBUF_342
);
msg_block_in_IBUF_343_inst : IBUF
 port map (
   I => msg_block_in_343,
   O => msg_block_in_IBUF_343
);
msg_block_in_IBUF_344_inst : IBUF
 port map (
   I => msg_block_in_344,
   O => msg_block_in_IBUF_344
);
msg_block_in_IBUF_345_inst : IBUF
 port map (
   I => msg_block_in_345,
   O => msg_block_in_IBUF_345
);
msg_block_in_IBUF_346_inst : IBUF
 port map (
   I => msg_block_in_346,
   O => msg_block_in_IBUF_346
);
msg_block_in_IBUF_347_inst : IBUF
 port map (
   I => msg_block_in_347,
   O => msg_block_in_IBUF_347
);
msg_block_in_IBUF_348_inst : IBUF
 port map (
   I => msg_block_in_348,
   O => msg_block_in_IBUF_348
);
msg_block_in_IBUF_349_inst : IBUF
 port map (
   I => msg_block_in_349,
   O => msg_block_in_IBUF_349
);
msg_block_in_IBUF_34_inst : IBUF
 port map (
   I => msg_block_in_34,
   O => msg_block_in_IBUF_34
);
msg_block_in_IBUF_350_inst : IBUF
 port map (
   I => msg_block_in_350,
   O => msg_block_in_IBUF_350
);
msg_block_in_IBUF_351_inst : IBUF
 port map (
   I => msg_block_in_351,
   O => msg_block_in_IBUF_351
);
msg_block_in_IBUF_352_inst : IBUF
 port map (
   I => msg_block_in_352,
   O => msg_block_in_IBUF_352
);
msg_block_in_IBUF_353_inst : IBUF
 port map (
   I => msg_block_in_353,
   O => msg_block_in_IBUF_353
);
msg_block_in_IBUF_354_inst : IBUF
 port map (
   I => msg_block_in_354,
   O => msg_block_in_IBUF_354
);
msg_block_in_IBUF_355_inst : IBUF
 port map (
   I => msg_block_in_355,
   O => msg_block_in_IBUF_355
);
msg_block_in_IBUF_356_inst : IBUF
 port map (
   I => msg_block_in_356,
   O => msg_block_in_IBUF_356
);
msg_block_in_IBUF_357_inst : IBUF
 port map (
   I => msg_block_in_357,
   O => msg_block_in_IBUF_357
);
msg_block_in_IBUF_358_inst : IBUF
 port map (
   I => msg_block_in_358,
   O => msg_block_in_IBUF_358
);
msg_block_in_IBUF_359_inst : IBUF
 port map (
   I => msg_block_in_359,
   O => msg_block_in_IBUF_359
);
msg_block_in_IBUF_35_inst : IBUF
 port map (
   I => msg_block_in_35,
   O => msg_block_in_IBUF_35
);
msg_block_in_IBUF_360_inst : IBUF
 port map (
   I => msg_block_in_360,
   O => msg_block_in_IBUF_360
);
msg_block_in_IBUF_361_inst : IBUF
 port map (
   I => msg_block_in_361,
   O => msg_block_in_IBUF_361
);
msg_block_in_IBUF_362_inst : IBUF
 port map (
   I => msg_block_in_362,
   O => msg_block_in_IBUF_362
);
msg_block_in_IBUF_363_inst : IBUF
 port map (
   I => msg_block_in_363,
   O => msg_block_in_IBUF_363
);
msg_block_in_IBUF_364_inst : IBUF
 port map (
   I => msg_block_in_364,
   O => msg_block_in_IBUF_364
);
msg_block_in_IBUF_365_inst : IBUF
 port map (
   I => msg_block_in_365,
   O => msg_block_in_IBUF_365
);
msg_block_in_IBUF_366_inst : IBUF
 port map (
   I => msg_block_in_366,
   O => msg_block_in_IBUF_366
);
msg_block_in_IBUF_367_inst : IBUF
 port map (
   I => msg_block_in_367,
   O => msg_block_in_IBUF_367
);
msg_block_in_IBUF_368_inst : IBUF
 port map (
   I => msg_block_in_368,
   O => msg_block_in_IBUF_368
);
msg_block_in_IBUF_369_inst : IBUF
 port map (
   I => msg_block_in_369,
   O => msg_block_in_IBUF_369
);
msg_block_in_IBUF_36_inst : IBUF
 port map (
   I => msg_block_in_36,
   O => msg_block_in_IBUF_36
);
msg_block_in_IBUF_370_inst : IBUF
 port map (
   I => msg_block_in_370,
   O => msg_block_in_IBUF_370
);
msg_block_in_IBUF_371_inst : IBUF
 port map (
   I => msg_block_in_371,
   O => msg_block_in_IBUF_371
);
msg_block_in_IBUF_372_inst : IBUF
 port map (
   I => msg_block_in_372,
   O => msg_block_in_IBUF_372
);
msg_block_in_IBUF_373_inst : IBUF
 port map (
   I => msg_block_in_373,
   O => msg_block_in_IBUF_373
);
msg_block_in_IBUF_374_inst : IBUF
 port map (
   I => msg_block_in_374,
   O => msg_block_in_IBUF_374
);
msg_block_in_IBUF_375_inst : IBUF
 port map (
   I => msg_block_in_375,
   O => msg_block_in_IBUF_375
);
msg_block_in_IBUF_376_inst : IBUF
 port map (
   I => msg_block_in_376,
   O => msg_block_in_IBUF_376
);
msg_block_in_IBUF_377_inst : IBUF
 port map (
   I => msg_block_in_377,
   O => msg_block_in_IBUF_377
);
msg_block_in_IBUF_378_inst : IBUF
 port map (
   I => msg_block_in_378,
   O => msg_block_in_IBUF_378
);
msg_block_in_IBUF_379_inst : IBUF
 port map (
   I => msg_block_in_379,
   O => msg_block_in_IBUF_379
);
msg_block_in_IBUF_37_inst : IBUF
 port map (
   I => msg_block_in_37,
   O => msg_block_in_IBUF_37
);
msg_block_in_IBUF_380_inst : IBUF
 port map (
   I => msg_block_in_380,
   O => msg_block_in_IBUF_380
);
msg_block_in_IBUF_381_inst : IBUF
 port map (
   I => msg_block_in_381,
   O => msg_block_in_IBUF_381
);
msg_block_in_IBUF_382_inst : IBUF
 port map (
   I => msg_block_in_382,
   O => msg_block_in_IBUF_382
);
msg_block_in_IBUF_383_inst : IBUF
 port map (
   I => msg_block_in_383,
   O => msg_block_in_IBUF_383
);
msg_block_in_IBUF_384_inst : IBUF
 port map (
   I => msg_block_in_384,
   O => msg_block_in_IBUF_384
);
msg_block_in_IBUF_385_inst : IBUF
 port map (
   I => msg_block_in_385,
   O => msg_block_in_IBUF_385
);
msg_block_in_IBUF_386_inst : IBUF
 port map (
   I => msg_block_in_386,
   O => msg_block_in_IBUF_386
);
msg_block_in_IBUF_387_inst : IBUF
 port map (
   I => msg_block_in_387,
   O => msg_block_in_IBUF_387
);
msg_block_in_IBUF_388_inst : IBUF
 port map (
   I => msg_block_in_388,
   O => msg_block_in_IBUF_388
);
msg_block_in_IBUF_389_inst : IBUF
 port map (
   I => msg_block_in_389,
   O => msg_block_in_IBUF_389
);
msg_block_in_IBUF_38_inst : IBUF
 port map (
   I => msg_block_in_38,
   O => msg_block_in_IBUF_38
);
msg_block_in_IBUF_390_inst : IBUF
 port map (
   I => msg_block_in_390,
   O => msg_block_in_IBUF_390
);
msg_block_in_IBUF_391_inst : IBUF
 port map (
   I => msg_block_in_391,
   O => msg_block_in_IBUF_391
);
msg_block_in_IBUF_392_inst : IBUF
 port map (
   I => msg_block_in_392,
   O => msg_block_in_IBUF_392
);
msg_block_in_IBUF_393_inst : IBUF
 port map (
   I => msg_block_in_393,
   O => msg_block_in_IBUF_393
);
msg_block_in_IBUF_394_inst : IBUF
 port map (
   I => msg_block_in_394,
   O => msg_block_in_IBUF_394
);
msg_block_in_IBUF_395_inst : IBUF
 port map (
   I => msg_block_in_395,
   O => msg_block_in_IBUF_395
);
msg_block_in_IBUF_396_inst : IBUF
 port map (
   I => msg_block_in_396,
   O => msg_block_in_IBUF_396
);
msg_block_in_IBUF_397_inst : IBUF
 port map (
   I => msg_block_in_397,
   O => msg_block_in_IBUF_397
);
msg_block_in_IBUF_398_inst : IBUF
 port map (
   I => msg_block_in_398,
   O => msg_block_in_IBUF_398
);
msg_block_in_IBUF_399_inst : IBUF
 port map (
   I => msg_block_in_399,
   O => msg_block_in_IBUF_399
);
msg_block_in_IBUF_39_inst : IBUF
 port map (
   I => msg_block_in_39,
   O => msg_block_in_IBUF_39
);
msg_block_in_IBUF_3_inst : IBUF
 port map (
   I => msg_block_in_3,
   O => msg_block_in_IBUF_3
);
msg_block_in_IBUF_400_inst : IBUF
 port map (
   I => msg_block_in_400,
   O => msg_block_in_IBUF_400
);
msg_block_in_IBUF_401_inst : IBUF
 port map (
   I => msg_block_in_401,
   O => msg_block_in_IBUF_401
);
msg_block_in_IBUF_402_inst : IBUF
 port map (
   I => msg_block_in_402,
   O => msg_block_in_IBUF_402
);
msg_block_in_IBUF_403_inst : IBUF
 port map (
   I => msg_block_in_403,
   O => msg_block_in_IBUF_403
);
msg_block_in_IBUF_404_inst : IBUF
 port map (
   I => msg_block_in_404,
   O => msg_block_in_IBUF_404
);
msg_block_in_IBUF_405_inst : IBUF
 port map (
   I => msg_block_in_405,
   O => msg_block_in_IBUF_405
);
msg_block_in_IBUF_406_inst : IBUF
 port map (
   I => msg_block_in_406,
   O => msg_block_in_IBUF_406
);
msg_block_in_IBUF_407_inst : IBUF
 port map (
   I => msg_block_in_407,
   O => msg_block_in_IBUF_407
);
msg_block_in_IBUF_408_inst : IBUF
 port map (
   I => msg_block_in_408,
   O => msg_block_in_IBUF_408
);
msg_block_in_IBUF_409_inst : IBUF
 port map (
   I => msg_block_in_409,
   O => msg_block_in_IBUF_409
);
msg_block_in_IBUF_40_inst : IBUF
 port map (
   I => msg_block_in_40,
   O => msg_block_in_IBUF_40
);
msg_block_in_IBUF_410_inst : IBUF
 port map (
   I => msg_block_in_410,
   O => msg_block_in_IBUF_410
);
msg_block_in_IBUF_411_inst : IBUF
 port map (
   I => msg_block_in_411,
   O => msg_block_in_IBUF_411
);
msg_block_in_IBUF_412_inst : IBUF
 port map (
   I => msg_block_in_412,
   O => msg_block_in_IBUF_412
);
msg_block_in_IBUF_413_inst : IBUF
 port map (
   I => msg_block_in_413,
   O => msg_block_in_IBUF_413
);
msg_block_in_IBUF_414_inst : IBUF
 port map (
   I => msg_block_in_414,
   O => msg_block_in_IBUF_414
);
msg_block_in_IBUF_415_inst : IBUF
 port map (
   I => msg_block_in_415,
   O => msg_block_in_IBUF_415
);
msg_block_in_IBUF_416_inst : IBUF
 port map (
   I => msg_block_in_416,
   O => msg_block_in_IBUF_416
);
msg_block_in_IBUF_417_inst : IBUF
 port map (
   I => msg_block_in_417,
   O => msg_block_in_IBUF_417
);
msg_block_in_IBUF_418_inst : IBUF
 port map (
   I => msg_block_in_418,
   O => msg_block_in_IBUF_418
);
msg_block_in_IBUF_419_inst : IBUF
 port map (
   I => msg_block_in_419,
   O => msg_block_in_IBUF_419
);
msg_block_in_IBUF_41_inst : IBUF
 port map (
   I => msg_block_in_41,
   O => msg_block_in_IBUF_41
);
msg_block_in_IBUF_420_inst : IBUF
 port map (
   I => msg_block_in_420,
   O => msg_block_in_IBUF_420
);
msg_block_in_IBUF_421_inst : IBUF
 port map (
   I => msg_block_in_421,
   O => msg_block_in_IBUF_421
);
msg_block_in_IBUF_422_inst : IBUF
 port map (
   I => msg_block_in_422,
   O => msg_block_in_IBUF_422
);
msg_block_in_IBUF_423_inst : IBUF
 port map (
   I => msg_block_in_423,
   O => msg_block_in_IBUF_423
);
msg_block_in_IBUF_424_inst : IBUF
 port map (
   I => msg_block_in_424,
   O => msg_block_in_IBUF_424
);
msg_block_in_IBUF_425_inst : IBUF
 port map (
   I => msg_block_in_425,
   O => msg_block_in_IBUF_425
);
msg_block_in_IBUF_426_inst : IBUF
 port map (
   I => msg_block_in_426,
   O => msg_block_in_IBUF_426
);
msg_block_in_IBUF_427_inst : IBUF
 port map (
   I => msg_block_in_427,
   O => msg_block_in_IBUF_427
);
msg_block_in_IBUF_428_inst : IBUF
 port map (
   I => msg_block_in_428,
   O => msg_block_in_IBUF_428
);
msg_block_in_IBUF_429_inst : IBUF
 port map (
   I => msg_block_in_429,
   O => msg_block_in_IBUF_429
);
msg_block_in_IBUF_42_inst : IBUF
 port map (
   I => msg_block_in_42,
   O => msg_block_in_IBUF_42
);
msg_block_in_IBUF_430_inst : IBUF
 port map (
   I => msg_block_in_430,
   O => msg_block_in_IBUF_430
);
msg_block_in_IBUF_431_inst : IBUF
 port map (
   I => msg_block_in_431,
   O => msg_block_in_IBUF_431
);
msg_block_in_IBUF_432_inst : IBUF
 port map (
   I => msg_block_in_432,
   O => msg_block_in_IBUF_432
);
msg_block_in_IBUF_433_inst : IBUF
 port map (
   I => msg_block_in_433,
   O => msg_block_in_IBUF_433
);
msg_block_in_IBUF_434_inst : IBUF
 port map (
   I => msg_block_in_434,
   O => msg_block_in_IBUF_434
);
msg_block_in_IBUF_435_inst : IBUF
 port map (
   I => msg_block_in_435,
   O => msg_block_in_IBUF_435
);
msg_block_in_IBUF_436_inst : IBUF
 port map (
   I => msg_block_in_436,
   O => msg_block_in_IBUF_436
);
msg_block_in_IBUF_437_inst : IBUF
 port map (
   I => msg_block_in_437,
   O => msg_block_in_IBUF_437
);
msg_block_in_IBUF_438_inst : IBUF
 port map (
   I => msg_block_in_438,
   O => msg_block_in_IBUF_438
);
msg_block_in_IBUF_439_inst : IBUF
 port map (
   I => msg_block_in_439,
   O => msg_block_in_IBUF_439
);
msg_block_in_IBUF_43_inst : IBUF
 port map (
   I => msg_block_in_43,
   O => msg_block_in_IBUF_43
);
msg_block_in_IBUF_440_inst : IBUF
 port map (
   I => msg_block_in_440,
   O => msg_block_in_IBUF_440
);
msg_block_in_IBUF_441_inst : IBUF
 port map (
   I => msg_block_in_441,
   O => msg_block_in_IBUF_441
);
msg_block_in_IBUF_442_inst : IBUF
 port map (
   I => msg_block_in_442,
   O => msg_block_in_IBUF_442
);
msg_block_in_IBUF_443_inst : IBUF
 port map (
   I => msg_block_in_443,
   O => msg_block_in_IBUF_443
);
msg_block_in_IBUF_444_inst : IBUF
 port map (
   I => msg_block_in_444,
   O => msg_block_in_IBUF_444
);
msg_block_in_IBUF_445_inst : IBUF
 port map (
   I => msg_block_in_445,
   O => msg_block_in_IBUF_445
);
msg_block_in_IBUF_446_inst : IBUF
 port map (
   I => msg_block_in_446,
   O => msg_block_in_IBUF_446
);
msg_block_in_IBUF_447_inst : IBUF
 port map (
   I => msg_block_in_447,
   O => msg_block_in_IBUF_447
);
msg_block_in_IBUF_448_inst : IBUF
 port map (
   I => msg_block_in_448,
   O => msg_block_in_IBUF_448
);
msg_block_in_IBUF_449_inst : IBUF
 port map (
   I => msg_block_in_449,
   O => msg_block_in_IBUF_449
);
msg_block_in_IBUF_44_inst : IBUF
 port map (
   I => msg_block_in_44,
   O => msg_block_in_IBUF_44
);
msg_block_in_IBUF_450_inst : IBUF
 port map (
   I => msg_block_in_450,
   O => msg_block_in_IBUF_450
);
msg_block_in_IBUF_451_inst : IBUF
 port map (
   I => msg_block_in_451,
   O => msg_block_in_IBUF_451
);
msg_block_in_IBUF_452_inst : IBUF
 port map (
   I => msg_block_in_452,
   O => msg_block_in_IBUF_452
);
msg_block_in_IBUF_453_inst : IBUF
 port map (
   I => msg_block_in_453,
   O => msg_block_in_IBUF_453
);
msg_block_in_IBUF_454_inst : IBUF
 port map (
   I => msg_block_in_454,
   O => msg_block_in_IBUF_454
);
msg_block_in_IBUF_455_inst : IBUF
 port map (
   I => msg_block_in_455,
   O => msg_block_in_IBUF_455
);
msg_block_in_IBUF_456_inst : IBUF
 port map (
   I => msg_block_in_456,
   O => msg_block_in_IBUF_456
);
msg_block_in_IBUF_457_inst : IBUF
 port map (
   I => msg_block_in_457,
   O => msg_block_in_IBUF_457
);
msg_block_in_IBUF_458_inst : IBUF
 port map (
   I => msg_block_in_458,
   O => msg_block_in_IBUF_458
);
msg_block_in_IBUF_459_inst : IBUF
 port map (
   I => msg_block_in_459,
   O => msg_block_in_IBUF_459
);
msg_block_in_IBUF_45_inst : IBUF
 port map (
   I => msg_block_in_45,
   O => msg_block_in_IBUF_45
);
msg_block_in_IBUF_460_inst : IBUF
 port map (
   I => msg_block_in_460,
   O => msg_block_in_IBUF_460
);
msg_block_in_IBUF_461_inst : IBUF
 port map (
   I => msg_block_in_461,
   O => msg_block_in_IBUF_461
);
msg_block_in_IBUF_462_inst : IBUF
 port map (
   I => msg_block_in_462,
   O => msg_block_in_IBUF_462
);
msg_block_in_IBUF_463_inst : IBUF
 port map (
   I => msg_block_in_463,
   O => msg_block_in_IBUF_463
);
msg_block_in_IBUF_464_inst : IBUF
 port map (
   I => msg_block_in_464,
   O => msg_block_in_IBUF_464
);
msg_block_in_IBUF_465_inst : IBUF
 port map (
   I => msg_block_in_465,
   O => msg_block_in_IBUF_465
);
msg_block_in_IBUF_466_inst : IBUF
 port map (
   I => msg_block_in_466,
   O => msg_block_in_IBUF_466
);
msg_block_in_IBUF_467_inst : IBUF
 port map (
   I => msg_block_in_467,
   O => msg_block_in_IBUF_467
);
msg_block_in_IBUF_468_inst : IBUF
 port map (
   I => msg_block_in_468,
   O => msg_block_in_IBUF_468
);
msg_block_in_IBUF_469_inst : IBUF
 port map (
   I => msg_block_in_469,
   O => msg_block_in_IBUF_469
);
msg_block_in_IBUF_46_inst : IBUF
 port map (
   I => msg_block_in_46,
   O => msg_block_in_IBUF_46
);
msg_block_in_IBUF_470_inst : IBUF
 port map (
   I => msg_block_in_470,
   O => msg_block_in_IBUF_470
);
msg_block_in_IBUF_471_inst : IBUF
 port map (
   I => msg_block_in_471,
   O => msg_block_in_IBUF_471
);
msg_block_in_IBUF_472_inst : IBUF
 port map (
   I => msg_block_in_472,
   O => msg_block_in_IBUF_472
);
msg_block_in_IBUF_473_inst : IBUF
 port map (
   I => msg_block_in_473,
   O => msg_block_in_IBUF_473
);
msg_block_in_IBUF_474_inst : IBUF
 port map (
   I => msg_block_in_474,
   O => msg_block_in_IBUF_474
);
msg_block_in_IBUF_475_inst : IBUF
 port map (
   I => msg_block_in_475,
   O => msg_block_in_IBUF_475
);
msg_block_in_IBUF_476_inst : IBUF
 port map (
   I => msg_block_in_476,
   O => msg_block_in_IBUF_476
);
msg_block_in_IBUF_477_inst : IBUF
 port map (
   I => msg_block_in_477,
   O => msg_block_in_IBUF_477
);
msg_block_in_IBUF_478_inst : IBUF
 port map (
   I => msg_block_in_478,
   O => msg_block_in_IBUF_478
);
msg_block_in_IBUF_479_inst : IBUF
 port map (
   I => msg_block_in_479,
   O => msg_block_in_IBUF_479
);
msg_block_in_IBUF_47_inst : IBUF
 port map (
   I => msg_block_in_47,
   O => msg_block_in_IBUF_47
);
msg_block_in_IBUF_480_inst : IBUF
 port map (
   I => msg_block_in_480,
   O => msg_block_in_IBUF_480
);
msg_block_in_IBUF_481_inst : IBUF
 port map (
   I => msg_block_in_481,
   O => msg_block_in_IBUF_481
);
msg_block_in_IBUF_482_inst : IBUF
 port map (
   I => msg_block_in_482,
   O => msg_block_in_IBUF_482
);
msg_block_in_IBUF_483_inst : IBUF
 port map (
   I => msg_block_in_483,
   O => msg_block_in_IBUF_483
);
msg_block_in_IBUF_484_inst : IBUF
 port map (
   I => msg_block_in_484,
   O => msg_block_in_IBUF_484
);
msg_block_in_IBUF_485_inst : IBUF
 port map (
   I => msg_block_in_485,
   O => msg_block_in_IBUF_485
);
msg_block_in_IBUF_486_inst : IBUF
 port map (
   I => msg_block_in_486,
   O => msg_block_in_IBUF_486
);
msg_block_in_IBUF_487_inst : IBUF
 port map (
   I => msg_block_in_487,
   O => msg_block_in_IBUF_487
);
msg_block_in_IBUF_488_inst : IBUF
 port map (
   I => msg_block_in_488,
   O => msg_block_in_IBUF_488
);
msg_block_in_IBUF_489_inst : IBUF
 port map (
   I => msg_block_in_489,
   O => msg_block_in_IBUF_489
);
msg_block_in_IBUF_48_inst : IBUF
 port map (
   I => msg_block_in_48,
   O => msg_block_in_IBUF_48
);
msg_block_in_IBUF_490_inst : IBUF
 port map (
   I => msg_block_in_490,
   O => msg_block_in_IBUF_490
);
msg_block_in_IBUF_491_inst : IBUF
 port map (
   I => msg_block_in_491,
   O => msg_block_in_IBUF_491
);
msg_block_in_IBUF_492_inst : IBUF
 port map (
   I => msg_block_in_492,
   O => msg_block_in_IBUF_492
);
msg_block_in_IBUF_493_inst : IBUF
 port map (
   I => msg_block_in_493,
   O => msg_block_in_IBUF_493
);
msg_block_in_IBUF_494_inst : IBUF
 port map (
   I => msg_block_in_494,
   O => msg_block_in_IBUF_494
);
msg_block_in_IBUF_495_inst : IBUF
 port map (
   I => msg_block_in_495,
   O => msg_block_in_IBUF_495
);
msg_block_in_IBUF_496_inst : IBUF
 port map (
   I => msg_block_in_496,
   O => msg_block_in_IBUF_496
);
msg_block_in_IBUF_497_inst : IBUF
 port map (
   I => msg_block_in_497,
   O => msg_block_in_IBUF_497
);
msg_block_in_IBUF_498_inst : IBUF
 port map (
   I => msg_block_in_498,
   O => msg_block_in_IBUF_498
);
msg_block_in_IBUF_499_inst : IBUF
 port map (
   I => msg_block_in_499,
   O => msg_block_in_IBUF_499
);
msg_block_in_IBUF_49_inst : IBUF
 port map (
   I => msg_block_in_49,
   O => msg_block_in_IBUF_49
);
msg_block_in_IBUF_4_inst : IBUF
 port map (
   I => msg_block_in_4,
   O => msg_block_in_IBUF_4
);
msg_block_in_IBUF_500_inst : IBUF
 port map (
   I => msg_block_in_500,
   O => msg_block_in_IBUF_500
);
msg_block_in_IBUF_501_inst : IBUF
 port map (
   I => msg_block_in_501,
   O => msg_block_in_IBUF_501
);
msg_block_in_IBUF_502_inst : IBUF
 port map (
   I => msg_block_in_502,
   O => msg_block_in_IBUF_502
);
msg_block_in_IBUF_503_inst : IBUF
 port map (
   I => msg_block_in_503,
   O => msg_block_in_IBUF_503
);
msg_block_in_IBUF_504_inst : IBUF
 port map (
   I => msg_block_in_504,
   O => msg_block_in_IBUF_504
);
msg_block_in_IBUF_505_inst : IBUF
 port map (
   I => msg_block_in_505,
   O => msg_block_in_IBUF_505
);
msg_block_in_IBUF_506_inst : IBUF
 port map (
   I => msg_block_in_506,
   O => msg_block_in_IBUF_506
);
msg_block_in_IBUF_507_inst : IBUF
 port map (
   I => msg_block_in_507,
   O => msg_block_in_IBUF_507
);
msg_block_in_IBUF_508_inst : IBUF
 port map (
   I => msg_block_in_508,
   O => msg_block_in_IBUF_508
);
msg_block_in_IBUF_509_inst : IBUF
 port map (
   I => msg_block_in_509,
   O => msg_block_in_IBUF_509
);
msg_block_in_IBUF_50_inst : IBUF
 port map (
   I => msg_block_in_50,
   O => msg_block_in_IBUF_50
);
msg_block_in_IBUF_510_inst : IBUF
 port map (
   I => msg_block_in_510,
   O => msg_block_in_IBUF_510
);
msg_block_in_IBUF_511_inst : IBUF
 port map (
   I => msg_block_in_511,
   O => msg_block_in_IBUF_511
);
msg_block_in_IBUF_51_inst : IBUF
 port map (
   I => msg_block_in_51,
   O => msg_block_in_IBUF_51
);
msg_block_in_IBUF_52_inst : IBUF
 port map (
   I => msg_block_in_52,
   O => msg_block_in_IBUF_52
);
msg_block_in_IBUF_53_inst : IBUF
 port map (
   I => msg_block_in_53,
   O => msg_block_in_IBUF_53
);
msg_block_in_IBUF_54_inst : IBUF
 port map (
   I => msg_block_in_54,
   O => msg_block_in_IBUF_54
);
msg_block_in_IBUF_55_inst : IBUF
 port map (
   I => msg_block_in_55,
   O => msg_block_in_IBUF_55
);
msg_block_in_IBUF_56_inst : IBUF
 port map (
   I => msg_block_in_56,
   O => msg_block_in_IBUF_56
);
msg_block_in_IBUF_57_inst : IBUF
 port map (
   I => msg_block_in_57,
   O => msg_block_in_IBUF_57
);
msg_block_in_IBUF_58_inst : IBUF
 port map (
   I => msg_block_in_58,
   O => msg_block_in_IBUF_58
);
msg_block_in_IBUF_59_inst : IBUF
 port map (
   I => msg_block_in_59,
   O => msg_block_in_IBUF_59
);
msg_block_in_IBUF_5_inst : IBUF
 port map (
   I => msg_block_in_5,
   O => msg_block_in_IBUF_5
);
msg_block_in_IBUF_60_inst : IBUF
 port map (
   I => msg_block_in_60,
   O => msg_block_in_IBUF_60
);
msg_block_in_IBUF_61_inst : IBUF
 port map (
   I => msg_block_in_61,
   O => msg_block_in_IBUF_61
);
msg_block_in_IBUF_62_inst : IBUF
 port map (
   I => msg_block_in_62,
   O => msg_block_in_IBUF_62
);
msg_block_in_IBUF_63_inst : IBUF
 port map (
   I => msg_block_in_63,
   O => msg_block_in_IBUF_63
);
msg_block_in_IBUF_64_inst : IBUF
 port map (
   I => msg_block_in_64,
   O => msg_block_in_IBUF_64
);
msg_block_in_IBUF_65_inst : IBUF
 port map (
   I => msg_block_in_65,
   O => msg_block_in_IBUF_65
);
msg_block_in_IBUF_66_inst : IBUF
 port map (
   I => msg_block_in_66,
   O => msg_block_in_IBUF_66
);
msg_block_in_IBUF_67_inst : IBUF
 port map (
   I => msg_block_in_67,
   O => msg_block_in_IBUF_67
);
msg_block_in_IBUF_68_inst : IBUF
 port map (
   I => msg_block_in_68,
   O => msg_block_in_IBUF_68
);
msg_block_in_IBUF_69_inst : IBUF
 port map (
   I => msg_block_in_69,
   O => msg_block_in_IBUF_69
);
msg_block_in_IBUF_6_inst : IBUF
 port map (
   I => msg_block_in_6,
   O => msg_block_in_IBUF_6
);
msg_block_in_IBUF_70_inst : IBUF
 port map (
   I => msg_block_in_70,
   O => msg_block_in_IBUF_70
);
msg_block_in_IBUF_71_inst : IBUF
 port map (
   I => msg_block_in_71,
   O => msg_block_in_IBUF_71
);
msg_block_in_IBUF_72_inst : IBUF
 port map (
   I => msg_block_in_72,
   O => msg_block_in_IBUF_72
);
msg_block_in_IBUF_73_inst : IBUF
 port map (
   I => msg_block_in_73,
   O => msg_block_in_IBUF_73
);
msg_block_in_IBUF_74_inst : IBUF
 port map (
   I => msg_block_in_74,
   O => msg_block_in_IBUF_74
);
msg_block_in_IBUF_75_inst : IBUF
 port map (
   I => msg_block_in_75,
   O => msg_block_in_IBUF_75
);
msg_block_in_IBUF_76_inst : IBUF
 port map (
   I => msg_block_in_76,
   O => msg_block_in_IBUF_76
);
msg_block_in_IBUF_77_inst : IBUF
 port map (
   I => msg_block_in_77,
   O => msg_block_in_IBUF_77
);
msg_block_in_IBUF_78_inst : IBUF
 port map (
   I => msg_block_in_78,
   O => msg_block_in_IBUF_78
);
msg_block_in_IBUF_79_inst : IBUF
 port map (
   I => msg_block_in_79,
   O => msg_block_in_IBUF_79
);
msg_block_in_IBUF_7_inst : IBUF
 port map (
   I => msg_block_in_7,
   O => msg_block_in_IBUF_7
);
msg_block_in_IBUF_80_inst : IBUF
 port map (
   I => msg_block_in_80,
   O => msg_block_in_IBUF_80
);
msg_block_in_IBUF_81_inst : IBUF
 port map (
   I => msg_block_in_81,
   O => msg_block_in_IBUF_81
);
msg_block_in_IBUF_82_inst : IBUF
 port map (
   I => msg_block_in_82,
   O => msg_block_in_IBUF_82
);
msg_block_in_IBUF_83_inst : IBUF
 port map (
   I => msg_block_in_83,
   O => msg_block_in_IBUF_83
);
msg_block_in_IBUF_84_inst : IBUF
 port map (
   I => msg_block_in_84,
   O => msg_block_in_IBUF_84
);
msg_block_in_IBUF_85_inst : IBUF
 port map (
   I => msg_block_in_85,
   O => msg_block_in_IBUF_85
);
msg_block_in_IBUF_86_inst : IBUF
 port map (
   I => msg_block_in_86,
   O => msg_block_in_IBUF_86
);
msg_block_in_IBUF_87_inst : IBUF
 port map (
   I => msg_block_in_87,
   O => msg_block_in_IBUF_87
);
msg_block_in_IBUF_88_inst : IBUF
 port map (
   I => msg_block_in_88,
   O => msg_block_in_IBUF_88
);
msg_block_in_IBUF_89_inst : IBUF
 port map (
   I => msg_block_in_89,
   O => msg_block_in_IBUF_89
);
msg_block_in_IBUF_8_inst : IBUF
 port map (
   I => msg_block_in_8,
   O => msg_block_in_IBUF_8
);
msg_block_in_IBUF_90_inst : IBUF
 port map (
   I => msg_block_in_90,
   O => msg_block_in_IBUF_90
);
msg_block_in_IBUF_91_inst : IBUF
 port map (
   I => msg_block_in_91,
   O => msg_block_in_IBUF_91
);
msg_block_in_IBUF_92_inst : IBUF
 port map (
   I => msg_block_in_92,
   O => msg_block_in_IBUF_92
);
msg_block_in_IBUF_93_inst : IBUF
 port map (
   I => msg_block_in_93,
   O => msg_block_in_IBUF_93
);
msg_block_in_IBUF_94_inst : IBUF
 port map (
   I => msg_block_in_94,
   O => msg_block_in_IBUF_94
);
msg_block_in_IBUF_95_inst : IBUF
 port map (
   I => msg_block_in_95,
   O => msg_block_in_IBUF_95
);
msg_block_in_IBUF_96_inst : IBUF
 port map (
   I => msg_block_in_96,
   O => msg_block_in_IBUF_96
);
msg_block_in_IBUF_97_inst : IBUF
 port map (
   I => msg_block_in_97,
   O => msg_block_in_IBUF_97
);
msg_block_in_IBUF_98_inst : IBUF
 port map (
   I => msg_block_in_98,
   O => msg_block_in_IBUF_98
);
msg_block_in_IBUF_99_inst : IBUF
 port map (
   I => msg_block_in_99,
   O => msg_block_in_IBUF_99
);
msg_block_in_IBUF_9_inst : IBUF
 port map (
   I => msg_block_in_9,
   O => msg_block_in_IBUF_9
);
M_0_31_i_1 : LUT2
  generic map(
   INIT => X"2"
  )
 port map (
   I0 => M_0,
   I1 => rst_IBUF,
   O => M_reg_0_0
);
M_reg_0_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_31,
   R => '0',
   Q => M_reg_0_0
);
M_reg_0_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_21,
   R => '0',
   Q => M_reg_0_10
);
M_reg_0_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_20,
   R => '0',
   Q => M_reg_0_11
);
M_reg_0_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_19,
   R => '0',
   Q => M_reg_0_12
);
M_reg_0_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_18,
   R => '0',
   Q => M_reg_0_13
);
M_reg_0_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_17,
   R => '0',
   Q => M_reg_0_14
);
M_reg_0_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_16,
   R => '0',
   Q => M_reg_0_15
);
M_reg_0_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_15,
   R => '0',
   Q => M_reg_0_16
);
M_reg_0_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_14,
   R => '0',
   Q => M_reg_0_17
);
M_reg_0_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_13,
   R => '0',
   Q => M_reg_0_18
);
M_reg_0_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_12,
   R => '0',
   Q => M_reg_0_19
);
M_reg_0_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_30,
   R => '0',
   Q => M_reg_0_1
);
M_reg_0_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_11,
   R => '0',
   Q => M_reg_0_20
);
M_reg_0_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_10,
   R => '0',
   Q => M_reg_0_21
);
M_reg_0_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_9,
   R => '0',
   Q => M_reg_0_22
);
M_reg_0_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_8,
   R => '0',
   Q => M_reg_0_23
);
M_reg_0_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_7,
   R => '0',
   Q => M_reg_0_24
);
M_reg_0_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_6,
   R => '0',
   Q => M_reg_0_25
);
M_reg_0_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_5,
   R => '0',
   Q => M_reg_0_26
);
M_reg_0_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_4,
   R => '0',
   Q => M_reg_0_27
);
M_reg_0_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_3,
   R => '0',
   Q => M_reg_0_28
);
M_reg_0_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_2,
   R => '0',
   Q => M_reg_0_29
);
M_reg_0_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_29,
   R => '0',
   Q => M_reg_0_2
);
M_reg_0_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_1,
   R => '0',
   Q => M_reg_0_30
);
M_reg_0_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_0,
   R => '0',
   Q => M_reg_0_31
);
M_reg_0_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_28,
   R => '0',
   Q => M_reg_0_3
);
M_reg_0_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_27,
   R => '0',
   Q => M_reg_0_4
);
M_reg_0_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_26,
   R => '0',
   Q => M_reg_0_5
);
M_reg_0_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_25,
   R => '0',
   Q => M_reg_0_6
);
M_reg_0_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_24,
   R => '0',
   Q => M_reg_0_7
);
M_reg_0_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_23,
   R => '0',
   Q => M_reg_0_8
);
M_reg_0_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_22,
   R => '0',
   Q => M_reg_0_9
);
M_reg_10_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_351,
   R => '0',
   Q => M_reg_10_0
);
M_reg_10_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_341,
   R => '0',
   Q => M_reg_10_10
);
M_reg_10_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_340,
   R => '0',
   Q => M_reg_10_11
);
M_reg_10_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_339,
   R => '0',
   Q => M_reg_10_12
);
M_reg_10_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_338,
   R => '0',
   Q => M_reg_10_13
);
M_reg_10_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_337,
   R => '0',
   Q => M_reg_10_14
);
M_reg_10_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_336,
   R => '0',
   Q => M_reg_10_15
);
M_reg_10_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_335,
   R => '0',
   Q => M_reg_10_16
);
M_reg_10_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_334,
   R => '0',
   Q => M_reg_10_17
);
M_reg_10_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_333,
   R => '0',
   Q => M_reg_10_18
);
M_reg_10_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_332,
   R => '0',
   Q => M_reg_10_19
);
M_reg_10_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_350,
   R => '0',
   Q => M_reg_10_1
);
M_reg_10_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_331,
   R => '0',
   Q => M_reg_10_20
);
M_reg_10_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_330,
   R => '0',
   Q => M_reg_10_21
);
M_reg_10_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_329,
   R => '0',
   Q => M_reg_10_22
);
M_reg_10_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_328,
   R => '0',
   Q => M_reg_10_23
);
M_reg_10_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_327,
   R => '0',
   Q => M_reg_10_24
);
M_reg_10_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_326,
   R => '0',
   Q => M_reg_10_25
);
M_reg_10_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_325,
   R => '0',
   Q => M_reg_10_26
);
M_reg_10_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_324,
   R => '0',
   Q => M_reg_10_27
);
M_reg_10_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_323,
   R => '0',
   Q => M_reg_10_28
);
M_reg_10_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_322,
   R => '0',
   Q => M_reg_10_29
);
M_reg_10_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_349,
   R => '0',
   Q => M_reg_10_2
);
M_reg_10_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_321,
   R => '0',
   Q => M_reg_10_30
);
M_reg_10_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_320,
   R => '0',
   Q => M_reg_10_31
);
M_reg_10_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_348,
   R => '0',
   Q => M_reg_10_3
);
M_reg_10_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_347,
   R => '0',
   Q => M_reg_10_4
);
M_reg_10_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_346,
   R => '0',
   Q => M_reg_10_5
);
M_reg_10_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_345,
   R => '0',
   Q => M_reg_10_6
);
M_reg_10_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_344,
   R => '0',
   Q => M_reg_10_7
);
M_reg_10_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_343,
   R => '0',
   Q => M_reg_10_8
);
M_reg_10_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_342,
   R => '0',
   Q => M_reg_10_9
);
M_reg_11_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_383,
   R => '0',
   Q => M_reg_11_0
);
M_reg_11_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_373,
   R => '0',
   Q => M_reg_11_10
);
M_reg_11_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_372,
   R => '0',
   Q => M_reg_11_11
);
M_reg_11_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_371,
   R => '0',
   Q => M_reg_11_12
);
M_reg_11_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_370,
   R => '0',
   Q => M_reg_11_13
);
M_reg_11_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_369,
   R => '0',
   Q => M_reg_11_14
);
M_reg_11_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_368,
   R => '0',
   Q => M_reg_11_15
);
M_reg_11_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_367,
   R => '0',
   Q => M_reg_11_16
);
M_reg_11_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_366,
   R => '0',
   Q => M_reg_11_17
);
M_reg_11_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_365,
   R => '0',
   Q => M_reg_11_18
);
M_reg_11_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_364,
   R => '0',
   Q => M_reg_11_19
);
M_reg_11_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_382,
   R => '0',
   Q => M_reg_11_1
);
M_reg_11_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_363,
   R => '0',
   Q => M_reg_11_20
);
M_reg_11_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_362,
   R => '0',
   Q => M_reg_11_21
);
M_reg_11_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_361,
   R => '0',
   Q => M_reg_11_22
);
M_reg_11_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_360,
   R => '0',
   Q => M_reg_11_23
);
M_reg_11_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_359,
   R => '0',
   Q => M_reg_11_24
);
M_reg_11_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_358,
   R => '0',
   Q => M_reg_11_25
);
M_reg_11_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_357,
   R => '0',
   Q => M_reg_11_26
);
M_reg_11_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_356,
   R => '0',
   Q => M_reg_11_27
);
M_reg_11_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_355,
   R => '0',
   Q => M_reg_11_28
);
M_reg_11_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_354,
   R => '0',
   Q => M_reg_11_29
);
M_reg_11_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_381,
   R => '0',
   Q => M_reg_11_2
);
M_reg_11_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_353,
   R => '0',
   Q => M_reg_11_30
);
M_reg_11_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_352,
   R => '0',
   Q => M_reg_11_31
);
M_reg_11_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_380,
   R => '0',
   Q => M_reg_11_3
);
M_reg_11_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_379,
   R => '0',
   Q => M_reg_11_4
);
M_reg_11_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_378,
   R => '0',
   Q => M_reg_11_5
);
M_reg_11_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_377,
   R => '0',
   Q => M_reg_11_6
);
M_reg_11_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_376,
   R => '0',
   Q => M_reg_11_7
);
M_reg_11_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_375,
   R => '0',
   Q => M_reg_11_8
);
M_reg_11_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_374,
   R => '0',
   Q => M_reg_11_9
);
M_reg_12_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_415,
   R => '0',
   Q => M_reg_12_0
);
M_reg_12_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_405,
   R => '0',
   Q => M_reg_12_10
);
M_reg_12_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_404,
   R => '0',
   Q => M_reg_12_11
);
M_reg_12_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_403,
   R => '0',
   Q => M_reg_12_12
);
M_reg_12_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_402,
   R => '0',
   Q => M_reg_12_13
);
M_reg_12_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_401,
   R => '0',
   Q => M_reg_12_14
);
M_reg_12_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_400,
   R => '0',
   Q => M_reg_12_15
);
M_reg_12_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_399,
   R => '0',
   Q => M_reg_12_16
);
M_reg_12_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_398,
   R => '0',
   Q => M_reg_12_17
);
M_reg_12_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_397,
   R => '0',
   Q => M_reg_12_18
);
M_reg_12_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_396,
   R => '0',
   Q => M_reg_12_19
);
M_reg_12_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_414,
   R => '0',
   Q => M_reg_12_1
);
M_reg_12_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_395,
   R => '0',
   Q => M_reg_12_20
);
M_reg_12_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_394,
   R => '0',
   Q => M_reg_12_21
);
M_reg_12_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_393,
   R => '0',
   Q => M_reg_12_22
);
M_reg_12_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_392,
   R => '0',
   Q => M_reg_12_23
);
M_reg_12_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_391,
   R => '0',
   Q => M_reg_12_24
);
M_reg_12_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_390,
   R => '0',
   Q => M_reg_12_25
);
M_reg_12_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_389,
   R => '0',
   Q => M_reg_12_26
);
M_reg_12_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_388,
   R => '0',
   Q => M_reg_12_27
);
M_reg_12_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_387,
   R => '0',
   Q => M_reg_12_28
);
M_reg_12_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_386,
   R => '0',
   Q => M_reg_12_29
);
M_reg_12_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_413,
   R => '0',
   Q => M_reg_12_2
);
M_reg_12_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_385,
   R => '0',
   Q => M_reg_12_30
);
M_reg_12_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_384,
   R => '0',
   Q => M_reg_12_31
);
M_reg_12_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_412,
   R => '0',
   Q => M_reg_12_3
);
M_reg_12_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_411,
   R => '0',
   Q => M_reg_12_4
);
M_reg_12_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_410,
   R => '0',
   Q => M_reg_12_5
);
M_reg_12_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_409,
   R => '0',
   Q => M_reg_12_6
);
M_reg_12_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_408,
   R => '0',
   Q => M_reg_12_7
);
M_reg_12_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_407,
   R => '0',
   Q => M_reg_12_8
);
M_reg_12_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_406,
   R => '0',
   Q => M_reg_12_9
);
M_reg_13_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_447,
   R => '0',
   Q => M_reg_13_0
);
M_reg_13_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_437,
   R => '0',
   Q => M_reg_13_10
);
M_reg_13_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_436,
   R => '0',
   Q => M_reg_13_11
);
M_reg_13_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_435,
   R => '0',
   Q => M_reg_13_12
);
M_reg_13_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_434,
   R => '0',
   Q => M_reg_13_13
);
M_reg_13_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_433,
   R => '0',
   Q => M_reg_13_14
);
M_reg_13_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_432,
   R => '0',
   Q => M_reg_13_15
);
M_reg_13_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_431,
   R => '0',
   Q => M_reg_13_16
);
M_reg_13_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_430,
   R => '0',
   Q => M_reg_13_17
);
M_reg_13_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_429,
   R => '0',
   Q => M_reg_13_18
);
M_reg_13_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_428,
   R => '0',
   Q => M_reg_13_19
);
M_reg_13_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_446,
   R => '0',
   Q => M_reg_13_1
);
M_reg_13_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_427,
   R => '0',
   Q => M_reg_13_20
);
M_reg_13_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_426,
   R => '0',
   Q => M_reg_13_21
);
M_reg_13_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_425,
   R => '0',
   Q => M_reg_13_22
);
M_reg_13_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_424,
   R => '0',
   Q => M_reg_13_23
);
M_reg_13_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_423,
   R => '0',
   Q => M_reg_13_24
);
M_reg_13_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_422,
   R => '0',
   Q => M_reg_13_25
);
M_reg_13_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_421,
   R => '0',
   Q => M_reg_13_26
);
M_reg_13_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_420,
   R => '0',
   Q => M_reg_13_27
);
M_reg_13_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_419,
   R => '0',
   Q => M_reg_13_28
);
M_reg_13_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_418,
   R => '0',
   Q => M_reg_13_29
);
M_reg_13_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_445,
   R => '0',
   Q => M_reg_13_2
);
M_reg_13_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_417,
   R => '0',
   Q => M_reg_13_30
);
M_reg_13_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_416,
   R => '0',
   Q => M_reg_13_31
);
M_reg_13_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_444,
   R => '0',
   Q => M_reg_13_3
);
M_reg_13_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_443,
   R => '0',
   Q => M_reg_13_4
);
M_reg_13_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_442,
   R => '0',
   Q => M_reg_13_5
);
M_reg_13_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_441,
   R => '0',
   Q => M_reg_13_6
);
M_reg_13_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_440,
   R => '0',
   Q => M_reg_13_7
);
M_reg_13_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_439,
   R => '0',
   Q => M_reg_13_8
);
M_reg_13_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_438,
   R => '0',
   Q => M_reg_13_9
);
M_reg_14_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_479,
   R => '0',
   Q => M_reg_14_0
);
M_reg_14_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_469,
   R => '0',
   Q => M_reg_14_10
);
M_reg_14_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_468,
   R => '0',
   Q => M_reg_14_11
);
M_reg_14_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_467,
   R => '0',
   Q => M_reg_14_12
);
M_reg_14_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_466,
   R => '0',
   Q => M_reg_14_13
);
M_reg_14_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_465,
   R => '0',
   Q => M_reg_14_14
);
M_reg_14_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_464,
   R => '0',
   Q => M_reg_14_15
);
M_reg_14_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_463,
   R => '0',
   Q => M_reg_14_16
);
M_reg_14_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_462,
   R => '0',
   Q => M_reg_14_17
);
M_reg_14_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_461,
   R => '0',
   Q => M_reg_14_18
);
M_reg_14_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_460,
   R => '0',
   Q => M_reg_14_19
);
M_reg_14_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_478,
   R => '0',
   Q => M_reg_14_1
);
M_reg_14_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_459,
   R => '0',
   Q => M_reg_14_20
);
M_reg_14_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_458,
   R => '0',
   Q => M_reg_14_21
);
M_reg_14_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_457,
   R => '0',
   Q => M_reg_14_22
);
M_reg_14_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_456,
   R => '0',
   Q => M_reg_14_23
);
M_reg_14_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_455,
   R => '0',
   Q => M_reg_14_24
);
M_reg_14_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_454,
   R => '0',
   Q => M_reg_14_25
);
M_reg_14_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_453,
   R => '0',
   Q => M_reg_14_26
);
M_reg_14_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_452,
   R => '0',
   Q => M_reg_14_27
);
M_reg_14_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_451,
   R => '0',
   Q => M_reg_14_28
);
M_reg_14_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_450,
   R => '0',
   Q => M_reg_14_29
);
M_reg_14_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_477,
   R => '0',
   Q => M_reg_14_2
);
M_reg_14_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_449,
   R => '0',
   Q => M_reg_14_30
);
M_reg_14_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_448,
   R => '0',
   Q => M_reg_14_31
);
M_reg_14_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_476,
   R => '0',
   Q => M_reg_14_3
);
M_reg_14_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_475,
   R => '0',
   Q => M_reg_14_4
);
M_reg_14_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_474,
   R => '0',
   Q => M_reg_14_5
);
M_reg_14_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_473,
   R => '0',
   Q => M_reg_14_6
);
M_reg_14_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_472,
   R => '0',
   Q => M_reg_14_7
);
M_reg_14_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_471,
   R => '0',
   Q => M_reg_14_8
);
M_reg_14_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_470,
   R => '0',
   Q => M_reg_14_9
);
M_reg_15_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_511,
   R => '0',
   Q => M_reg_15_0
);
M_reg_15_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_501,
   R => '0',
   Q => M_reg_15_10
);
M_reg_15_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_500,
   R => '0',
   Q => M_reg_15_11
);
M_reg_15_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_499,
   R => '0',
   Q => M_reg_15_12
);
M_reg_15_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_498,
   R => '0',
   Q => M_reg_15_13
);
M_reg_15_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_497,
   R => '0',
   Q => M_reg_15_14
);
M_reg_15_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_496,
   R => '0',
   Q => M_reg_15_15
);
M_reg_15_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_495,
   R => '0',
   Q => M_reg_15_16
);
M_reg_15_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_494,
   R => '0',
   Q => M_reg_15_17
);
M_reg_15_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_493,
   R => '0',
   Q => M_reg_15_18
);
M_reg_15_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_492,
   R => '0',
   Q => M_reg_15_19
);
M_reg_15_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_510,
   R => '0',
   Q => M_reg_15_1
);
M_reg_15_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_491,
   R => '0',
   Q => M_reg_15_20
);
M_reg_15_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_490,
   R => '0',
   Q => M_reg_15_21
);
M_reg_15_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_489,
   R => '0',
   Q => M_reg_15_22
);
M_reg_15_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_488,
   R => '0',
   Q => M_reg_15_23
);
M_reg_15_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_487,
   R => '0',
   Q => M_reg_15_24
);
M_reg_15_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_486,
   R => '0',
   Q => M_reg_15_25
);
M_reg_15_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_485,
   R => '0',
   Q => M_reg_15_26
);
M_reg_15_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_484,
   R => '0',
   Q => M_reg_15_27
);
M_reg_15_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_483,
   R => '0',
   Q => M_reg_15_28
);
M_reg_15_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_482,
   R => '0',
   Q => M_reg_15_29
);
M_reg_15_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_509,
   R => '0',
   Q => M_reg_15_2
);
M_reg_15_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_481,
   R => '0',
   Q => M_reg_15_30
);
M_reg_15_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_480,
   R => '0',
   Q => M_reg_15_31
);
M_reg_15_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_508,
   R => '0',
   Q => M_reg_15_3
);
M_reg_15_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_507,
   R => '0',
   Q => M_reg_15_4
);
M_reg_15_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_506,
   R => '0',
   Q => M_reg_15_5
);
M_reg_15_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_505,
   R => '0',
   Q => M_reg_15_6
);
M_reg_15_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_504,
   R => '0',
   Q => M_reg_15_7
);
M_reg_15_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_503,
   R => '0',
   Q => M_reg_15_8
);
M_reg_15_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_502,
   R => '0',
   Q => M_reg_15_9
);
M_reg_1_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_63,
   R => '0',
   Q => M_reg_1_0
);
M_reg_1_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_53,
   R => '0',
   Q => M_reg_1_10
);
M_reg_1_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_52,
   R => '0',
   Q => M_reg_1_11
);
M_reg_1_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_51,
   R => '0',
   Q => M_reg_1_12
);
M_reg_1_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_50,
   R => '0',
   Q => M_reg_1_13
);
M_reg_1_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_49,
   R => '0',
   Q => M_reg_1_14
);
M_reg_1_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_48,
   R => '0',
   Q => M_reg_1_15
);
M_reg_1_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_47,
   R => '0',
   Q => M_reg_1_16
);
M_reg_1_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_46,
   R => '0',
   Q => M_reg_1_17
);
M_reg_1_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_45,
   R => '0',
   Q => M_reg_1_18
);
M_reg_1_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_44,
   R => '0',
   Q => M_reg_1_19
);
M_reg_1_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_62,
   R => '0',
   Q => M_reg_1_1
);
M_reg_1_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_43,
   R => '0',
   Q => M_reg_1_20
);
M_reg_1_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_42,
   R => '0',
   Q => M_reg_1_21
);
M_reg_1_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_41,
   R => '0',
   Q => M_reg_1_22
);
M_reg_1_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_40,
   R => '0',
   Q => M_reg_1_23
);
M_reg_1_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_39,
   R => '0',
   Q => M_reg_1_24
);
M_reg_1_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_38,
   R => '0',
   Q => M_reg_1_25
);
M_reg_1_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_37,
   R => '0',
   Q => M_reg_1_26
);
M_reg_1_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_36,
   R => '0',
   Q => M_reg_1_27
);
M_reg_1_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_35,
   R => '0',
   Q => M_reg_1_28
);
M_reg_1_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_34,
   R => '0',
   Q => M_reg_1_29
);
M_reg_1_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_61,
   R => '0',
   Q => M_reg_1_2
);
M_reg_1_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_33,
   R => '0',
   Q => M_reg_1_30
);
M_reg_1_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_32,
   R => '0',
   Q => M_reg_1_31
);
M_reg_1_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_60,
   R => '0',
   Q => M_reg_1_3
);
M_reg_1_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_59,
   R => '0',
   Q => M_reg_1_4
);
M_reg_1_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_58,
   R => '0',
   Q => M_reg_1_5
);
M_reg_1_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_57,
   R => '0',
   Q => M_reg_1_6
);
M_reg_1_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_56,
   R => '0',
   Q => M_reg_1_7
);
M_reg_1_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_55,
   R => '0',
   Q => M_reg_1_8
);
M_reg_1_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_54,
   R => '0',
   Q => M_reg_1_9
);
M_reg_2_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_95,
   R => '0',
   Q => M_reg_2_0
);
M_reg_2_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_85,
   R => '0',
   Q => M_reg_2_10
);
M_reg_2_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_84,
   R => '0',
   Q => M_reg_2_11
);
M_reg_2_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_83,
   R => '0',
   Q => M_reg_2_12
);
M_reg_2_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_82,
   R => '0',
   Q => M_reg_2_13
);
M_reg_2_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_81,
   R => '0',
   Q => M_reg_2_14
);
M_reg_2_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_80,
   R => '0',
   Q => M_reg_2_15
);
M_reg_2_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_79,
   R => '0',
   Q => M_reg_2_16
);
M_reg_2_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_78,
   R => '0',
   Q => M_reg_2_17
);
M_reg_2_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_77,
   R => '0',
   Q => M_reg_2_18
);
M_reg_2_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_76,
   R => '0',
   Q => M_reg_2_19
);
M_reg_2_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_94,
   R => '0',
   Q => M_reg_2_1
);
M_reg_2_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_75,
   R => '0',
   Q => M_reg_2_20
);
M_reg_2_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_74,
   R => '0',
   Q => M_reg_2_21
);
M_reg_2_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_73,
   R => '0',
   Q => M_reg_2_22
);
M_reg_2_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_72,
   R => '0',
   Q => M_reg_2_23
);
M_reg_2_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_71,
   R => '0',
   Q => M_reg_2_24
);
M_reg_2_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_70,
   R => '0',
   Q => M_reg_2_25
);
M_reg_2_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_69,
   R => '0',
   Q => M_reg_2_26
);
M_reg_2_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_68,
   R => '0',
   Q => M_reg_2_27
);
M_reg_2_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_67,
   R => '0',
   Q => M_reg_2_28
);
M_reg_2_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_66,
   R => '0',
   Q => M_reg_2_29
);
M_reg_2_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_93,
   R => '0',
   Q => M_reg_2_2
);
M_reg_2_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_65,
   R => '0',
   Q => M_reg_2_30
);
M_reg_2_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_64,
   R => '0',
   Q => M_reg_2_31
);
M_reg_2_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_92,
   R => '0',
   Q => M_reg_2_3
);
M_reg_2_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_91,
   R => '0',
   Q => M_reg_2_4
);
M_reg_2_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_90,
   R => '0',
   Q => M_reg_2_5
);
M_reg_2_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_89,
   R => '0',
   Q => M_reg_2_6
);
M_reg_2_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_88,
   R => '0',
   Q => M_reg_2_7
);
M_reg_2_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_87,
   R => '0',
   Q => M_reg_2_8
);
M_reg_2_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_86,
   R => '0',
   Q => M_reg_2_9
);
M_reg_3_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_127,
   R => '0',
   Q => M_reg_3_0
);
M_reg_3_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_117,
   R => '0',
   Q => M_reg_3_10
);
M_reg_3_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_116,
   R => '0',
   Q => M_reg_3_11
);
M_reg_3_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_115,
   R => '0',
   Q => M_reg_3_12
);
M_reg_3_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_114,
   R => '0',
   Q => M_reg_3_13
);
M_reg_3_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_113,
   R => '0',
   Q => M_reg_3_14
);
M_reg_3_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_112,
   R => '0',
   Q => M_reg_3_15
);
M_reg_3_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_111,
   R => '0',
   Q => M_reg_3_16
);
M_reg_3_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_110,
   R => '0',
   Q => M_reg_3_17
);
M_reg_3_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_109,
   R => '0',
   Q => M_reg_3_18
);
M_reg_3_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_108,
   R => '0',
   Q => M_reg_3_19
);
M_reg_3_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_126,
   R => '0',
   Q => M_reg_3_1
);
M_reg_3_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_107,
   R => '0',
   Q => M_reg_3_20
);
M_reg_3_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_106,
   R => '0',
   Q => M_reg_3_21
);
M_reg_3_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_105,
   R => '0',
   Q => M_reg_3_22
);
M_reg_3_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_104,
   R => '0',
   Q => M_reg_3_23
);
M_reg_3_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_103,
   R => '0',
   Q => M_reg_3_24
);
M_reg_3_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_102,
   R => '0',
   Q => M_reg_3_25
);
M_reg_3_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_101,
   R => '0',
   Q => M_reg_3_26
);
M_reg_3_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_100,
   R => '0',
   Q => M_reg_3_27
);
M_reg_3_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_99,
   R => '0',
   Q => M_reg_3_28
);
M_reg_3_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_98,
   R => '0',
   Q => M_reg_3_29
);
M_reg_3_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_125,
   R => '0',
   Q => M_reg_3_2
);
M_reg_3_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_97,
   R => '0',
   Q => M_reg_3_30
);
M_reg_3_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_96,
   R => '0',
   Q => M_reg_3_31
);
M_reg_3_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_124,
   R => '0',
   Q => M_reg_3_3
);
M_reg_3_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_123,
   R => '0',
   Q => M_reg_3_4
);
M_reg_3_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_122,
   R => '0',
   Q => M_reg_3_5
);
M_reg_3_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_121,
   R => '0',
   Q => M_reg_3_6
);
M_reg_3_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_120,
   R => '0',
   Q => M_reg_3_7
);
M_reg_3_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_119,
   R => '0',
   Q => M_reg_3_8
);
M_reg_3_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_118,
   R => '0',
   Q => M_reg_3_9
);
M_reg_4_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_159,
   R => '0',
   Q => M_reg_4_0
);
M_reg_4_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_149,
   R => '0',
   Q => M_reg_4_10
);
M_reg_4_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_148,
   R => '0',
   Q => M_reg_4_11
);
M_reg_4_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_147,
   R => '0',
   Q => M_reg_4_12
);
M_reg_4_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_146,
   R => '0',
   Q => M_reg_4_13
);
M_reg_4_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_145,
   R => '0',
   Q => M_reg_4_14
);
M_reg_4_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_144,
   R => '0',
   Q => M_reg_4_15
);
M_reg_4_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_143,
   R => '0',
   Q => M_reg_4_16
);
M_reg_4_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_142,
   R => '0',
   Q => M_reg_4_17
);
M_reg_4_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_141,
   R => '0',
   Q => M_reg_4_18
);
M_reg_4_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_140,
   R => '0',
   Q => M_reg_4_19
);
M_reg_4_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_158,
   R => '0',
   Q => M_reg_4_1
);
M_reg_4_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_139,
   R => '0',
   Q => M_reg_4_20
);
M_reg_4_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_138,
   R => '0',
   Q => M_reg_4_21
);
M_reg_4_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_137,
   R => '0',
   Q => M_reg_4_22
);
M_reg_4_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_136,
   R => '0',
   Q => M_reg_4_23
);
M_reg_4_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_135,
   R => '0',
   Q => M_reg_4_24
);
M_reg_4_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_134,
   R => '0',
   Q => M_reg_4_25
);
M_reg_4_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_133,
   R => '0',
   Q => M_reg_4_26
);
M_reg_4_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_132,
   R => '0',
   Q => M_reg_4_27
);
M_reg_4_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_131,
   R => '0',
   Q => M_reg_4_28
);
M_reg_4_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_130,
   R => '0',
   Q => M_reg_4_29
);
M_reg_4_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_157,
   R => '0',
   Q => M_reg_4_2
);
M_reg_4_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_129,
   R => '0',
   Q => M_reg_4_30
);
M_reg_4_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_128,
   R => '0',
   Q => M_reg_4_31
);
M_reg_4_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_156,
   R => '0',
   Q => M_reg_4_3
);
M_reg_4_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_155,
   R => '0',
   Q => M_reg_4_4
);
M_reg_4_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_154,
   R => '0',
   Q => M_reg_4_5
);
M_reg_4_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_153,
   R => '0',
   Q => M_reg_4_6
);
M_reg_4_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_152,
   R => '0',
   Q => M_reg_4_7
);
M_reg_4_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_151,
   R => '0',
   Q => M_reg_4_8
);
M_reg_4_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_150,
   R => '0',
   Q => M_reg_4_9
);
M_reg_5_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_191,
   R => '0',
   Q => M_reg_5_0
);
M_reg_5_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_181,
   R => '0',
   Q => M_reg_5_10
);
M_reg_5_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_180,
   R => '0',
   Q => M_reg_5_11
);
M_reg_5_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_179,
   R => '0',
   Q => M_reg_5_12
);
M_reg_5_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_178,
   R => '0',
   Q => M_reg_5_13
);
M_reg_5_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_177,
   R => '0',
   Q => M_reg_5_14
);
M_reg_5_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_176,
   R => '0',
   Q => M_reg_5_15
);
M_reg_5_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_175,
   R => '0',
   Q => M_reg_5_16
);
M_reg_5_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_174,
   R => '0',
   Q => M_reg_5_17
);
M_reg_5_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_173,
   R => '0',
   Q => M_reg_5_18
);
M_reg_5_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_172,
   R => '0',
   Q => M_reg_5_19
);
M_reg_5_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_190,
   R => '0',
   Q => M_reg_5_1
);
M_reg_5_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_171,
   R => '0',
   Q => M_reg_5_20
);
M_reg_5_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_170,
   R => '0',
   Q => M_reg_5_21
);
M_reg_5_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_169,
   R => '0',
   Q => M_reg_5_22
);
M_reg_5_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_168,
   R => '0',
   Q => M_reg_5_23
);
M_reg_5_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_167,
   R => '0',
   Q => M_reg_5_24
);
M_reg_5_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_166,
   R => '0',
   Q => M_reg_5_25
);
M_reg_5_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_165,
   R => '0',
   Q => M_reg_5_26
);
M_reg_5_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_164,
   R => '0',
   Q => M_reg_5_27
);
M_reg_5_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_163,
   R => '0',
   Q => M_reg_5_28
);
M_reg_5_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_162,
   R => '0',
   Q => M_reg_5_29
);
M_reg_5_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_189,
   R => '0',
   Q => M_reg_5_2
);
M_reg_5_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_161,
   R => '0',
   Q => M_reg_5_30
);
M_reg_5_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_160,
   R => '0',
   Q => M_reg_5_31
);
M_reg_5_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_188,
   R => '0',
   Q => M_reg_5_3
);
M_reg_5_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_187,
   R => '0',
   Q => M_reg_5_4
);
M_reg_5_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_186,
   R => '0',
   Q => M_reg_5_5
);
M_reg_5_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_185,
   R => '0',
   Q => M_reg_5_6
);
M_reg_5_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_184,
   R => '0',
   Q => M_reg_5_7
);
M_reg_5_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_183,
   R => '0',
   Q => M_reg_5_8
);
M_reg_5_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_182,
   R => '0',
   Q => M_reg_5_9
);
M_reg_6_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_223,
   R => '0',
   Q => M_reg_6_0
);
M_reg_6_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_213,
   R => '0',
   Q => M_reg_6_10
);
M_reg_6_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_212,
   R => '0',
   Q => M_reg_6_11
);
M_reg_6_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_211,
   R => '0',
   Q => M_reg_6_12
);
M_reg_6_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_210,
   R => '0',
   Q => M_reg_6_13
);
M_reg_6_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_209,
   R => '0',
   Q => M_reg_6_14
);
M_reg_6_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_208,
   R => '0',
   Q => M_reg_6_15
);
M_reg_6_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_207,
   R => '0',
   Q => M_reg_6_16
);
M_reg_6_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_206,
   R => '0',
   Q => M_reg_6_17
);
M_reg_6_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_205,
   R => '0',
   Q => M_reg_6_18
);
M_reg_6_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_204,
   R => '0',
   Q => M_reg_6_19
);
M_reg_6_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_222,
   R => '0',
   Q => M_reg_6_1
);
M_reg_6_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_203,
   R => '0',
   Q => M_reg_6_20
);
M_reg_6_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_202,
   R => '0',
   Q => M_reg_6_21
);
M_reg_6_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_201,
   R => '0',
   Q => M_reg_6_22
);
M_reg_6_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_200,
   R => '0',
   Q => M_reg_6_23
);
M_reg_6_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_199,
   R => '0',
   Q => M_reg_6_24
);
M_reg_6_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_198,
   R => '0',
   Q => M_reg_6_25
);
M_reg_6_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_197,
   R => '0',
   Q => M_reg_6_26
);
M_reg_6_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_196,
   R => '0',
   Q => M_reg_6_27
);
M_reg_6_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_195,
   R => '0',
   Q => M_reg_6_28
);
M_reg_6_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_194,
   R => '0',
   Q => M_reg_6_29
);
M_reg_6_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_221,
   R => '0',
   Q => M_reg_6_2
);
M_reg_6_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_193,
   R => '0',
   Q => M_reg_6_30
);
M_reg_6_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_192,
   R => '0',
   Q => M_reg_6_31
);
M_reg_6_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_220,
   R => '0',
   Q => M_reg_6_3
);
M_reg_6_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_219,
   R => '0',
   Q => M_reg_6_4
);
M_reg_6_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_218,
   R => '0',
   Q => M_reg_6_5
);
M_reg_6_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_217,
   R => '0',
   Q => M_reg_6_6
);
M_reg_6_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_216,
   R => '0',
   Q => M_reg_6_7
);
M_reg_6_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_215,
   R => '0',
   Q => M_reg_6_8
);
M_reg_6_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_214,
   R => '0',
   Q => M_reg_6_9
);
M_reg_7_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_255,
   R => '0',
   Q => M_reg_7_0
);
M_reg_7_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_245,
   R => '0',
   Q => M_reg_7_10
);
M_reg_7_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_244,
   R => '0',
   Q => M_reg_7_11
);
M_reg_7_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_243,
   R => '0',
   Q => M_reg_7_12
);
M_reg_7_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_242,
   R => '0',
   Q => M_reg_7_13
);
M_reg_7_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_241,
   R => '0',
   Q => M_reg_7_14
);
M_reg_7_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_240,
   R => '0',
   Q => M_reg_7_15
);
M_reg_7_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_239,
   R => '0',
   Q => M_reg_7_16
);
M_reg_7_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_238,
   R => '0',
   Q => M_reg_7_17
);
M_reg_7_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_237,
   R => '0',
   Q => M_reg_7_18
);
M_reg_7_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_236,
   R => '0',
   Q => M_reg_7_19
);
M_reg_7_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_254,
   R => '0',
   Q => M_reg_7_1
);
M_reg_7_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_235,
   R => '0',
   Q => M_reg_7_20
);
M_reg_7_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_234,
   R => '0',
   Q => M_reg_7_21
);
M_reg_7_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_233,
   R => '0',
   Q => M_reg_7_22
);
M_reg_7_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_232,
   R => '0',
   Q => M_reg_7_23
);
M_reg_7_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_231,
   R => '0',
   Q => M_reg_7_24
);
M_reg_7_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_230,
   R => '0',
   Q => M_reg_7_25
);
M_reg_7_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_229,
   R => '0',
   Q => M_reg_7_26
);
M_reg_7_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_228,
   R => '0',
   Q => M_reg_7_27
);
M_reg_7_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_227,
   R => '0',
   Q => M_reg_7_28
);
M_reg_7_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_226,
   R => '0',
   Q => M_reg_7_29
);
M_reg_7_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_253,
   R => '0',
   Q => M_reg_7_2
);
M_reg_7_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_225,
   R => '0',
   Q => M_reg_7_30
);
M_reg_7_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_224,
   R => '0',
   Q => M_reg_7_31
);
M_reg_7_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_252,
   R => '0',
   Q => M_reg_7_3
);
M_reg_7_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_251,
   R => '0',
   Q => M_reg_7_4
);
M_reg_7_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_250,
   R => '0',
   Q => M_reg_7_5
);
M_reg_7_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_249,
   R => '0',
   Q => M_reg_7_6
);
M_reg_7_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_248,
   R => '0',
   Q => M_reg_7_7
);
M_reg_7_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_247,
   R => '0',
   Q => M_reg_7_8
);
M_reg_7_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_246,
   R => '0',
   Q => M_reg_7_9
);
M_reg_8_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_287,
   R => '0',
   Q => M_reg_8_0
);
M_reg_8_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_277,
   R => '0',
   Q => M_reg_8_10
);
M_reg_8_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_276,
   R => '0',
   Q => M_reg_8_11
);
M_reg_8_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_275,
   R => '0',
   Q => M_reg_8_12
);
M_reg_8_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_274,
   R => '0',
   Q => M_reg_8_13
);
M_reg_8_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_273,
   R => '0',
   Q => M_reg_8_14
);
M_reg_8_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_272,
   R => '0',
   Q => M_reg_8_15
);
M_reg_8_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_271,
   R => '0',
   Q => M_reg_8_16
);
M_reg_8_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_270,
   R => '0',
   Q => M_reg_8_17
);
M_reg_8_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_269,
   R => '0',
   Q => M_reg_8_18
);
M_reg_8_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_268,
   R => '0',
   Q => M_reg_8_19
);
M_reg_8_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_286,
   R => '0',
   Q => M_reg_8_1
);
M_reg_8_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_267,
   R => '0',
   Q => M_reg_8_20
);
M_reg_8_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_266,
   R => '0',
   Q => M_reg_8_21
);
M_reg_8_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_265,
   R => '0',
   Q => M_reg_8_22
);
M_reg_8_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_264,
   R => '0',
   Q => M_reg_8_23
);
M_reg_8_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_263,
   R => '0',
   Q => M_reg_8_24
);
M_reg_8_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_262,
   R => '0',
   Q => M_reg_8_25
);
M_reg_8_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_261,
   R => '0',
   Q => M_reg_8_26
);
M_reg_8_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_260,
   R => '0',
   Q => M_reg_8_27
);
M_reg_8_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_259,
   R => '0',
   Q => M_reg_8_28
);
M_reg_8_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_258,
   R => '0',
   Q => M_reg_8_29
);
M_reg_8_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_285,
   R => '0',
   Q => M_reg_8_2
);
M_reg_8_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_257,
   R => '0',
   Q => M_reg_8_30
);
M_reg_8_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_256,
   R => '0',
   Q => M_reg_8_31
);
M_reg_8_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_284,
   R => '0',
   Q => M_reg_8_3
);
M_reg_8_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_283,
   R => '0',
   Q => M_reg_8_4
);
M_reg_8_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_282,
   R => '0',
   Q => M_reg_8_5
);
M_reg_8_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_281,
   R => '0',
   Q => M_reg_8_6
);
M_reg_8_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_280,
   R => '0',
   Q => M_reg_8_7
);
M_reg_8_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_279,
   R => '0',
   Q => M_reg_8_8
);
M_reg_8_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_278,
   R => '0',
   Q => M_reg_8_9
);
M_reg_9_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_319,
   R => '0',
   Q => M_reg_9_0
);
M_reg_9_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_309,
   R => '0',
   Q => M_reg_9_10
);
M_reg_9_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_308,
   R => '0',
   Q => M_reg_9_11
);
M_reg_9_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_307,
   R => '0',
   Q => M_reg_9_12
);
M_reg_9_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_306,
   R => '0',
   Q => M_reg_9_13
);
M_reg_9_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_305,
   R => '0',
   Q => M_reg_9_14
);
M_reg_9_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_304,
   R => '0',
   Q => M_reg_9_15
);
M_reg_9_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_303,
   R => '0',
   Q => M_reg_9_16
);
M_reg_9_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_302,
   R => '0',
   Q => M_reg_9_17
);
M_reg_9_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_301,
   R => '0',
   Q => M_reg_9_18
);
M_reg_9_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_300,
   R => '0',
   Q => M_reg_9_19
);
M_reg_9_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_318,
   R => '0',
   Q => M_reg_9_1
);
M_reg_9_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_299,
   R => '0',
   Q => M_reg_9_20
);
M_reg_9_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_298,
   R => '0',
   Q => M_reg_9_21
);
M_reg_9_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_297,
   R => '0',
   Q => M_reg_9_22
);
M_reg_9_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_296,
   R => '0',
   Q => M_reg_9_23
);
M_reg_9_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_295,
   R => '0',
   Q => M_reg_9_24
);
M_reg_9_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_294,
   R => '0',
   Q => M_reg_9_25
);
M_reg_9_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_293,
   R => '0',
   Q => M_reg_9_26
);
M_reg_9_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_292,
   R => '0',
   Q => M_reg_9_27
);
M_reg_9_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_291,
   R => '0',
   Q => M_reg_9_28
);
M_reg_9_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_290,
   R => '0',
   Q => M_reg_9_29
);
M_reg_9_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_317,
   R => '0',
   Q => M_reg_9_2
);
M_reg_9_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_289,
   R => '0',
   Q => M_reg_9_30
);
M_reg_9_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_288,
   R => '0',
   Q => M_reg_9_31
);
M_reg_9_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_316,
   R => '0',
   Q => M_reg_9_3
);
M_reg_9_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_315,
   R => '0',
   Q => M_reg_9_4
);
M_reg_9_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_314,
   R => '0',
   Q => M_reg_9_5
);
M_reg_9_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_313,
   R => '0',
   Q => M_reg_9_6
);
M_reg_9_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_312,
   R => '0',
   Q => M_reg_9_7
);
M_reg_9_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_311,
   R => '0',
   Q => M_reg_9_8
);
M_reg_9_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => M_reg_0_0,
   D => msg_block_in_IBUF_310,
   R => '0',
   Q => M_reg_9_9
);
rst_IBUF_inst : IBUF
 port map (
   I => rst,
   O => rst_IBUF
);
T1_11_i_10 : LUT3
  generic map(
   INIT => X"b8"
  )
 port map (
   I0 => f_reg_n_0_10,
   I1 => ROTR11_out_1,
   I2 => g_reg_n_0_10,
   O => T1_11_i_10_n_0
);
T1_11_i_100 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_27_3,
   I1 => W_reg_26_3,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_25_3,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_24_3,
   O => T1_11_i_100_n_0
);
T1_11_i_101 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_19_3,
   I1 => W_reg_18_3,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_17_3,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_16_3,
   O => T1_11_i_101_n_0
);
T1_11_i_102 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_23_3,
   I1 => W_reg_22_3,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_21_3,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_20_3,
   O => T1_11_i_102_n_0
);
T1_11_i_103 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_11_3,
   I1 => W_reg_10_3,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_9_3,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_8_3,
   O => T1_11_i_103_n_0
);
T1_11_i_104 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_15_3,
   I1 => W_reg_14_3,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_13_3,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_12_3,
   O => T1_11_i_104_n_0
);
T1_11_i_105 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_3_3,
   I1 => W_reg_2_3,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_1_3,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_0_3,
   O => T1_11_i_105_n_0
);
T1_11_i_106 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_7_3,
   I1 => W_reg_6_3,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_5_3,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_4_3,
   O => T1_11_i_106_n_0
);
T1_11_i_11 : LUT3
  generic map(
   INIT => X"b8"
  )
 port map (
   I0 => f_reg_n_0_9,
   I1 => ROTR11_out_2,
   I2 => g_reg_n_0_9,
   O => T1_11_i_11_n_0
);
T1_11_i_12 : LUT3
  generic map(
   INIT => X"b8"
  )
 port map (
   I0 => f_reg_n_0_8,
   I1 => ROTR11_out_3,
   I2 => g_reg_n_0_8,
   O => T1_11_i_12_n_0
);
T1_11_i_14 : LUT3
  generic map(
   INIT => X"b8"
  )
 port map (
   I0 => f_reg_n_0_7,
   I1 => ROTR11_out_4,
   I2 => g_reg_n_0_7,
   O => T1_11_i_14_n_0
);
T1_11_i_15 : LUT3
  generic map(
   INIT => X"e8"
  )
 port map (
   I0 => g0_b6_n_0,
   I1 => T1_11_i_23_n_0,
   I2 => h_6,
   O => T1_11_i_15_n_0
);
T1_11_i_16 : LUT3
  generic map(
   INIT => X"e8"
  )
 port map (
   I0 => g0_b5_n_0,
   I1 => T1_11_i_24_n_0,
   I2 => h_5,
   O => T1_11_i_16_n_0
);
T1_11_i_17 : LUT3
  generic map(
   INIT => X"e8"
  )
 port map (
   I0 => g0_b4_n_0,
   I1 => T1_11_i_25_n_0,
   I2 => h_4,
   O => T1_11_i_17_n_0
);
T1_11_i_18 : LUT3
  generic map(
   INIT => X"e8"
  )
 port map (
   I0 => g0_b3_n_0,
   I1 => T1_11_i_26_n_0,
   I2 => h_3,
   O => T1_11_i_18_n_0
);
T1_11_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => g0_b7_n_0,
   I1 => T1_15_i_26_n_0,
   I2 => h_7,
   I3 => T1_11_i_15_n_0,
   O => T1_11_i_19_n_0
);
T1_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => ROTR11_out_27,
   I1 => ROTR11_out_22,
   I2 => ROTR11_out_8,
   I3 => T1_reg_15_i_13_n_5,
   I4 => T1_11_i_10_n_0,
   O => T1_11_i_2_n_0
);
T1_11_i_20 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => g0_b6_n_0,
   I1 => T1_11_i_23_n_0,
   I2 => h_6,
   I3 => T1_11_i_16_n_0,
   O => T1_11_i_20_n_0
);
T1_11_i_21 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => g0_b5_n_0,
   I1 => T1_11_i_24_n_0,
   I2 => h_5,
   I3 => T1_11_i_17_n_0,
   O => T1_11_i_21_n_0
);
T1_11_i_22 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => g0_b4_n_0,
   I1 => T1_11_i_25_n_0,
   I2 => h_4,
   I3 => T1_11_i_18_n_0,
   O => T1_11_i_22_n_0
);
T1_11_i_23 : LUT6
  generic map(
   INIT => X"505f505f30303f3f"
  )
 port map (
   I0 => T1_11_i_27_n_0,
   I1 => T1_11_i_28_n_0,
   I2 => HASH_02_COUNTER_5,
   I3 => T1_11_i_29_n_0,
   I4 => T1_11_i_30_n_0,
   I5 => HASH_02_COUNTER_4,
   O => T1_11_i_23_n_0
);
T1_11_i_24 : LUT6
  generic map(
   INIT => X"505f505f30303f3f"
  )
 port map (
   I0 => T1_11_i_31_n_0,
   I1 => T1_11_i_32_n_0,
   I2 => HASH_02_COUNTER_5,
   I3 => T1_11_i_33_n_0,
   I4 => T1_11_i_34_n_0,
   I5 => HASH_02_COUNTER_4,
   O => T1_11_i_24_n_0
);
T1_11_i_25 : LUT6
  generic map(
   INIT => X"303f303f50505f5f"
  )
 port map (
   I0 => T1_11_i_35_n_0,
   I1 => T1_11_i_36_n_0,
   I2 => HASH_02_COUNTER_5,
   I3 => T1_11_i_37_n_0,
   I4 => T1_11_i_38_n_0,
   I5 => HASH_02_COUNTER_4,
   O => T1_11_i_25_n_0
);
T1_11_i_26 : LUT6
  generic map(
   INIT => X"303f303f50505f5f"
  )
 port map (
   I0 => T1_11_i_39_n_0,
   I1 => T1_11_i_40_n_0,
   I2 => HASH_02_COUNTER_5,
   I3 => T1_11_i_41_n_0,
   I4 => T1_11_i_42_n_0,
   I5 => HASH_02_COUNTER_4,
   O => T1_11_i_26_n_0
);
T1_11_i_27 : LUT6
  generic map(
   INIT => X"303f5050303f5f5f"
  )
 port map (
   I0 => T1_11_i_43_n_0,
   I1 => T1_11_i_44_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_11_i_45_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_11_i_46_n_0,
   O => T1_11_i_27_n_0
);
T1_11_i_28 : LUT6
  generic map(
   INIT => X"5050303f5f5f303f"
  )
 port map (
   I0 => T1_11_i_47_n_0,
   I1 => T1_11_i_48_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_11_i_49_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_11_i_50_n_0,
   O => T1_11_i_28_n_0
);
T1_11_i_29 : LUT6
  generic map(
   INIT => X"5050303f5f5f303f"
  )
 port map (
   I0 => T1_11_i_51_n_0,
   I1 => T1_11_i_52_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_11_i_53_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_11_i_54_n_0,
   O => T1_11_i_29_n_0
);
T1_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => ROTR11_out_28,
   I1 => ROTR11_out_23,
   I2 => ROTR11_out_9,
   I3 => T1_reg_15_i_13_n_6,
   I4 => T1_11_i_11_n_0,
   O => T1_11_i_3_n_0
);
T1_11_i_30 : LUT6
  generic map(
   INIT => X"303f5050303f5f5f"
  )
 port map (
   I0 => T1_11_i_55_n_0,
   I1 => T1_11_i_56_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_11_i_57_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_11_i_58_n_0,
   O => T1_11_i_30_n_0
);
T1_11_i_31 : LUT6
  generic map(
   INIT => X"303f5050303f5f5f"
  )
 port map (
   I0 => T1_11_i_59_n_0,
   I1 => T1_11_i_60_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_11_i_61_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_11_i_62_n_0,
   O => T1_11_i_31_n_0
);
T1_11_i_32 : LUT6
  generic map(
   INIT => X"3030505f3f3f505f"
  )
 port map (
   I0 => T1_11_i_63_n_0,
   I1 => T1_11_i_64_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_11_i_65_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_11_i_66_n_0,
   O => T1_11_i_32_n_0
);
T1_11_i_33 : LUT6
  generic map(
   INIT => X"5050303f5f5f303f"
  )
 port map (
   I0 => T1_11_i_67_n_0,
   I1 => T1_11_i_68_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_11_i_69_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_11_i_70_n_0,
   O => T1_11_i_33_n_0
);
T1_11_i_34 : LUT6
  generic map(
   INIT => X"303f5050303f5f5f"
  )
 port map (
   I0 => T1_11_i_71_n_0,
   I1 => T1_11_i_72_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_11_i_73_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_11_i_74_n_0,
   O => T1_11_i_34_n_0
);
T1_11_i_35 : LUT6
  generic map(
   INIT => X"5050303f5f5f303f"
  )
 port map (
   I0 => T1_11_i_75_n_0,
   I1 => T1_11_i_76_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_11_i_77_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_11_i_78_n_0,
   O => T1_11_i_35_n_0
);
T1_11_i_36 : LUT6
  generic map(
   INIT => X"303f5050303f5f5f"
  )
 port map (
   I0 => T1_11_i_79_n_0,
   I1 => T1_11_i_80_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_11_i_81_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_11_i_82_n_0,
   O => T1_11_i_36_n_0
);
T1_11_i_37 : LUT6
  generic map(
   INIT => X"5050303f5f5f303f"
  )
 port map (
   I0 => T1_11_i_83_n_0,
   I1 => T1_11_i_84_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_11_i_85_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_11_i_86_n_0,
   O => T1_11_i_37_n_0
);
T1_11_i_38 : LUT6
  generic map(
   INIT => X"505f3030505f3f3f"
  )
 port map (
   I0 => T1_11_i_87_n_0,
   I1 => T1_11_i_88_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_11_i_89_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_11_i_90_n_0,
   O => T1_11_i_38_n_0
);
T1_11_i_39 : LUT6
  generic map(
   INIT => X"303f5050303f5f5f"
  )
 port map (
   I0 => T1_11_i_91_n_0,
   I1 => T1_11_i_92_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_11_i_93_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_11_i_94_n_0,
   O => T1_11_i_39_n_0
);
T1_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => ROTR11_out_29,
   I1 => ROTR11_out_24,
   I2 => ROTR11_out_10,
   I3 => T1_reg_15_i_13_n_7,
   I4 => T1_11_i_12_n_0,
   O => T1_11_i_4_n_0
);
T1_11_i_40 : LUT6
  generic map(
   INIT => X"3030505f3f3f505f"
  )
 port map (
   I0 => T1_11_i_95_n_0,
   I1 => T1_11_i_96_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_11_i_97_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_11_i_98_n_0,
   O => T1_11_i_40_n_0
);
T1_11_i_41 : LUT6
  generic map(
   INIT => X"5050303f5f5f303f"
  )
 port map (
   I0 => T1_11_i_99_n_0,
   I1 => T1_11_i_100_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_11_i_101_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_11_i_102_n_0,
   O => T1_11_i_41_n_0
);
T1_11_i_42 : LUT6
  generic map(
   INIT => X"3030505f3f3f505f"
  )
 port map (
   I0 => T1_11_i_103_n_0,
   I1 => T1_11_i_104_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_11_i_105_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_11_i_106_n_0,
   O => T1_11_i_42_n_0
);
T1_11_i_43 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_59_6,
   I1 => W_reg_58_6,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_57_6,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_56_6,
   O => T1_11_i_43_n_0
);
T1_11_i_44 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_63_6,
   I1 => W_reg_62_6,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_61_6,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_60_6,
   O => T1_11_i_44_n_0
);
T1_11_i_45 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_55_6,
   I1 => W_reg_54_6,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_53_6,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_52_6,
   O => T1_11_i_45_n_0
);
T1_11_i_46 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_51_6,
   I1 => W_reg_50_6,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_49_6,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_48_6,
   O => T1_11_i_46_n_0
);
T1_11_i_47 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_47_6,
   I1 => W_reg_46_6,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_45_6,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_44_6,
   O => T1_11_i_47_n_0
);
T1_11_i_48 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_43_6,
   I1 => W_reg_42_6,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_41_6,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_40_6,
   O => T1_11_i_48_n_0
);
T1_11_i_49 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_35_6,
   I1 => W_reg_34_6,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_33_6,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_32_6,
   O => T1_11_i_49_n_0
);
T1_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => ROTR11_out_25,
   I1 => ROTR11_out_11,
   I2 => ROTR11_out_30,
   I3 => T1_reg_11_i_13_n_4,
   I4 => T1_11_i_14_n_0,
   O => T1_11_i_5_n_0
);
T1_11_i_50 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_39_6,
   I1 => W_reg_38_6,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_37_6,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_36_6,
   O => T1_11_i_50_n_0
);
T1_11_i_51 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_31_6,
   I1 => W_reg_30_6,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_29_6,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_28_6,
   O => T1_11_i_51_n_0
);
T1_11_i_52 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_27_6,
   I1 => W_reg_26_6,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_25_6,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_24_6,
   O => T1_11_i_52_n_0
);
T1_11_i_53 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_19_6,
   I1 => W_reg_18_6,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_17_6,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_16_6,
   O => T1_11_i_53_n_0
);
T1_11_i_54 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_23_6,
   I1 => W_reg_22_6,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_21_6,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_20_6,
   O => T1_11_i_54_n_0
);
T1_11_i_55 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_11_6,
   I1 => W_reg_10_6,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_9_6,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_8_6,
   O => T1_11_i_55_n_0
);
T1_11_i_56 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_15_6,
   I1 => W_reg_14_6,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_13_6,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_12_6,
   O => T1_11_i_56_n_0
);
T1_11_i_57 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_7_6,
   I1 => W_reg_6_6,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_5_6,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_4_6,
   O => T1_11_i_57_n_0
);
T1_11_i_58 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_3_6,
   I1 => W_reg_2_6,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_1_6,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_0_6,
   O => T1_11_i_58_n_0
);
T1_11_i_59 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_59_5,
   I1 => W_reg_58_5,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_57_5,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_56_5,
   O => T1_11_i_59_n_0
);
T1_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => T1_11_i_2_n_0,
   I1 => ROTR11_out_26,
   I2 => ROTR11_out_21,
   I3 => ROTR11_out_7,
   I4 => T1_reg_15_i_13_n_4,
   I5 => T1_15_i_14_n_0,
   O => T1_11_i_6_n_0
);
T1_11_i_60 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_63_5,
   I1 => W_reg_62_5,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_61_5,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_60_5,
   O => T1_11_i_60_n_0
);
T1_11_i_61 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_55_5,
   I1 => W_reg_54_5,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_53_5,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_52_5,
   O => T1_11_i_61_n_0
);
T1_11_i_62 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_51_5,
   I1 => W_reg_50_5,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_49_5,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_48_5,
   O => T1_11_i_62_n_0
);
T1_11_i_63 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_43_5,
   I1 => W_reg_42_5,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_41_5,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_40_5,
   O => T1_11_i_63_n_0
);
T1_11_i_64 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_47_5,
   I1 => W_reg_46_5,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_45_5,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_44_5,
   O => T1_11_i_64_n_0
);
T1_11_i_65 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_35_5,
   I1 => W_reg_34_5,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_33_5,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_32_5,
   O => T1_11_i_65_n_0
);
T1_11_i_66 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_39_5,
   I1 => W_reg_38_5,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_37_5,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_36_5,
   O => T1_11_i_66_n_0
);
T1_11_i_67 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_31_5,
   I1 => W_reg_30_5,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_29_5,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_28_5,
   O => T1_11_i_67_n_0
);
T1_11_i_68 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_27_5,
   I1 => W_reg_26_5,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_25_5,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_24_5,
   O => T1_11_i_68_n_0
);
T1_11_i_69 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_19_5,
   I1 => W_reg_18_5,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_17_5,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_16_5,
   O => T1_11_i_69_n_0
);
T1_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => T1_11_i_3_n_0,
   I1 => T1_reg_15_i_13_n_5,
   I2 => T1_11_i_10_n_0,
   I3 => ROTR11_out_27,
   I4 => ROTR11_out_22,
   I5 => ROTR11_out_8,
   O => T1_11_i_7_n_0
);
T1_11_i_70 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_23_5,
   I1 => W_reg_22_5,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_21_5,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_20_5,
   O => T1_11_i_70_n_0
);
T1_11_i_71 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_11_5,
   I1 => W_reg_10_5,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_9_5,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_8_5,
   O => T1_11_i_71_n_0
);
T1_11_i_72 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_15_5,
   I1 => W_reg_14_5,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_13_5,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_12_5,
   O => T1_11_i_72_n_0
);
T1_11_i_73 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_7_5,
   I1 => W_reg_6_5,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_5_5,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_4_5,
   O => T1_11_i_73_n_0
);
T1_11_i_74 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_3_5,
   I1 => W_reg_2_5,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_1_5,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_0_5,
   O => T1_11_i_74_n_0
);
T1_11_i_75 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_47_4,
   I1 => W_reg_46_4,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_45_4,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_44_4,
   O => T1_11_i_75_n_0
);
T1_11_i_76 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_43_4,
   I1 => W_reg_42_4,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_41_4,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_40_4,
   O => T1_11_i_76_n_0
);
T1_11_i_77 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_35_4,
   I1 => W_reg_34_4,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_33_4,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_32_4,
   O => T1_11_i_77_n_0
);
T1_11_i_78 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_39_4,
   I1 => W_reg_38_4,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_37_4,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_36_4,
   O => T1_11_i_78_n_0
);
T1_11_i_79 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_59_4,
   I1 => W_reg_58_4,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_57_4,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_56_4,
   O => T1_11_i_79_n_0
);
T1_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => T1_11_i_4_n_0,
   I1 => ROTR11_out_28,
   I2 => ROTR11_out_23,
   I3 => ROTR11_out_9,
   I4 => T1_reg_15_i_13_n_6,
   I5 => T1_11_i_11_n_0,
   O => T1_11_i_8_n_0
);
T1_11_i_80 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_63_4,
   I1 => W_reg_62_4,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_61_4,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_60_4,
   O => T1_11_i_80_n_0
);
T1_11_i_81 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_55_4,
   I1 => W_reg_54_4,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_53_4,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_52_4,
   O => T1_11_i_81_n_0
);
T1_11_i_82 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_51_4,
   I1 => W_reg_50_4,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_49_4,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_48_4,
   O => T1_11_i_82_n_0
);
T1_11_i_83 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_31_4,
   I1 => W_reg_30_4,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_29_4,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_28_4,
   O => T1_11_i_83_n_0
);
T1_11_i_84 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_27_4,
   I1 => W_reg_26_4,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_25_4,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_24_4,
   O => T1_11_i_84_n_0
);
T1_11_i_85 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_19_4,
   I1 => W_reg_18_4,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_17_4,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_16_4,
   O => T1_11_i_85_n_0
);
T1_11_i_86 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_23_4,
   I1 => W_reg_22_4,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_21_4,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_20_4,
   O => T1_11_i_86_n_0
);
T1_11_i_87 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_15_4,
   I1 => W_reg_14_4,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_13_4,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_12_4,
   O => T1_11_i_87_n_0
);
T1_11_i_88 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_11_4,
   I1 => W_reg_10_4,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_9_4,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_8_4,
   O => T1_11_i_88_n_0
);
T1_11_i_89 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_7_4,
   I1 => W_reg_6_4,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_5_4,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_4_4,
   O => T1_11_i_89_n_0
);
T1_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => T1_11_i_5_n_0,
   I1 => T1_reg_15_i_13_n_7,
   I2 => T1_11_i_12_n_0,
   I3 => ROTR11_out_29,
   I4 => ROTR11_out_24,
   I5 => ROTR11_out_10,
   O => T1_11_i_9_n_0
);
T1_11_i_90 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_3_4,
   I1 => W_reg_2_4,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_1_4,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_0_4,
   O => T1_11_i_90_n_0
);
T1_11_i_91 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_43_3,
   I1 => W_reg_42_3,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_41_3,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_40_3,
   O => T1_11_i_91_n_0
);
T1_11_i_92 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_47_3,
   I1 => W_reg_46_3,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_45_3,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_44_3,
   O => T1_11_i_92_n_0
);
T1_11_i_93 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_39_3,
   I1 => W_reg_38_3,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_37_3,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_36_3,
   O => T1_11_i_93_n_0
);
T1_11_i_94 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_35_3,
   I1 => W_reg_34_3,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_33_3,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_32_3,
   O => T1_11_i_94_n_0
);
T1_11_i_95 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_59_3,
   I1 => W_reg_58_3,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_57_3,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_56_3,
   O => T1_11_i_95_n_0
);
T1_11_i_96 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_63_3,
   I1 => W_reg_62_3,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_61_3,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_60_3,
   O => T1_11_i_96_n_0
);
T1_11_i_97 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_51_3,
   I1 => W_reg_50_3,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_49_3,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_48_3,
   O => T1_11_i_97_n_0
);
T1_11_i_98 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_55_3,
   I1 => W_reg_54_3,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_53_3,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_52_3,
   O => T1_11_i_98_n_0
);
T1_11_i_99 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_31_3,
   I1 => W_reg_30_3,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_29_3,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_28_3,
   O => T1_11_i_99_n_0
);
T1_15_i_10 : LUT3
  generic map(
   INIT => X"b8"
  )
 port map (
   I0 => f_reg_n_0_14,
   I1 => ROTR11_out_29,
   I2 => g_reg_n_0_14,
   O => T1_15_i_10_n_0
);
T1_15_i_100 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_3_7,
   I1 => W_reg_2_7,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_1_7,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_0_7,
   O => T1_15_i_100_n_0
);
T1_15_i_101 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_3_10,
   I1 => W_reg_2_10,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_1_10,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_0_10,
   O => T1_15_i_101_n_0
);
T1_15_i_102 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_7_10,
   I1 => W_reg_6_10,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_5_10,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_4_10,
   O => T1_15_i_102_n_0
);
T1_15_i_103 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_11_10,
   I1 => W_reg_10_10,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_9_10,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_8_10,
   O => T1_15_i_103_n_0
);
T1_15_i_104 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_15_10,
   I1 => W_reg_14_10,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_13_10,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_12_10,
   O => T1_15_i_104_n_0
);
T1_15_i_105 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_3_9,
   I1 => W_reg_2_9,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_1_9,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_0_9,
   O => T1_15_i_105_n_0
);
T1_15_i_106 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_7_9,
   I1 => W_reg_6_9,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_5_9,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_4_9,
   O => T1_15_i_106_n_0
);
T1_15_i_107 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_11_9,
   I1 => W_reg_10_9,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_9_9,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_8_9,
   O => T1_15_i_107_n_0
);
T1_15_i_108 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_15_9,
   I1 => W_reg_14_9,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_13_9,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_12_9,
   O => T1_15_i_108_n_0
);
T1_15_i_109 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_3_8,
   I1 => W_reg_2_8,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_1_8,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_0_8,
   O => T1_15_i_109_n_0
);
T1_15_i_11 : LUT3
  generic map(
   INIT => X"b8"
  )
 port map (
   I0 => f_reg_n_0_13,
   I1 => ROTR11_out_30,
   I2 => g_reg_n_0_13,
   O => T1_15_i_11_n_0
);
T1_15_i_110 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_7_8,
   I1 => W_reg_6_8,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_5_8,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_4_8,
   O => T1_15_i_110_n_0
);
T1_15_i_111 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_11_8,
   I1 => W_reg_10_8,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_9_8,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_8_8,
   O => T1_15_i_111_n_0
);
T1_15_i_112 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_15_8,
   I1 => W_reg_14_8,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_13_8,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_12_8,
   O => T1_15_i_112_n_0
);
T1_15_i_12 : LUT3
  generic map(
   INIT => X"b8"
  )
 port map (
   I0 => f_reg_n_0_12,
   I1 => ROTR11_out_31,
   I2 => g_reg_n_0_12,
   O => T1_15_i_12_n_0
);
T1_15_i_14 : LUT3
  generic map(
   INIT => X"b8"
  )
 port map (
   I0 => f_reg_n_0_11,
   I1 => ROTR11_out_32,
   I2 => g_reg_n_0_11,
   O => T1_15_i_14_n_0
);
T1_15_i_15 : LUT3
  generic map(
   INIT => X"e8"
  )
 port map (
   I0 => g0_b10_n_0,
   I1 => T1_15_i_23_n_0,
   I2 => h_10,
   O => T1_15_i_15_n_0
);
T1_15_i_16 : LUT3
  generic map(
   INIT => X"e8"
  )
 port map (
   I0 => g0_b9_n_0,
   I1 => T1_15_i_24_n_0,
   I2 => h_9,
   O => T1_15_i_16_n_0
);
T1_15_i_17 : LUT3
  generic map(
   INIT => X"e8"
  )
 port map (
   I0 => g0_b8_n_0,
   I1 => T1_15_i_25_n_0,
   I2 => h_8,
   O => T1_15_i_17_n_0
);
T1_15_i_18 : LUT3
  generic map(
   INIT => X"e8"
  )
 port map (
   I0 => g0_b7_n_0,
   I1 => T1_15_i_26_n_0,
   I2 => h_7,
   O => T1_15_i_18_n_0
);
T1_15_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => g0_b11_n_0,
   I1 => T1_19_i_26_n_0,
   I2 => h_11,
   I3 => T1_15_i_15_n_0,
   O => T1_15_i_19_n_0
);
T1_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => ROTR11_out_18,
   I1 => ROTR11_out_23,
   I2 => ROTR11_out_4,
   I3 => T1_reg_19_i_13_n_5,
   I4 => T1_15_i_10_n_0,
   O => T1_15_i_2_n_0
);
T1_15_i_20 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => g0_b10_n_0,
   I1 => T1_15_i_23_n_0,
   I2 => h_10,
   I3 => T1_15_i_16_n_0,
   O => T1_15_i_20_n_0
);
T1_15_i_21 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => g0_b9_n_0,
   I1 => T1_15_i_24_n_0,
   I2 => h_9,
   I3 => T1_15_i_17_n_0,
   O => T1_15_i_21_n_0
);
T1_15_i_22 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => g0_b8_n_0,
   I1 => T1_15_i_25_n_0,
   I2 => h_8,
   I3 => T1_15_i_18_n_0,
   O => T1_15_i_22_n_0
);
T1_15_i_23 : LUT6
  generic map(
   INIT => X"50505f5f3f303f30"
  )
 port map (
   I0 => T1_15_i_27_n_0,
   I1 => T1_15_i_28_n_0,
   I2 => HASH_02_COUNTER_5,
   I3 => T1_reg_15_i_29_n_0,
   I4 => T1_15_i_30_n_0,
   I5 => HASH_02_COUNTER_4,
   O => T1_15_i_23_n_0
);
T1_15_i_24 : LUT6
  generic map(
   INIT => X"50505f5f3f303f30"
  )
 port map (
   I0 => T1_15_i_31_n_0,
   I1 => T1_15_i_32_n_0,
   I2 => HASH_02_COUNTER_5,
   I3 => T1_reg_15_i_33_n_0,
   I4 => T1_15_i_34_n_0,
   I5 => HASH_02_COUNTER_4,
   O => T1_15_i_24_n_0
);
T1_15_i_25 : LUT6
  generic map(
   INIT => X"50505f5f3f303f30"
  )
 port map (
   I0 => T1_15_i_35_n_0,
   I1 => T1_15_i_36_n_0,
   I2 => HASH_02_COUNTER_5,
   I3 => T1_reg_15_i_37_n_0,
   I4 => T1_15_i_38_n_0,
   I5 => HASH_02_COUNTER_4,
   O => T1_15_i_25_n_0
);
T1_15_i_26 : LUT6
  generic map(
   INIT => X"505f505f30303f3f"
  )
 port map (
   I0 => T1_15_i_39_n_0,
   I1 => T1_15_i_40_n_0,
   I2 => HASH_02_COUNTER_5,
   I3 => T1_15_i_41_n_0,
   I4 => T1_15_i_42_n_0,
   I5 => HASH_02_COUNTER_4,
   O => T1_15_i_26_n_0
);
T1_15_i_27 : LUT6
  generic map(
   INIT => X"505f3030505f3f3f"
  )
 port map (
   I0 => T1_15_i_43_n_0,
   I1 => T1_15_i_44_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_15_i_45_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_15_i_46_n_0,
   O => T1_15_i_27_n_0
);
T1_15_i_28 : LUT6
  generic map(
   INIT => X"3030505f3f3f505f"
  )
 port map (
   I0 => T1_15_i_47_n_0,
   I1 => T1_15_i_48_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_15_i_49_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_15_i_50_n_0,
   O => T1_15_i_28_n_0
);
T1_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => ROTR11_out_5,
   I1 => ROTR11_out_19,
   I2 => ROTR11_out_24,
   I3 => T1_reg_19_i_13_n_6,
   I4 => T1_15_i_11_n_0,
   O => T1_15_i_3_n_0
);
T1_15_i_30 : LUT6
  generic map(
   INIT => X"3030505f3f3f505f"
  )
 port map (
   I0 => T1_15_i_53_n_0,
   I1 => T1_15_i_54_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_15_i_55_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_15_i_56_n_0,
   O => T1_15_i_30_n_0
);
T1_15_i_31 : LUT6
  generic map(
   INIT => X"303f5050303f5f5f"
  )
 port map (
   I0 => T1_15_i_57_n_0,
   I1 => T1_15_i_58_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_15_i_59_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_15_i_60_n_0,
   O => T1_15_i_31_n_0
);
T1_15_i_32 : LUT6
  generic map(
   INIT => X"3030505f3f3f505f"
  )
 port map (
   I0 => T1_15_i_61_n_0,
   I1 => T1_15_i_62_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_15_i_63_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_15_i_64_n_0,
   O => T1_15_i_32_n_0
);
T1_15_i_34 : LUT6
  generic map(
   INIT => X"3030505f3f3f505f"
  )
 port map (
   I0 => T1_15_i_67_n_0,
   I1 => T1_15_i_68_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_15_i_69_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_15_i_70_n_0,
   O => T1_15_i_34_n_0
);
T1_15_i_35 : LUT6
  generic map(
   INIT => X"303f5050303f5f5f"
  )
 port map (
   I0 => T1_15_i_71_n_0,
   I1 => T1_15_i_72_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_15_i_73_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_15_i_74_n_0,
   O => T1_15_i_35_n_0
);
T1_15_i_36 : LUT6
  generic map(
   INIT => X"5050303f5f5f303f"
  )
 port map (
   I0 => T1_15_i_75_n_0,
   I1 => T1_15_i_76_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_15_i_77_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_15_i_78_n_0,
   O => T1_15_i_36_n_0
);
T1_15_i_38 : LUT6
  generic map(
   INIT => X"3030505f3f3f505f"
  )
 port map (
   I0 => T1_15_i_81_n_0,
   I1 => T1_15_i_82_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_15_i_83_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_15_i_84_n_0,
   O => T1_15_i_38_n_0
);
T1_15_i_39 : LUT6
  generic map(
   INIT => X"303f5050303f5f5f"
  )
 port map (
   I0 => T1_15_i_85_n_0,
   I1 => T1_15_i_86_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_15_i_87_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_15_i_88_n_0,
   O => T1_15_i_39_n_0
);
T1_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => ROTR11_out_25,
   I1 => ROTR11_out_20,
   I2 => ROTR11_out_6,
   I3 => T1_reg_19_i_13_n_7,
   I4 => T1_15_i_12_n_0,
   O => T1_15_i_4_n_0
);
T1_15_i_40 : LUT6
  generic map(
   INIT => X"5050303f5f5f303f"
  )
 port map (
   I0 => T1_15_i_89_n_0,
   I1 => T1_15_i_90_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_15_i_91_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_15_i_92_n_0,
   O => T1_15_i_40_n_0
);
T1_15_i_41 : LUT6
  generic map(
   INIT => X"5050303f5f5f303f"
  )
 port map (
   I0 => T1_15_i_93_n_0,
   I1 => T1_15_i_94_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_15_i_95_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_15_i_96_n_0,
   O => T1_15_i_41_n_0
);
T1_15_i_42 : LUT6
  generic map(
   INIT => X"303f5050303f5f5f"
  )
 port map (
   I0 => T1_15_i_97_n_0,
   I1 => T1_15_i_98_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_15_i_99_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_15_i_100_n_0,
   O => T1_15_i_42_n_0
);
T1_15_i_43 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_63_10,
   I1 => W_reg_62_10,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_61_10,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_60_10,
   O => T1_15_i_43_n_0
);
T1_15_i_44 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_59_10,
   I1 => W_reg_58_10,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_57_10,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_56_10,
   O => T1_15_i_44_n_0
);
T1_15_i_45 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_55_10,
   I1 => W_reg_54_10,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_53_10,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_52_10,
   O => T1_15_i_45_n_0
);
T1_15_i_46 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_51_10,
   I1 => W_reg_50_10,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_49_10,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_48_10,
   O => T1_15_i_46_n_0
);
T1_15_i_47 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_43_10,
   I1 => W_reg_42_10,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_41_10,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_40_10,
   O => T1_15_i_47_n_0
);
T1_15_i_48 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_47_10,
   I1 => W_reg_46_10,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_45_10,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_44_10,
   O => T1_15_i_48_n_0
);
T1_15_i_49 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_35_10,
   I1 => W_reg_34_10,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_33_10,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_32_10,
   O => T1_15_i_49_n_0
);
T1_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => ROTR11_out_26,
   I1 => ROTR11_out_21,
   I2 => ROTR11_out_7,
   I3 => T1_reg_15_i_13_n_4,
   I4 => T1_15_i_14_n_0,
   O => T1_15_i_5_n_0
);
T1_15_i_50 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_39_10,
   I1 => W_reg_38_10,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_37_10,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_36_10,
   O => T1_15_i_50_n_0
);
T1_15_i_53 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_27_10,
   I1 => W_reg_26_10,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_25_10,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_24_10,
   O => T1_15_i_53_n_0
);
T1_15_i_54 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_31_10,
   I1 => W_reg_30_10,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_29_10,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_28_10,
   O => T1_15_i_54_n_0
);
T1_15_i_55 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_19_10,
   I1 => W_reg_18_10,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_17_10,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_16_10,
   O => T1_15_i_55_n_0
);
T1_15_i_56 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_23_10,
   I1 => W_reg_22_10,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_21_10,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_20_10,
   O => T1_15_i_56_n_0
);
T1_15_i_57 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_59_9,
   I1 => W_reg_58_9,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_57_9,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_56_9,
   O => T1_15_i_57_n_0
);
T1_15_i_58 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_63_9,
   I1 => W_reg_62_9,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_61_9,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_60_9,
   O => T1_15_i_58_n_0
);
T1_15_i_59 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_55_9,
   I1 => W_reg_54_9,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_53_9,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_52_9,
   O => T1_15_i_59_n_0
);
T1_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => T1_15_i_2_n_0,
   I1 => T1_reg_19_i_13_n_4,
   I2 => T1_19_i_14_n_0,
   I3 => ROTR11_out_17,
   I4 => ROTR11_out_22,
   I5 => ROTR11_out_3,
   O => T1_15_i_6_n_0
);
T1_15_i_60 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_51_9,
   I1 => W_reg_50_9,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_49_9,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_48_9,
   O => T1_15_i_60_n_0
);
T1_15_i_61 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_43_9,
   I1 => W_reg_42_9,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_41_9,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_40_9,
   O => T1_15_i_61_n_0
);
T1_15_i_62 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_47_9,
   I1 => W_reg_46_9,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_45_9,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_44_9,
   O => T1_15_i_62_n_0
);
T1_15_i_63 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_35_9,
   I1 => W_reg_34_9,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_33_9,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_32_9,
   O => T1_15_i_63_n_0
);
T1_15_i_64 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_39_9,
   I1 => W_reg_38_9,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_37_9,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_36_9,
   O => T1_15_i_64_n_0
);
T1_15_i_67 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_27_9,
   I1 => W_reg_26_9,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_25_9,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_24_9,
   O => T1_15_i_67_n_0
);
T1_15_i_68 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_31_9,
   I1 => W_reg_30_9,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_29_9,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_28_9,
   O => T1_15_i_68_n_0
);
T1_15_i_69 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_19_9,
   I1 => W_reg_18_9,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_17_9,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_16_9,
   O => T1_15_i_69_n_0
);
T1_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => T1_15_i_3_n_0,
   I1 => T1_reg_19_i_13_n_5,
   I2 => T1_15_i_10_n_0,
   I3 => ROTR11_out_18,
   I4 => ROTR11_out_23,
   I5 => ROTR11_out_4,
   O => T1_15_i_7_n_0
);
T1_15_i_70 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_23_9,
   I1 => W_reg_22_9,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_21_9,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_20_9,
   O => T1_15_i_70_n_0
);
T1_15_i_71 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_59_8,
   I1 => W_reg_58_8,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_57_8,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_56_8,
   O => T1_15_i_71_n_0
);
T1_15_i_72 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_63_8,
   I1 => W_reg_62_8,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_61_8,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_60_8,
   O => T1_15_i_72_n_0
);
T1_15_i_73 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_55_8,
   I1 => W_reg_54_8,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_53_8,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_52_8,
   O => T1_15_i_73_n_0
);
T1_15_i_74 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_51_8,
   I1 => W_reg_50_8,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_49_8,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_48_8,
   O => T1_15_i_74_n_0
);
T1_15_i_75 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_47_8,
   I1 => W_reg_46_8,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_45_8,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_44_8,
   O => T1_15_i_75_n_0
);
T1_15_i_76 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_43_8,
   I1 => W_reg_42_8,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_41_8,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_40_8,
   O => T1_15_i_76_n_0
);
T1_15_i_77 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_35_8,
   I1 => W_reg_34_8,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_33_8,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_32_8,
   O => T1_15_i_77_n_0
);
T1_15_i_78 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_39_8,
   I1 => W_reg_38_8,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_37_8,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_36_8,
   O => T1_15_i_78_n_0
);
T1_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => T1_15_i_4_n_0,
   I1 => ROTR11_out_5,
   I2 => ROTR11_out_19,
   I3 => ROTR11_out_24,
   I4 => T1_reg_19_i_13_n_6,
   I5 => T1_15_i_11_n_0,
   O => T1_15_i_8_n_0
);
T1_15_i_81 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_27_8,
   I1 => W_reg_26_8,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_25_8,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_24_8,
   O => T1_15_i_81_n_0
);
T1_15_i_82 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_31_8,
   I1 => W_reg_30_8,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_29_8,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_28_8,
   O => T1_15_i_82_n_0
);
T1_15_i_83 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_19_8,
   I1 => W_reg_18_8,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_17_8,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_16_8,
   O => T1_15_i_83_n_0
);
T1_15_i_84 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_23_8,
   I1 => W_reg_22_8,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_21_8,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_20_8,
   O => T1_15_i_84_n_0
);
T1_15_i_85 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_59_7,
   I1 => W_reg_58_7,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_57_7,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_56_7,
   O => T1_15_i_85_n_0
);
T1_15_i_86 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_63_7,
   I1 => W_reg_62_7,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_61_7,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_60_7,
   O => T1_15_i_86_n_0
);
T1_15_i_87 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_55_7,
   I1 => W_reg_54_7,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_53_7,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_52_7,
   O => T1_15_i_87_n_0
);
T1_15_i_88 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_51_7,
   I1 => W_reg_50_7,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_49_7,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_48_7,
   O => T1_15_i_88_n_0
);
T1_15_i_89 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_47_7,
   I1 => W_reg_46_7,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_45_7,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_44_7,
   O => T1_15_i_89_n_0
);
T1_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => T1_15_i_5_n_0,
   I1 => T1_reg_19_i_13_n_7,
   I2 => T1_15_i_12_n_0,
   I3 => ROTR11_out_25,
   I4 => ROTR11_out_20,
   I5 => ROTR11_out_6,
   O => T1_15_i_9_n_0
);
T1_15_i_90 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_43_7,
   I1 => W_reg_42_7,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_41_7,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_40_7,
   O => T1_15_i_90_n_0
);
T1_15_i_91 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_35_7,
   I1 => W_reg_34_7,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_33_7,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_32_7,
   O => T1_15_i_91_n_0
);
T1_15_i_92 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_39_7,
   I1 => W_reg_38_7,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_37_7,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_36_7,
   O => T1_15_i_92_n_0
);
T1_15_i_93 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_31_7,
   I1 => W_reg_30_7,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_29_7,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_28_7,
   O => T1_15_i_93_n_0
);
T1_15_i_94 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_27_7,
   I1 => W_reg_26_7,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_25_7,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_24_7,
   O => T1_15_i_94_n_0
);
T1_15_i_95 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_19_7,
   I1 => W_reg_18_7,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_17_7,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_16_7,
   O => T1_15_i_95_n_0
);
T1_15_i_96 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_23_7,
   I1 => W_reg_22_7,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_21_7,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_20_7,
   O => T1_15_i_96_n_0
);
T1_15_i_97 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_11_7,
   I1 => W_reg_10_7,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_9_7,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_8_7,
   O => T1_15_i_97_n_0
);
T1_15_i_98 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_15_7,
   I1 => W_reg_14_7,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_13_7,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_12_7,
   O => T1_15_i_98_n_0
);
T1_15_i_99 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_7_7,
   I1 => W_reg_6_7,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_5_7,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_4_7,
   O => T1_15_i_99_n_0
);
T1_19_i_10 : LUT3
  generic map(
   INIT => X"b8"
  )
 port map (
   I0 => f_reg_n_0_18,
   I1 => ROTR11_out_25,
   I2 => g_reg_n_0_18,
   O => T1_19_i_10_n_0
);
T1_19_i_101 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_31_11,
   I1 => W_reg_30_11,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_29_11,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_28_11,
   O => T1_19_i_101_n_0
);
T1_19_i_102 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_27_11,
   I1 => W_reg_26_11,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_25_11,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_24_11,
   O => T1_19_i_102_n_0
);
T1_19_i_103 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_19_11,
   I1 => W_reg_18_11,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_17_11,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_16_11,
   O => T1_19_i_103_n_0
);
T1_19_i_104 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_23_11,
   I1 => W_reg_22_11,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_21_11,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_20_11,
   O => T1_19_i_104_n_0
);
T1_19_i_105 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_3_11,
   I1 => W_reg_2_11,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_1_11,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_0_11,
   O => T1_19_i_105_n_0
);
T1_19_i_106 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_7_11,
   I1 => W_reg_6_11,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_5_11,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_4_11,
   O => T1_19_i_106_n_0
);
T1_19_i_107 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_11_11,
   I1 => W_reg_10_11,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_9_11,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_8_11,
   O => T1_19_i_107_n_0
);
T1_19_i_108 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_15_11,
   I1 => W_reg_14_11,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_13_11,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_12_11,
   O => T1_19_i_108_n_0
);
T1_19_i_11 : LUT3
  generic map(
   INIT => X"b8"
  )
 port map (
   I0 => f_reg_n_0_17,
   I1 => ROTR11_out_26,
   I2 => g_reg_n_0_17,
   O => T1_19_i_11_n_0
);
T1_19_i_12 : LUT3
  generic map(
   INIT => X"b8"
  )
 port map (
   I0 => f_reg_n_0_16,
   I1 => ROTR11_out_27,
   I2 => g_reg_n_0_16,
   O => T1_19_i_12_n_0
);
T1_19_i_14 : LUT3
  generic map(
   INIT => X"b8"
  )
 port map (
   I0 => f_reg_n_0_15,
   I1 => ROTR11_out_28,
   I2 => g_reg_n_0_15,
   O => T1_19_i_14_n_0
);
T1_19_i_15 : LUT3
  generic map(
   INIT => X"e8"
  )
 port map (
   I0 => g0_b14_n_0,
   I1 => T1_19_i_23_n_0,
   I2 => h_14,
   O => T1_19_i_15_n_0
);
T1_19_i_16 : LUT3
  generic map(
   INIT => X"e8"
  )
 port map (
   I0 => g0_b13_n_0,
   I1 => T1_19_i_24_n_0,
   I2 => h_13,
   O => T1_19_i_16_n_0
);
T1_19_i_17 : LUT3
  generic map(
   INIT => X"e8"
  )
 port map (
   I0 => g0_b12_n_0,
   I1 => T1_19_i_25_n_0,
   I2 => h_12,
   O => T1_19_i_17_n_0
);
T1_19_i_18 : LUT3
  generic map(
   INIT => X"e8"
  )
 port map (
   I0 => g0_b11_n_0,
   I1 => T1_19_i_26_n_0,
   I2 => h_11,
   O => T1_19_i_18_n_0
);
T1_19_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => g0_b15_n_0,
   I1 => T1_23_i_26_n_0,
   I2 => h_15,
   I3 => T1_19_i_15_n_0,
   O => T1_19_i_19_n_0
);
T1_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => ROTR11_out_32,
   I1 => ROTR11_out_19,
   I2 => ROTR11_out_14,
   I3 => T1_reg_23_i_13_n_5,
   I4 => T1_19_i_10_n_0,
   O => T1_19_i_2_n_0
);
T1_19_i_20 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => g0_b14_n_0,
   I1 => T1_19_i_23_n_0,
   I2 => h_14,
   I3 => T1_19_i_16_n_0,
   O => T1_19_i_20_n_0
);
T1_19_i_21 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => g0_b13_n_0,
   I1 => T1_19_i_24_n_0,
   I2 => h_13,
   I3 => T1_19_i_17_n_0,
   O => T1_19_i_21_n_0
);
T1_19_i_22 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => g0_b12_n_0,
   I1 => T1_19_i_25_n_0,
   I2 => h_12,
   I3 => T1_19_i_18_n_0,
   O => T1_19_i_22_n_0
);
T1_19_i_23 : LUT6
  generic map(
   INIT => X"505f505f30303f3f"
  )
 port map (
   I0 => T1_19_i_27_n_0,
   I1 => T1_19_i_28_n_0,
   I2 => HASH_02_COUNTER_5,
   I3 => T1_19_i_29_n_0,
   I4 => T1_19_i_30_n_0,
   I5 => HASH_02_COUNTER_4,
   O => T1_19_i_23_n_0
);
T1_19_i_24 : LUT6
  generic map(
   INIT => X"505f505f30303f3f"
  )
 port map (
   I0 => T1_19_i_31_n_0,
   I1 => T1_19_i_32_n_0,
   I2 => HASH_02_COUNTER_5,
   I3 => T1_19_i_33_n_0,
   I4 => T1_19_i_34_n_0,
   I5 => HASH_02_COUNTER_4,
   O => T1_19_i_24_n_0
);
T1_19_i_25 : LUT6
  generic map(
   INIT => X"303f303f50505f5f"
  )
 port map (
   I0 => T1_19_i_35_n_0,
   I1 => T1_19_i_36_n_0,
   I2 => HASH_02_COUNTER_5,
   I3 => T1_19_i_37_n_0,
   I4 => T1_19_i_38_n_0,
   I5 => HASH_02_COUNTER_4,
   O => T1_19_i_25_n_0
);
T1_19_i_26 : LUT6
  generic map(
   INIT => X"50505f5f3f303f30"
  )
 port map (
   I0 => T1_19_i_39_n_0,
   I1 => T1_19_i_40_n_0,
   I2 => HASH_02_COUNTER_5,
   I3 => T1_reg_19_i_41_n_0,
   I4 => T1_19_i_42_n_0,
   I5 => HASH_02_COUNTER_4,
   O => T1_19_i_26_n_0
);
T1_19_i_27 : LUT6
  generic map(
   INIT => X"303f5050303f5f5f"
  )
 port map (
   I0 => T1_19_i_43_n_0,
   I1 => T1_19_i_44_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_19_i_45_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_19_i_46_n_0,
   O => T1_19_i_27_n_0
);
T1_19_i_28 : LUT6
  generic map(
   INIT => X"3030505f3f3f505f"
  )
 port map (
   I0 => T1_19_i_47_n_0,
   I1 => T1_19_i_48_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_19_i_49_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_19_i_50_n_0,
   O => T1_19_i_28_n_0
);
T1_19_i_29 : LUT6
  generic map(
   INIT => X"3030505f3f3f505f"
  )
 port map (
   I0 => T1_19_i_51_n_0,
   I1 => T1_19_i_52_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_19_i_53_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_19_i_54_n_0,
   O => T1_19_i_29_n_0
);
T1_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => ROTR11_out_15,
   I1 => ROTR11_out_20,
   I2 => ROTR11_out_1,
   I3 => T1_reg_23_i_13_n_6,
   I4 => T1_19_i_11_n_0,
   O => T1_19_i_3_n_0
);
T1_19_i_30 : LUT6
  generic map(
   INIT => X"303f5050303f5f5f"
  )
 port map (
   I0 => T1_19_i_55_n_0,
   I1 => T1_19_i_56_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_19_i_57_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_19_i_58_n_0,
   O => T1_19_i_30_n_0
);
T1_19_i_31 : LUT6
  generic map(
   INIT => X"5050303f5f5f303f"
  )
 port map (
   I0 => T1_19_i_59_n_0,
   I1 => T1_19_i_60_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_19_i_61_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_19_i_62_n_0,
   O => T1_19_i_31_n_0
);
T1_19_i_32 : LUT6
  generic map(
   INIT => X"505f3030505f3f3f"
  )
 port map (
   I0 => T1_19_i_63_n_0,
   I1 => T1_19_i_64_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_19_i_65_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_19_i_66_n_0,
   O => T1_19_i_32_n_0
);
T1_19_i_33 : LUT6
  generic map(
   INIT => X"5050303f5f5f303f"
  )
 port map (
   I0 => T1_19_i_67_n_0,
   I1 => T1_19_i_68_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_19_i_69_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_19_i_70_n_0,
   O => T1_19_i_33_n_0
);
T1_19_i_34 : LUT6
  generic map(
   INIT => X"505f3030505f3f3f"
  )
 port map (
   I0 => T1_19_i_71_n_0,
   I1 => T1_19_i_72_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_19_i_73_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_19_i_74_n_0,
   O => T1_19_i_34_n_0
);
T1_19_i_35 : LUT6
  generic map(
   INIT => X"5050303f5f5f303f"
  )
 port map (
   I0 => T1_19_i_75_n_0,
   I1 => T1_19_i_76_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_19_i_77_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_19_i_78_n_0,
   O => T1_19_i_35_n_0
);
T1_19_i_36 : LUT6
  generic map(
   INIT => X"505f3030505f3f3f"
  )
 port map (
   I0 => T1_19_i_79_n_0,
   I1 => T1_19_i_80_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_19_i_81_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_19_i_82_n_0,
   O => T1_19_i_36_n_0
);
T1_19_i_37 : LUT6
  generic map(
   INIT => X"5050303f5f5f303f"
  )
 port map (
   I0 => T1_19_i_83_n_0,
   I1 => T1_19_i_84_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_19_i_85_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_19_i_86_n_0,
   O => T1_19_i_37_n_0
);
T1_19_i_38 : LUT6
  generic map(
   INIT => X"303f5050303f5f5f"
  )
 port map (
   I0 => T1_19_i_87_n_0,
   I1 => T1_19_i_88_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_19_i_89_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_19_i_90_n_0,
   O => T1_19_i_38_n_0
);
T1_19_i_39 : LUT6
  generic map(
   INIT => X"505f3030505f3f3f"
  )
 port map (
   I0 => T1_19_i_91_n_0,
   I1 => T1_19_i_92_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_19_i_93_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_19_i_94_n_0,
   O => T1_19_i_39_n_0
);
T1_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => ROTR11_out_16,
   I1 => ROTR11_out_21,
   I2 => ROTR11_out_2,
   I3 => T1_reg_23_i_13_n_7,
   I4 => T1_19_i_12_n_0,
   O => T1_19_i_4_n_0
);
T1_19_i_40 : LUT6
  generic map(
   INIT => X"5050303f5f5f303f"
  )
 port map (
   I0 => T1_19_i_95_n_0,
   I1 => T1_19_i_96_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_19_i_97_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_19_i_98_n_0,
   O => T1_19_i_40_n_0
);
T1_19_i_42 : LUT6
  generic map(
   INIT => X"5050303f5f5f303f"
  )
 port map (
   I0 => T1_19_i_101_n_0,
   I1 => T1_19_i_102_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_19_i_103_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_19_i_104_n_0,
   O => T1_19_i_42_n_0
);
T1_19_i_43 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_59_14,
   I1 => W_reg_58_14,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_57_14,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_56_14,
   O => T1_19_i_43_n_0
);
T1_19_i_44 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_63_14,
   I1 => W_reg_62_14,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_61_14,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_60_14,
   O => T1_19_i_44_n_0
);
T1_19_i_45 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_55_14,
   I1 => W_reg_54_14,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_53_14,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_52_14,
   O => T1_19_i_45_n_0
);
T1_19_i_46 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_51_14,
   I1 => W_reg_50_14,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_49_14,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_48_14,
   O => T1_19_i_46_n_0
);
T1_19_i_47 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_43_14,
   I1 => W_reg_42_14,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_41_14,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_40_14,
   O => T1_19_i_47_n_0
);
T1_19_i_48 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_47_14,
   I1 => W_reg_46_14,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_45_14,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_44_14,
   O => T1_19_i_48_n_0
);
T1_19_i_49 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_35_14,
   I1 => W_reg_34_14,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_33_14,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_32_14,
   O => T1_19_i_49_n_0
);
T1_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => ROTR11_out_17,
   I1 => ROTR11_out_22,
   I2 => ROTR11_out_3,
   I3 => T1_reg_19_i_13_n_4,
   I4 => T1_19_i_14_n_0,
   O => T1_19_i_5_n_0
);
T1_19_i_50 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_39_14,
   I1 => W_reg_38_14,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_37_14,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_36_14,
   O => T1_19_i_50_n_0
);
T1_19_i_51 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_27_14,
   I1 => W_reg_26_14,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_25_14,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_24_14,
   O => T1_19_i_51_n_0
);
T1_19_i_52 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_31_14,
   I1 => W_reg_30_14,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_29_14,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_28_14,
   O => T1_19_i_52_n_0
);
T1_19_i_53 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_19_14,
   I1 => W_reg_18_14,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_17_14,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_16_14,
   O => T1_19_i_53_n_0
);
T1_19_i_54 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_23_14,
   I1 => W_reg_22_14,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_21_14,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_20_14,
   O => T1_19_i_54_n_0
);
T1_19_i_55 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_11_14,
   I1 => W_reg_10_14,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_9_14,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_8_14,
   O => T1_19_i_55_n_0
);
T1_19_i_56 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_15_14,
   I1 => W_reg_14_14,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_13_14,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_12_14,
   O => T1_19_i_56_n_0
);
T1_19_i_57 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_7_14,
   I1 => W_reg_6_14,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_5_14,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_4_14,
   O => T1_19_i_57_n_0
);
T1_19_i_58 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_3_14,
   I1 => W_reg_2_14,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_1_14,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_0_14,
   O => T1_19_i_58_n_0
);
T1_19_i_59 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_63_13,
   I1 => W_reg_62_13,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_61_13,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_60_13,
   O => T1_19_i_59_n_0
);
T1_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => T1_19_i_2_n_0,
   I1 => ROTR11_out_18,
   I2 => ROTR11_out_13,
   I3 => ROTR11_out_31,
   I4 => T1_reg_23_i_13_n_4,
   I5 => T1_23_i_14_n_0,
   O => T1_19_i_6_n_0
);
T1_19_i_60 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_59_13,
   I1 => W_reg_58_13,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_57_13,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_56_13,
   O => T1_19_i_60_n_0
);
T1_19_i_61 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_51_13,
   I1 => W_reg_50_13,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_49_13,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_48_13,
   O => T1_19_i_61_n_0
);
T1_19_i_62 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_55_13,
   I1 => W_reg_54_13,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_53_13,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_52_13,
   O => T1_19_i_62_n_0
);
T1_19_i_63 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_47_13,
   I1 => W_reg_46_13,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_45_13,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_44_13,
   O => T1_19_i_63_n_0
);
T1_19_i_64 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_43_13,
   I1 => W_reg_42_13,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_41_13,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_40_13,
   O => T1_19_i_64_n_0
);
T1_19_i_65 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_39_13,
   I1 => W_reg_38_13,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_37_13,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_36_13,
   O => T1_19_i_65_n_0
);
T1_19_i_66 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_35_13,
   I1 => W_reg_34_13,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_33_13,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_32_13,
   O => T1_19_i_66_n_0
);
T1_19_i_67 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_31_13,
   I1 => W_reg_30_13,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_29_13,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_28_13,
   O => T1_19_i_67_n_0
);
T1_19_i_68 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_27_13,
   I1 => W_reg_26_13,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_25_13,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_24_13,
   O => T1_19_i_68_n_0
);
T1_19_i_69 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_19_13,
   I1 => W_reg_18_13,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_17_13,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_16_13,
   O => T1_19_i_69_n_0
);
T1_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => T1_19_i_3_n_0,
   I1 => ROTR11_out_32,
   I2 => ROTR11_out_19,
   I3 => ROTR11_out_14,
   I4 => T1_reg_23_i_13_n_5,
   I5 => T1_19_i_10_n_0,
   O => T1_19_i_7_n_0
);
T1_19_i_70 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_23_13,
   I1 => W_reg_22_13,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_21_13,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_20_13,
   O => T1_19_i_70_n_0
);
T1_19_i_71 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_15_13,
   I1 => W_reg_14_13,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_13_13,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_12_13,
   O => T1_19_i_71_n_0
);
T1_19_i_72 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_11_13,
   I1 => W_reg_10_13,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_9_13,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_8_13,
   O => T1_19_i_72_n_0
);
T1_19_i_73 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_7_13,
   I1 => W_reg_6_13,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_5_13,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_4_13,
   O => T1_19_i_73_n_0
);
T1_19_i_74 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_3_13,
   I1 => W_reg_2_13,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_1_13,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_0_13,
   O => T1_19_i_74_n_0
);
T1_19_i_75 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_47_12,
   I1 => W_reg_46_12,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_45_12,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_44_12,
   O => T1_19_i_75_n_0
);
T1_19_i_76 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_43_12,
   I1 => W_reg_42_12,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_41_12,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_40_12,
   O => T1_19_i_76_n_0
);
T1_19_i_77 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_35_12,
   I1 => W_reg_34_12,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_33_12,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_32_12,
   O => T1_19_i_77_n_0
);
T1_19_i_78 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_39_12,
   I1 => W_reg_38_12,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_37_12,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_36_12,
   O => T1_19_i_78_n_0
);
T1_19_i_79 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_63_12,
   I1 => W_reg_62_12,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_61_12,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_60_12,
   O => T1_19_i_79_n_0
);
T1_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => T1_19_i_4_n_0,
   I1 => T1_reg_23_i_13_n_6,
   I2 => T1_19_i_11_n_0,
   I3 => ROTR11_out_15,
   I4 => ROTR11_out_20,
   I5 => ROTR11_out_1,
   O => T1_19_i_8_n_0
);
T1_19_i_80 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_59_12,
   I1 => W_reg_58_12,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_57_12,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_56_12,
   O => T1_19_i_80_n_0
);
T1_19_i_81 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_55_12,
   I1 => W_reg_54_12,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_53_12,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_52_12,
   O => T1_19_i_81_n_0
);
T1_19_i_82 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_51_12,
   I1 => W_reg_50_12,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_49_12,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_48_12,
   O => T1_19_i_82_n_0
);
T1_19_i_83 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_31_12,
   I1 => W_reg_30_12,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_29_12,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_28_12,
   O => T1_19_i_83_n_0
);
T1_19_i_84 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_27_12,
   I1 => W_reg_26_12,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_25_12,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_24_12,
   O => T1_19_i_84_n_0
);
T1_19_i_85 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_19_12,
   I1 => W_reg_18_12,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_17_12,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_16_12,
   O => T1_19_i_85_n_0
);
T1_19_i_86 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_23_12,
   I1 => W_reg_22_12,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_21_12,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_20_12,
   O => T1_19_i_86_n_0
);
T1_19_i_87 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_11_12,
   I1 => W_reg_10_12,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_9_12,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_8_12,
   O => T1_19_i_87_n_0
);
T1_19_i_88 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_15_12,
   I1 => W_reg_14_12,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_13_12,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_12_12,
   O => T1_19_i_88_n_0
);
T1_19_i_89 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_7_12,
   I1 => W_reg_6_12,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_5_12,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_4_12,
   O => T1_19_i_89_n_0
);
T1_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => T1_19_i_5_n_0,
   I1 => ROTR11_out_16,
   I2 => ROTR11_out_21,
   I3 => ROTR11_out_2,
   I4 => T1_reg_23_i_13_n_7,
   I5 => T1_19_i_12_n_0,
   O => T1_19_i_9_n_0
);
T1_19_i_90 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_3_12,
   I1 => W_reg_2_12,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_1_12,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_0_12,
   O => T1_19_i_90_n_0
);
T1_19_i_91 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_63_11,
   I1 => W_reg_62_11,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_61_11,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_60_11,
   O => T1_19_i_91_n_0
);
T1_19_i_92 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_59_11,
   I1 => W_reg_58_11,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_57_11,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_56_11,
   O => T1_19_i_92_n_0
);
T1_19_i_93 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_55_11,
   I1 => W_reg_54_11,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_53_11,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_52_11,
   O => T1_19_i_93_n_0
);
T1_19_i_94 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_51_11,
   I1 => W_reg_50_11,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_49_11,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_48_11,
   O => T1_19_i_94_n_0
);
T1_19_i_95 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_47_11,
   I1 => W_reg_46_11,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_45_11,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_44_11,
   O => T1_19_i_95_n_0
);
T1_19_i_96 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_43_11,
   I1 => W_reg_42_11,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_41_11,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_40_11,
   O => T1_19_i_96_n_0
);
T1_19_i_97 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_35_11,
   I1 => W_reg_34_11,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_33_11,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_32_11,
   O => T1_19_i_97_n_0
);
T1_19_i_98 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_39_11,
   I1 => W_reg_38_11,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_37_11,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_36_11,
   O => T1_19_i_98_n_0
);
T1_23_i_10 : LUT3
  generic map(
   INIT => X"b8"
  )
 port map (
   I0 => f_reg_n_0_22,
   I1 => ROTR11_out_21,
   I2 => g_reg_n_0_22,
   O => T1_23_i_10_n_0
);
T1_23_i_100 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_23_15,
   I1 => W_reg_22_15,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_21_15,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_20_15,
   O => T1_23_i_100_n_0
);
T1_23_i_101 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_15_15,
   I1 => W_reg_14_15,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_13_15,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_12_15,
   O => T1_23_i_101_n_0
);
T1_23_i_102 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_11_15,
   I1 => W_reg_10_15,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_9_15,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_8_15,
   O => T1_23_i_102_n_0
);
T1_23_i_103 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_3_15,
   I1 => W_reg_2_15,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_1_15,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_0_15,
   O => T1_23_i_103_n_0
);
T1_23_i_104 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_7_15,
   I1 => W_reg_6_15,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_5_15,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_4_15,
   O => T1_23_i_104_n_0
);
T1_23_i_105 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_35_15,
   I1 => W_reg_34_15,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_33_15,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_32_15,
   O => T1_23_i_105_n_0
);
T1_23_i_106 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_39_15,
   I1 => W_reg_38_15,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_37_15,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_36_15,
   O => T1_23_i_106_n_0
);
T1_23_i_107 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_43_15,
   I1 => W_reg_42_15,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_41_15,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_40_15,
   O => T1_23_i_107_n_0
);
T1_23_i_108 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_47_15,
   I1 => W_reg_46_15,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_45_15,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_44_15,
   O => T1_23_i_108_n_0
);
T1_23_i_11 : LUT3
  generic map(
   INIT => X"b8"
  )
 port map (
   I0 => f_reg_n_0_21,
   I1 => ROTR11_out_22,
   I2 => g_reg_n_0_21,
   O => T1_23_i_11_n_0
);
T1_23_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => ROTR11_out_12,
   I1 => ROTR11_out_30,
   I2 => ROTR11_out_17,
   O => T1_23_i_12_n_0
);
T1_23_i_14 : LUT3
  generic map(
   INIT => X"b8"
  )
 port map (
   I0 => f_reg_n_0_19,
   I1 => ROTR11_out_24,
   I2 => g_reg_n_0_19,
   O => T1_23_i_14_n_0
);
T1_23_i_15 : LUT3
  generic map(
   INIT => X"e8"
  )
 port map (
   I0 => g0_b18_n_0,
   I1 => T1_23_i_23_n_0,
   I2 => h_18,
   O => T1_23_i_15_n_0
);
T1_23_i_16 : LUT3
  generic map(
   INIT => X"e8"
  )
 port map (
   I0 => g0_b17_n_0,
   I1 => T1_23_i_24_n_0,
   I2 => h_17,
   O => T1_23_i_16_n_0
);
T1_23_i_17 : LUT3
  generic map(
   INIT => X"e8"
  )
 port map (
   I0 => g0_b16_n_0,
   I1 => T1_23_i_25_n_0,
   I2 => h_16,
   O => T1_23_i_17_n_0
);
T1_23_i_18 : LUT3
  generic map(
   INIT => X"e8"
  )
 port map (
   I0 => g0_b15_n_0,
   I1 => T1_23_i_26_n_0,
   I2 => h_15,
   O => T1_23_i_18_n_0
);
T1_23_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => g0_b19_n_0,
   I1 => T1_27_i_26_n_0,
   I2 => h_19,
   I3 => T1_23_i_15_n_0,
   O => T1_23_i_19_n_0
);
T1_23_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => ROTR11_out_15,
   I1 => ROTR11_out_10,
   I2 => ROTR11_out_28,
   I3 => T1_reg_27_i_13_n_5,
   I4 => T1_23_i_10_n_0,
   O => T1_23_i_2_n_0
);
T1_23_i_20 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => g0_b18_n_0,
   I1 => T1_23_i_23_n_0,
   I2 => h_18,
   I3 => T1_23_i_16_n_0,
   O => T1_23_i_20_n_0
);
T1_23_i_21 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => g0_b17_n_0,
   I1 => T1_23_i_24_n_0,
   I2 => h_17,
   I3 => T1_23_i_17_n_0,
   O => T1_23_i_21_n_0
);
T1_23_i_22 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => g0_b16_n_0,
   I1 => T1_23_i_25_n_0,
   I2 => h_16,
   I3 => T1_23_i_18_n_0,
   O => T1_23_i_22_n_0
);
T1_23_i_23 : LUT6
  generic map(
   INIT => X"505f505f30303f3f"
  )
 port map (
   I0 => T1_23_i_27_n_0,
   I1 => T1_23_i_28_n_0,
   I2 => HASH_02_COUNTER_5,
   I3 => T1_23_i_29_n_0,
   I4 => T1_23_i_30_n_0,
   I5 => HASH_02_COUNTER_4,
   O => T1_23_i_23_n_0
);
T1_23_i_24 : LUT6
  generic map(
   INIT => X"505f505f30303f3f"
  )
 port map (
   I0 => T1_23_i_31_n_0,
   I1 => T1_23_i_32_n_0,
   I2 => HASH_02_COUNTER_5,
   I3 => T1_23_i_33_n_0,
   I4 => T1_23_i_34_n_0,
   I5 => HASH_02_COUNTER_4,
   O => T1_23_i_24_n_0
);
T1_23_i_25 : LUT6
  generic map(
   INIT => X"505f505f30303f3f"
  )
 port map (
   I0 => T1_23_i_35_n_0,
   I1 => T1_23_i_36_n_0,
   I2 => HASH_02_COUNTER_5,
   I3 => T1_23_i_37_n_0,
   I4 => T1_23_i_38_n_0,
   I5 => HASH_02_COUNTER_4,
   O => T1_23_i_25_n_0
);
T1_23_i_26 : LUT6
  generic map(
   INIT => X"505f505fc0c0cfcf"
  )
 port map (
   I0 => T1_23_i_39_n_0,
   I1 => T1_reg_23_i_40_n_0,
   I2 => HASH_02_COUNTER_5,
   I3 => T1_23_i_41_n_0,
   I4 => T1_23_i_42_n_0,
   I5 => HASH_02_COUNTER_4,
   O => T1_23_i_26_n_0
);
T1_23_i_27 : LUT6
  generic map(
   INIT => X"303f5050303f5f5f"
  )
 port map (
   I0 => T1_23_i_43_n_0,
   I1 => T1_23_i_44_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_23_i_45_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_23_i_46_n_0,
   O => T1_23_i_27_n_0
);
T1_23_i_28 : LUT6
  generic map(
   INIT => X"05f5030305f5f3f3"
  )
 port map (
   I0 => T1_23_i_47_n_0,
   I1 => T1_23_i_48_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_23_i_49_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_23_i_50_n_0,
   O => T1_23_i_28_n_0
);
T1_23_i_29 : LUT6
  generic map(
   INIT => X"5050303f5f5f303f"
  )
 port map (
   I0 => T1_23_i_51_n_0,
   I1 => T1_23_i_52_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_23_i_53_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_23_i_54_n_0,
   O => T1_23_i_29_n_0
);
T1_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => ROTR11_out_16,
   I1 => ROTR11_out_11,
   I2 => ROTR11_out_29,
   I3 => T1_reg_27_i_13_n_6,
   I4 => T1_23_i_11_n_0,
   O => T1_23_i_3_n_0
);
T1_23_i_30 : LUT6
  generic map(
   INIT => X"303f5050303f5f5f"
  )
 port map (
   I0 => T1_23_i_55_n_0,
   I1 => T1_23_i_56_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_23_i_57_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_23_i_58_n_0,
   O => T1_23_i_30_n_0
);
T1_23_i_31 : LUT6
  generic map(
   INIT => X"5050303f5f5f303f"
  )
 port map (
   I0 => T1_23_i_59_n_0,
   I1 => T1_23_i_60_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_23_i_61_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_23_i_62_n_0,
   O => T1_23_i_31_n_0
);
T1_23_i_32 : LUT6
  generic map(
   INIT => X"5050303f5f5f303f"
  )
 port map (
   I0 => T1_23_i_63_n_0,
   I1 => T1_23_i_64_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_23_i_65_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_23_i_66_n_0,
   O => T1_23_i_32_n_0
);
T1_23_i_33 : LUT6
  generic map(
   INIT => X"3030505f3f3f505f"
  )
 port map (
   I0 => T1_23_i_67_n_0,
   I1 => T1_23_i_68_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_23_i_69_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_23_i_70_n_0,
   O => T1_23_i_33_n_0
);
T1_23_i_34 : LUT6
  generic map(
   INIT => X"303f5050303f5f5f"
  )
 port map (
   I0 => T1_23_i_71_n_0,
   I1 => T1_23_i_72_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_23_i_73_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_23_i_74_n_0,
   O => T1_23_i_34_n_0
);
T1_23_i_35 : LUT6
  generic map(
   INIT => X"3030505f3f3f505f"
  )
 port map (
   I0 => T1_23_i_75_n_0,
   I1 => T1_23_i_76_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_23_i_77_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_23_i_78_n_0,
   O => T1_23_i_35_n_0
);
T1_23_i_36 : LUT6
  generic map(
   INIT => X"303f5050303f5f5f"
  )
 port map (
   I0 => T1_23_i_79_n_0,
   I1 => T1_23_i_80_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_23_i_81_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_23_i_82_n_0,
   O => T1_23_i_36_n_0
);
T1_23_i_37 : LUT6
  generic map(
   INIT => X"303f5050303f5f5f"
  )
 port map (
   I0 => T1_23_i_83_n_0,
   I1 => T1_23_i_84_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_23_i_85_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_23_i_86_n_0,
   O => T1_23_i_37_n_0
);
T1_23_i_38 : LUT6
  generic map(
   INIT => X"5050303f5f5f303f"
  )
 port map (
   I0 => T1_23_i_87_n_0,
   I1 => T1_23_i_88_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_23_i_89_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_23_i_90_n_0,
   O => T1_23_i_38_n_0
);
T1_23_i_39 : LUT6
  generic map(
   INIT => X"303f5050303f5f5f"
  )
 port map (
   I0 => T1_23_i_91_n_0,
   I1 => T1_23_i_92_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_23_i_93_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_23_i_94_n_0,
   O => T1_23_i_39_n_0
);
T1_23_i_4 : LUT5
  generic map(
   INIT => X"ffb8b800"
  )
 port map (
   I0 => f_reg_n_0_20,
   I1 => ROTR11_out_23,
   I2 => g_reg_n_0_20,
   I3 => T1_reg_27_i_13_n_7,
   I4 => T1_23_i_12_n_0,
   O => T1_23_i_4_n_0
);
T1_23_i_41 : LUT6
  generic map(
   INIT => X"3030505f3f3f505f"
  )
 port map (
   I0 => T1_23_i_97_n_0,
   I1 => T1_23_i_98_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_23_i_99_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_23_i_100_n_0,
   O => T1_23_i_41_n_0
);
T1_23_i_42 : LUT6
  generic map(
   INIT => X"5050303f5f5f303f"
  )
 port map (
   I0 => T1_23_i_101_n_0,
   I1 => T1_23_i_102_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_23_i_103_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_23_i_104_n_0,
   O => T1_23_i_42_n_0
);
T1_23_i_43 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_59_18,
   I1 => W_reg_58_18,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_57_18,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_56_18,
   O => T1_23_i_43_n_0
);
T1_23_i_44 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_63_18,
   I1 => W_reg_62_18,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_61_18,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_60_18,
   O => T1_23_i_44_n_0
);
T1_23_i_45 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_55_18,
   I1 => W_reg_54_18,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_53_18,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_52_18,
   O => T1_23_i_45_n_0
);
T1_23_i_46 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_51_18,
   I1 => W_reg_50_18,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_49_18,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_48_18,
   O => T1_23_i_46_n_0
);
T1_23_i_47 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_39_18,
   I1 => W_reg_38_18,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_37_18,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_36_18,
   O => T1_23_i_47_n_0
);
T1_23_i_48 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_35_18,
   I1 => W_reg_34_18,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_33_18,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_32_18,
   O => T1_23_i_48_n_0
);
T1_23_i_49 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_47_18,
   I1 => W_reg_46_18,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_45_18,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_44_18,
   O => T1_23_i_49_n_0
);
T1_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => ROTR11_out_18,
   I1 => ROTR11_out_13,
   I2 => ROTR11_out_31,
   I3 => T1_reg_23_i_13_n_4,
   I4 => T1_23_i_14_n_0,
   O => T1_23_i_5_n_0
);
T1_23_i_50 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_43_18,
   I1 => W_reg_42_18,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_41_18,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_40_18,
   O => T1_23_i_50_n_0
);
T1_23_i_51 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_31_18,
   I1 => W_reg_30_18,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_29_18,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_28_18,
   O => T1_23_i_51_n_0
);
T1_23_i_52 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_27_18,
   I1 => W_reg_26_18,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_25_18,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_24_18,
   O => T1_23_i_52_n_0
);
T1_23_i_53 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_19_18,
   I1 => W_reg_18_18,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_17_18,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_16_18,
   O => T1_23_i_53_n_0
);
T1_23_i_54 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_23_18,
   I1 => W_reg_22_18,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_21_18,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_20_18,
   O => T1_23_i_54_n_0
);
T1_23_i_55 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_11_18,
   I1 => W_reg_10_18,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_9_18,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_8_18,
   O => T1_23_i_55_n_0
);
T1_23_i_56 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_15_18,
   I1 => W_reg_14_18,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_13_18,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_12_18,
   O => T1_23_i_56_n_0
);
T1_23_i_57 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_7_18,
   I1 => W_reg_6_18,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_5_18,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_4_18,
   O => T1_23_i_57_n_0
);
T1_23_i_58 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_3_18,
   I1 => W_reg_2_18,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_1_18,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_0_18,
   O => T1_23_i_58_n_0
);
T1_23_i_59 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_63_17,
   I1 => W_reg_62_17,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_61_17,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_60_17,
   O => T1_23_i_59_n_0
);
T1_23_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => T1_23_i_2_n_0,
   I1 => ROTR11_out_14,
   I2 => ROTR11_out_9,
   I3 => ROTR11_out_27,
   I4 => T1_reg_27_i_13_n_4,
   I5 => T1_27_i_14_n_0,
   O => T1_23_i_6_n_0
);
T1_23_i_60 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_59_17,
   I1 => W_reg_58_17,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_57_17,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_56_17,
   O => T1_23_i_60_n_0
);
T1_23_i_61 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_51_17,
   I1 => W_reg_50_17,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_49_17,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_48_17,
   O => T1_23_i_61_n_0
);
T1_23_i_62 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_55_17,
   I1 => W_reg_54_17,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_53_17,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_52_17,
   O => T1_23_i_62_n_0
);
T1_23_i_63 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_47_17,
   I1 => W_reg_46_17,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_45_17,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_44_17,
   O => T1_23_i_63_n_0
);
T1_23_i_64 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_43_17,
   I1 => W_reg_42_17,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_41_17,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_40_17,
   O => T1_23_i_64_n_0
);
T1_23_i_65 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_35_17,
   I1 => W_reg_34_17,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_33_17,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_32_17,
   O => T1_23_i_65_n_0
);
T1_23_i_66 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_39_17,
   I1 => W_reg_38_17,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_37_17,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_36_17,
   O => T1_23_i_66_n_0
);
T1_23_i_67 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_27_17,
   I1 => W_reg_26_17,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_25_17,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_24_17,
   O => T1_23_i_67_n_0
);
T1_23_i_68 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_31_17,
   I1 => W_reg_30_17,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_29_17,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_28_17,
   O => T1_23_i_68_n_0
);
T1_23_i_69 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_19_17,
   I1 => W_reg_18_17,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_17_17,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_16_17,
   O => T1_23_i_69_n_0
);
T1_23_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => T1_23_i_3_n_0,
   I1 => T1_reg_27_i_13_n_5,
   I2 => T1_23_i_10_n_0,
   I3 => ROTR11_out_15,
   I4 => ROTR11_out_10,
   I5 => ROTR11_out_28,
   O => T1_23_i_7_n_0
);
T1_23_i_70 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_23_17,
   I1 => W_reg_22_17,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_21_17,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_20_17,
   O => T1_23_i_70_n_0
);
T1_23_i_71 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_11_17,
   I1 => W_reg_10_17,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_9_17,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_8_17,
   O => T1_23_i_71_n_0
);
T1_23_i_72 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_15_17,
   I1 => W_reg_14_17,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_13_17,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_12_17,
   O => T1_23_i_72_n_0
);
T1_23_i_73 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_7_17,
   I1 => W_reg_6_17,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_5_17,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_4_17,
   O => T1_23_i_73_n_0
);
T1_23_i_74 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_3_17,
   I1 => W_reg_2_17,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_1_17,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_0_17,
   O => T1_23_i_74_n_0
);
T1_23_i_75 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_59_16,
   I1 => W_reg_58_16,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_57_16,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_56_16,
   O => T1_23_i_75_n_0
);
T1_23_i_76 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_63_16,
   I1 => W_reg_62_16,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_61_16,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_60_16,
   O => T1_23_i_76_n_0
);
T1_23_i_77 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_51_16,
   I1 => W_reg_50_16,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_49_16,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_48_16,
   O => T1_23_i_77_n_0
);
T1_23_i_78 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_55_16,
   I1 => W_reg_54_16,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_53_16,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_52_16,
   O => T1_23_i_78_n_0
);
T1_23_i_79 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_43_16,
   I1 => W_reg_42_16,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_41_16,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_40_16,
   O => T1_23_i_79_n_0
);
T1_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => T1_23_i_4_n_0,
   I1 => T1_reg_27_i_13_n_6,
   I2 => T1_23_i_11_n_0,
   I3 => ROTR11_out_16,
   I4 => ROTR11_out_11,
   I5 => ROTR11_out_29,
   O => T1_23_i_8_n_0
);
T1_23_i_80 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_47_16,
   I1 => W_reg_46_16,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_45_16,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_44_16,
   O => T1_23_i_80_n_0
);
T1_23_i_81 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_39_16,
   I1 => W_reg_38_16,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_37_16,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_36_16,
   O => T1_23_i_81_n_0
);
T1_23_i_82 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_35_16,
   I1 => W_reg_34_16,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_33_16,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_32_16,
   O => T1_23_i_82_n_0
);
T1_23_i_83 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_27_16,
   I1 => W_reg_26_16,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_25_16,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_24_16,
   O => T1_23_i_83_n_0
);
T1_23_i_84 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_31_16,
   I1 => W_reg_30_16,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_29_16,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_28_16,
   O => T1_23_i_84_n_0
);
T1_23_i_85 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_23_16,
   I1 => W_reg_22_16,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_21_16,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_20_16,
   O => T1_23_i_85_n_0
);
T1_23_i_86 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_19_16,
   I1 => W_reg_18_16,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_17_16,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_16_16,
   O => T1_23_i_86_n_0
);
T1_23_i_87 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_15_16,
   I1 => W_reg_14_16,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_13_16,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_12_16,
   O => T1_23_i_87_n_0
);
T1_23_i_88 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_11_16,
   I1 => W_reg_10_16,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_9_16,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_8_16,
   O => T1_23_i_88_n_0
);
T1_23_i_89 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_3_16,
   I1 => W_reg_2_16,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_1_16,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_0_16,
   O => T1_23_i_89_n_0
);
T1_23_i_9 : LUT6
  generic map(
   INIT => X"656a9a959a95656a"
  )
 port map (
   I0 => T1_23_i_5_n_0,
   I1 => f_reg_n_0_20,
   I2 => ROTR11_out_23,
   I3 => g_reg_n_0_20,
   I4 => T1_reg_27_i_13_n_7,
   I5 => T1_23_i_12_n_0,
   O => T1_23_i_9_n_0
);
T1_23_i_90 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_7_16,
   I1 => W_reg_6_16,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_5_16,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_4_16,
   O => T1_23_i_90_n_0
);
T1_23_i_91 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_59_15,
   I1 => W_reg_58_15,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_57_15,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_56_15,
   O => T1_23_i_91_n_0
);
T1_23_i_92 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_63_15,
   I1 => W_reg_62_15,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_61_15,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_60_15,
   O => T1_23_i_92_n_0
);
T1_23_i_93 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_55_15,
   I1 => W_reg_54_15,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_53_15,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_52_15,
   O => T1_23_i_93_n_0
);
T1_23_i_94 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_51_15,
   I1 => W_reg_50_15,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_49_15,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_48_15,
   O => T1_23_i_94_n_0
);
T1_23_i_97 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_27_15,
   I1 => W_reg_26_15,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_25_15,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_24_15,
   O => T1_23_i_97_n_0
);
T1_23_i_98 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_31_15,
   I1 => W_reg_30_15,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_29_15,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_28_15,
   O => T1_23_i_98_n_0
);
T1_23_i_99 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_19_15,
   I1 => W_reg_18_15,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_17_15,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_16_15,
   O => T1_23_i_99_n_0
);
T1_27_i_10 : LUT3
  generic map(
   INIT => X"b8"
  )
 port map (
   I0 => f_reg_n_0_26,
   I1 => ROTR11_out_17,
   I2 => g_reg_n_0_26,
   O => T1_27_i_10_n_0
);
T1_27_i_100 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_19_19,
   I1 => W_reg_18_19,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_17_19,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_16_19,
   O => T1_27_i_100_n_0
);
T1_27_i_101 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_15_19,
   I1 => W_reg_14_19,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_13_19,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_12_19,
   O => T1_27_i_101_n_0
);
T1_27_i_102 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_11_19,
   I1 => W_reg_10_19,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_9_19,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_8_19,
   O => T1_27_i_102_n_0
);
T1_27_i_103 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_7_19,
   I1 => W_reg_6_19,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_5_19,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_4_19,
   O => T1_27_i_103_n_0
);
T1_27_i_104 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_3_19,
   I1 => W_reg_2_19,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_1_19,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_0_19,
   O => T1_27_i_104_n_0
);
T1_27_i_105 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_35_22,
   I1 => W_reg_34_22,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_33_22,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_32_22,
   O => T1_27_i_105_n_0
);
T1_27_i_106 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_39_22,
   I1 => W_reg_38_22,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_37_22,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_36_22,
   O => T1_27_i_106_n_0
);
T1_27_i_107 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_43_22,
   I1 => W_reg_42_22,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_41_22,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_40_22,
   O => T1_27_i_107_n_0
);
T1_27_i_108 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_47_22,
   I1 => W_reg_46_22,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_45_22,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_44_22,
   O => T1_27_i_108_n_0
);
T1_27_i_11 : LUT3
  generic map(
   INIT => X"b8"
  )
 port map (
   I0 => f_reg_n_0_25,
   I1 => ROTR11_out_18,
   I2 => g_reg_n_0_25,
   O => T1_27_i_11_n_0
);
T1_27_i_12 : LUT3
  generic map(
   INIT => X"b8"
  )
 port map (
   I0 => f_reg_n_0_24,
   I1 => ROTR11_out_19,
   I2 => g_reg_n_0_24,
   O => T1_27_i_12_n_0
);
T1_27_i_14 : LUT3
  generic map(
   INIT => X"b8"
  )
 port map (
   I0 => f_reg_n_0_23,
   I1 => ROTR11_out_20,
   I2 => g_reg_n_0_23,
   O => T1_27_i_14_n_0
);
T1_27_i_15 : LUT3
  generic map(
   INIT => X"e8"
  )
 port map (
   I0 => g0_b22_n_0,
   I1 => T1_27_i_23_n_0,
   I2 => h_22,
   O => T1_27_i_15_n_0
);
T1_27_i_16 : LUT3
  generic map(
   INIT => X"e8"
  )
 port map (
   I0 => g0_b21_n_0,
   I1 => T1_27_i_24_n_0,
   I2 => h_21,
   O => T1_27_i_16_n_0
);
T1_27_i_17 : LUT3
  generic map(
   INIT => X"e8"
  )
 port map (
   I0 => g0_b20_n_0,
   I1 => T1_27_i_25_n_0,
   I2 => h_20,
   O => T1_27_i_17_n_0
);
T1_27_i_18 : LUT3
  generic map(
   INIT => X"e8"
  )
 port map (
   I0 => g0_b19_n_0,
   I1 => T1_27_i_26_n_0,
   I2 => h_19,
   O => T1_27_i_18_n_0
);
T1_27_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => g0_b23_n_0,
   I1 => T1_31_i_41_n_0,
   I2 => h_23,
   I3 => T1_27_i_15_n_0,
   O => T1_27_i_19_n_0
);
T1_27_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => ROTR11_out_11,
   I1 => ROTR11_out_6,
   I2 => ROTR11_out_24,
   I3 => T1_reg_31_i_13_n_5,
   I4 => T1_27_i_10_n_0,
   O => T1_27_i_2_n_0
);
T1_27_i_20 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => g0_b22_n_0,
   I1 => T1_27_i_23_n_0,
   I2 => h_22,
   I3 => T1_27_i_16_n_0,
   O => T1_27_i_20_n_0
);
T1_27_i_21 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => g0_b21_n_0,
   I1 => T1_27_i_24_n_0,
   I2 => h_21,
   I3 => T1_27_i_17_n_0,
   O => T1_27_i_21_n_0
);
T1_27_i_22 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => g0_b20_n_0,
   I1 => T1_27_i_25_n_0,
   I2 => h_20,
   I3 => T1_27_i_18_n_0,
   O => T1_27_i_22_n_0
);
T1_27_i_23 : LUT6
  generic map(
   INIT => X"505f505fc0c0cfcf"
  )
 port map (
   I0 => T1_27_i_27_n_0,
   I1 => T1_reg_27_i_28_n_0,
   I2 => HASH_02_COUNTER_5,
   I3 => T1_27_i_29_n_0,
   I4 => T1_27_i_30_n_0,
   I5 => HASH_02_COUNTER_4,
   O => T1_27_i_23_n_0
);
T1_27_i_24 : LUT6
  generic map(
   INIT => X"303f303f50505f5f"
  )
 port map (
   I0 => T1_27_i_31_n_0,
   I1 => T1_27_i_32_n_0,
   I2 => HASH_02_COUNTER_5,
   I3 => T1_27_i_33_n_0,
   I4 => T1_27_i_34_n_0,
   I5 => HASH_02_COUNTER_4,
   O => T1_27_i_24_n_0
);
T1_27_i_25 : LUT6
  generic map(
   INIT => X"505f505f30303f3f"
  )
 port map (
   I0 => T1_27_i_35_n_0,
   I1 => T1_27_i_36_n_0,
   I2 => HASH_02_COUNTER_5,
   I3 => T1_27_i_37_n_0,
   I4 => T1_27_i_38_n_0,
   I5 => HASH_02_COUNTER_4,
   O => T1_27_i_25_n_0
);
T1_27_i_26 : LUT6
  generic map(
   INIT => X"505f505f30303f3f"
  )
 port map (
   I0 => T1_27_i_39_n_0,
   I1 => T1_27_i_40_n_0,
   I2 => HASH_02_COUNTER_5,
   I3 => T1_27_i_41_n_0,
   I4 => T1_27_i_42_n_0,
   I5 => HASH_02_COUNTER_4,
   O => T1_27_i_26_n_0
);
T1_27_i_27 : LUT6
  generic map(
   INIT => X"505f3030505f3f3f"
  )
 port map (
   I0 => T1_27_i_43_n_0,
   I1 => T1_27_i_44_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_27_i_45_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_27_i_46_n_0,
   O => T1_27_i_27_n_0
);
T1_27_i_29 : LUT6
  generic map(
   INIT => X"3030505f3f3f505f"
  )
 port map (
   I0 => T1_27_i_49_n_0,
   I1 => T1_27_i_50_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_27_i_51_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_27_i_52_n_0,
   O => T1_27_i_29_n_0
);
T1_27_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => ROTR11_out_12,
   I1 => ROTR11_out_7,
   I2 => ROTR11_out_25,
   I3 => T1_reg_31_i_13_n_6,
   I4 => T1_27_i_11_n_0,
   O => T1_27_i_3_n_0
);
T1_27_i_30 : LUT6
  generic map(
   INIT => X"5050303f5f5f303f"
  )
 port map (
   I0 => T1_27_i_53_n_0,
   I1 => T1_27_i_54_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_27_i_55_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_27_i_56_n_0,
   O => T1_27_i_30_n_0
);
T1_27_i_31 : LUT6
  generic map(
   INIT => X"505f3030505f3f3f"
  )
 port map (
   I0 => T1_27_i_57_n_0,
   I1 => T1_27_i_58_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_27_i_59_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_27_i_60_n_0,
   O => T1_27_i_31_n_0
);
T1_27_i_32 : LUT6
  generic map(
   INIT => X"3030505f3f3f505f"
  )
 port map (
   I0 => T1_27_i_61_n_0,
   I1 => T1_27_i_62_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_27_i_63_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_27_i_64_n_0,
   O => T1_27_i_32_n_0
);
T1_27_i_33 : LUT6
  generic map(
   INIT => X"3030505f3f3f505f"
  )
 port map (
   I0 => T1_27_i_65_n_0,
   I1 => T1_27_i_66_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_27_i_67_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_27_i_68_n_0,
   O => T1_27_i_33_n_0
);
T1_27_i_34 : LUT6
  generic map(
   INIT => X"505f3030505f3f3f"
  )
 port map (
   I0 => T1_27_i_69_n_0,
   I1 => T1_27_i_70_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_27_i_71_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_27_i_72_n_0,
   O => T1_27_i_34_n_0
);
T1_27_i_35 : LUT6
  generic map(
   INIT => X"3030505f3f3f505f"
  )
 port map (
   I0 => T1_27_i_73_n_0,
   I1 => T1_27_i_74_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_27_i_75_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_27_i_76_n_0,
   O => T1_27_i_35_n_0
);
T1_27_i_36 : LUT6
  generic map(
   INIT => X"505f3030505f3f3f"
  )
 port map (
   I0 => T1_27_i_77_n_0,
   I1 => T1_27_i_78_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_27_i_79_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_27_i_80_n_0,
   O => T1_27_i_36_n_0
);
T1_27_i_37 : LUT6
  generic map(
   INIT => X"505f3030505f3f3f"
  )
 port map (
   I0 => T1_27_i_81_n_0,
   I1 => T1_27_i_82_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_27_i_83_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_27_i_84_n_0,
   O => T1_27_i_37_n_0
);
T1_27_i_38 : LUT6
  generic map(
   INIT => X"5050303f5f5f303f"
  )
 port map (
   I0 => T1_27_i_85_n_0,
   I1 => T1_27_i_86_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_27_i_87_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_27_i_88_n_0,
   O => T1_27_i_38_n_0
);
T1_27_i_39 : LUT6
  generic map(
   INIT => X"5050303f5f5f303f"
  )
 port map (
   I0 => T1_27_i_89_n_0,
   I1 => T1_27_i_90_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_27_i_91_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_27_i_92_n_0,
   O => T1_27_i_39_n_0
);
T1_27_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => ROTR11_out_13,
   I1 => ROTR11_out_8,
   I2 => ROTR11_out_26,
   I3 => T1_reg_31_i_13_n_7,
   I4 => T1_27_i_12_n_0,
   O => T1_27_i_4_n_0
);
T1_27_i_40 : LUT6
  generic map(
   INIT => X"3030505f3f3f505f"
  )
 port map (
   I0 => T1_27_i_93_n_0,
   I1 => T1_27_i_94_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_27_i_95_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_27_i_96_n_0,
   O => T1_27_i_40_n_0
);
T1_27_i_41 : LUT6
  generic map(
   INIT => X"303f5050303f5f5f"
  )
 port map (
   I0 => T1_27_i_97_n_0,
   I1 => T1_27_i_98_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_27_i_99_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_27_i_100_n_0,
   O => T1_27_i_41_n_0
);
T1_27_i_42 : LUT6
  generic map(
   INIT => X"505f3030505f3f3f"
  )
 port map (
   I0 => T1_27_i_101_n_0,
   I1 => T1_27_i_102_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_27_i_103_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_27_i_104_n_0,
   O => T1_27_i_42_n_0
);
T1_27_i_43 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_63_22,
   I1 => W_reg_62_22,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_61_22,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_60_22,
   O => T1_27_i_43_n_0
);
T1_27_i_44 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_59_22,
   I1 => W_reg_58_22,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_57_22,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_56_22,
   O => T1_27_i_44_n_0
);
T1_27_i_45 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_55_22,
   I1 => W_reg_54_22,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_53_22,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_52_22,
   O => T1_27_i_45_n_0
);
T1_27_i_46 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_51_22,
   I1 => W_reg_50_22,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_49_22,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_48_22,
   O => T1_27_i_46_n_0
);
T1_27_i_49 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_27_22,
   I1 => W_reg_26_22,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_25_22,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_24_22,
   O => T1_27_i_49_n_0
);
T1_27_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => ROTR11_out_14,
   I1 => ROTR11_out_9,
   I2 => ROTR11_out_27,
   I3 => T1_reg_27_i_13_n_4,
   I4 => T1_27_i_14_n_0,
   O => T1_27_i_5_n_0
);
T1_27_i_50 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_31_22,
   I1 => W_reg_30_22,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_29_22,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_28_22,
   O => T1_27_i_50_n_0
);
T1_27_i_51 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_19_22,
   I1 => W_reg_18_22,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_17_22,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_16_22,
   O => T1_27_i_51_n_0
);
T1_27_i_52 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_23_22,
   I1 => W_reg_22_22,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_21_22,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_20_22,
   O => T1_27_i_52_n_0
);
T1_27_i_53 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_15_22,
   I1 => W_reg_14_22,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_13_22,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_12_22,
   O => T1_27_i_53_n_0
);
T1_27_i_54 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_11_22,
   I1 => W_reg_10_22,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_9_22,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_8_22,
   O => T1_27_i_54_n_0
);
T1_27_i_55 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_3_22,
   I1 => W_reg_2_22,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_1_22,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_0_22,
   O => T1_27_i_55_n_0
);
T1_27_i_56 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_7_22,
   I1 => W_reg_6_22,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_5_22,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_4_22,
   O => T1_27_i_56_n_0
);
T1_27_i_57 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_47_21,
   I1 => W_reg_46_21,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_45_21,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_44_21,
   O => T1_27_i_57_n_0
);
T1_27_i_58 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_43_21,
   I1 => W_reg_42_21,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_41_21,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_40_21,
   O => T1_27_i_58_n_0
);
T1_27_i_59 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_39_21,
   I1 => W_reg_38_21,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_37_21,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_36_21,
   O => T1_27_i_59_n_0
);
T1_27_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => T1_27_i_2_n_0,
   I1 => T1_reg_31_i_13_n_4,
   I2 => T1_31_i_14_n_0,
   I3 => ROTR11_out_5,
   I4 => ROTR11_out_23,
   I5 => ROTR11_out_10,
   O => T1_27_i_6_n_0
);
T1_27_i_60 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_35_21,
   I1 => W_reg_34_21,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_33_21,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_32_21,
   O => T1_27_i_60_n_0
);
T1_27_i_61 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_59_21,
   I1 => W_reg_58_21,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_57_21,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_56_21,
   O => T1_27_i_61_n_0
);
T1_27_i_62 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_63_21,
   I1 => W_reg_62_21,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_61_21,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_60_21,
   O => T1_27_i_62_n_0
);
T1_27_i_63 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_51_21,
   I1 => W_reg_50_21,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_49_21,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_48_21,
   O => T1_27_i_63_n_0
);
T1_27_i_64 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_55_21,
   I1 => W_reg_54_21,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_53_21,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_52_21,
   O => T1_27_i_64_n_0
);
T1_27_i_65 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_27_21,
   I1 => W_reg_26_21,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_25_21,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_24_21,
   O => T1_27_i_65_n_0
);
T1_27_i_66 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_31_21,
   I1 => W_reg_30_21,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_29_21,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_28_21,
   O => T1_27_i_66_n_0
);
T1_27_i_67 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_19_21,
   I1 => W_reg_18_21,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_17_21,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_16_21,
   O => T1_27_i_67_n_0
);
T1_27_i_68 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_23_21,
   I1 => W_reg_22_21,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_21_21,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_20_21,
   O => T1_27_i_68_n_0
);
T1_27_i_69 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_15_21,
   I1 => W_reg_14_21,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_13_21,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_12_21,
   O => T1_27_i_69_n_0
);
T1_27_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => T1_27_i_3_n_0,
   I1 => ROTR11_out_11,
   I2 => ROTR11_out_6,
   I3 => ROTR11_out_24,
   I4 => T1_reg_31_i_13_n_5,
   I5 => T1_27_i_10_n_0,
   O => T1_27_i_7_n_0
);
T1_27_i_70 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_11_21,
   I1 => W_reg_10_21,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_9_21,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_8_21,
   O => T1_27_i_70_n_0
);
T1_27_i_71 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_7_21,
   I1 => W_reg_6_21,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_5_21,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_4_21,
   O => T1_27_i_71_n_0
);
T1_27_i_72 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_3_21,
   I1 => W_reg_2_21,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_1_21,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_0_21,
   O => T1_27_i_72_n_0
);
T1_27_i_73 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_59_20,
   I1 => W_reg_58_20,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_57_20,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_56_20,
   O => T1_27_i_73_n_0
);
T1_27_i_74 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_63_20,
   I1 => W_reg_62_20,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_61_20,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_60_20,
   O => T1_27_i_74_n_0
);
T1_27_i_75 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_51_20,
   I1 => W_reg_50_20,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_49_20,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_48_20,
   O => T1_27_i_75_n_0
);
T1_27_i_76 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_55_20,
   I1 => W_reg_54_20,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_53_20,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_52_20,
   O => T1_27_i_76_n_0
);
T1_27_i_77 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_47_20,
   I1 => W_reg_46_20,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_45_20,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_44_20,
   O => T1_27_i_77_n_0
);
T1_27_i_78 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_43_20,
   I1 => W_reg_42_20,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_41_20,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_40_20,
   O => T1_27_i_78_n_0
);
T1_27_i_79 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_39_20,
   I1 => W_reg_38_20,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_37_20,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_36_20,
   O => T1_27_i_79_n_0
);
T1_27_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => T1_27_i_4_n_0,
   I1 => ROTR11_out_12,
   I2 => ROTR11_out_7,
   I3 => ROTR11_out_25,
   I4 => T1_reg_31_i_13_n_6,
   I5 => T1_27_i_11_n_0,
   O => T1_27_i_8_n_0
);
T1_27_i_80 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_35_20,
   I1 => W_reg_34_20,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_33_20,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_32_20,
   O => T1_27_i_80_n_0
);
T1_27_i_81 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_31_20,
   I1 => W_reg_30_20,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_29_20,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_28_20,
   O => T1_27_i_81_n_0
);
T1_27_i_82 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_27_20,
   I1 => W_reg_26_20,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_25_20,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_24_20,
   O => T1_27_i_82_n_0
);
T1_27_i_83 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_23_20,
   I1 => W_reg_22_20,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_21_20,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_20_20,
   O => T1_27_i_83_n_0
);
T1_27_i_84 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_19_20,
   I1 => W_reg_18_20,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_17_20,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_16_20,
   O => T1_27_i_84_n_0
);
T1_27_i_85 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_15_20,
   I1 => W_reg_14_20,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_13_20,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_12_20,
   O => T1_27_i_85_n_0
);
T1_27_i_86 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_11_20,
   I1 => W_reg_10_20,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_9_20,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_8_20,
   O => T1_27_i_86_n_0
);
T1_27_i_87 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_3_20,
   I1 => W_reg_2_20,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_1_20,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_0_20,
   O => T1_27_i_87_n_0
);
T1_27_i_88 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_7_20,
   I1 => W_reg_6_20,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_5_20,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_4_20,
   O => T1_27_i_88_n_0
);
T1_27_i_89 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_63_19,
   I1 => W_reg_62_19,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_61_19,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_60_19,
   O => T1_27_i_89_n_0
);
T1_27_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => T1_27_i_5_n_0,
   I1 => ROTR11_out_13,
   I2 => ROTR11_out_8,
   I3 => ROTR11_out_26,
   I4 => T1_reg_31_i_13_n_7,
   I5 => T1_27_i_12_n_0,
   O => T1_27_i_9_n_0
);
T1_27_i_90 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_59_19,
   I1 => W_reg_58_19,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_57_19,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_56_19,
   O => T1_27_i_90_n_0
);
T1_27_i_91 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_51_19,
   I1 => W_reg_50_19,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_49_19,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_48_19,
   O => T1_27_i_91_n_0
);
T1_27_i_92 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_55_19,
   I1 => W_reg_54_19,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_53_19,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_52_19,
   O => T1_27_i_92_n_0
);
T1_27_i_93 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_43_19,
   I1 => W_reg_42_19,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_41_19,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_40_19,
   O => T1_27_i_93_n_0
);
T1_27_i_94 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_47_19,
   I1 => W_reg_46_19,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_45_19,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_44_19,
   O => T1_27_i_94_n_0
);
T1_27_i_95 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_35_19,
   I1 => W_reg_34_19,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_33_19,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_32_19,
   O => T1_27_i_95_n_0
);
T1_27_i_96 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_39_19,
   I1 => W_reg_38_19,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_37_19,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_36_19,
   O => T1_27_i_96_n_0
);
T1_27_i_97 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_27_19,
   I1 => W_reg_26_19,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_25_19,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_24_19,
   O => T1_27_i_97_n_0
);
T1_27_i_98 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_31_19,
   I1 => W_reg_30_19,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_29_19,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_28_19,
   O => T1_27_i_98_n_0
);
T1_27_i_99 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_23_19,
   I1 => W_reg_22_19,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_21_19,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_20_19,
   O => T1_27_i_99_n_0
);
T1_31_i_1 : LUT5
  generic map(
   INIT => X"0000a8aa"
  )
 port map (
   I0 => FSM_onehot_CURRENT_STATE_reg_n_0_8,
   I1 => FSM_onehot_CURRENT_STATE_11_i_2_n_0,
   I2 => FSM_onehot_CURRENT_STATE_11_i_3_n_0,
   I3 => FSM_onehot_CURRENT_STATE_11_i_4_n_0,
   I4 => rst_IBUF,
   O => T1_31_i_1_n_0
);
T1_31_i_100 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_23_28,
   I1 => W_reg_22_28,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_21_28,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_20_28,
   O => T1_31_i_100_n_0
);
T1_31_i_101 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_19_28,
   I1 => W_reg_18_28,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_17_28,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_16_28,
   O => T1_31_i_101_n_0
);
T1_31_i_102 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_15_28,
   I1 => W_reg_14_28,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_13_28,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_12_28,
   O => T1_31_i_102_n_0
);
T1_31_i_103 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_11_28,
   I1 => W_reg_10_28,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_9_28,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_8_28,
   O => T1_31_i_103_n_0
);
T1_31_i_104 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_3_28,
   I1 => W_reg_2_28,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_1_28,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_0_28,
   O => T1_31_i_104_n_0
);
T1_31_i_105 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_7_28,
   I1 => W_reg_6_28,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_5_28,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_4_28,
   O => T1_31_i_105_n_0
);
T1_31_i_106 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_59_27,
   I1 => W_reg_58_27,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_57_27,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_56_27,
   O => T1_31_i_106_n_0
);
T1_31_i_107 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_63_27,
   I1 => W_reg_62_27,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_61_27,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_60_27,
   O => T1_31_i_107_n_0
);
T1_31_i_108 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_55_27,
   I1 => W_reg_54_27,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_53_27,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_52_27,
   O => T1_31_i_108_n_0
);
T1_31_i_109 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_51_27,
   I1 => W_reg_50_27,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_49_27,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_48_27,
   O => T1_31_i_109_n_0
);
T1_31_i_11 : LUT3
  generic map(
   INIT => X"b8"
  )
 port map (
   I0 => f_reg_n_0_29,
   I1 => ROTR11_out_14,
   I2 => g_reg_n_0_29,
   O => T1_31_i_11_n_0
);
T1_31_i_112 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_27_27,
   I1 => W_reg_26_27,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_25_27,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_24_27,
   O => T1_31_i_112_n_0
);
T1_31_i_113 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_31_27,
   I1 => W_reg_30_27,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_29_27,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_28_27,
   O => T1_31_i_113_n_0
);
T1_31_i_114 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_23_27,
   I1 => W_reg_22_27,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_21_27,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_20_27,
   O => T1_31_i_114_n_0
);
T1_31_i_115 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_19_27,
   I1 => W_reg_18_27,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_17_27,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_16_27,
   O => T1_31_i_115_n_0
);
T1_31_i_116 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_11_27,
   I1 => W_reg_10_27,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_9_27,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_8_27,
   O => T1_31_i_116_n_0
);
T1_31_i_117 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_15_27,
   I1 => W_reg_14_27,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_13_27,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_12_27,
   O => T1_31_i_117_n_0
);
T1_31_i_118 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_7_27,
   I1 => W_reg_6_27,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_5_27,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_4_27,
   O => T1_31_i_118_n_0
);
T1_31_i_119 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_3_27,
   I1 => W_reg_2_27,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_1_27,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_0_27,
   O => T1_31_i_119_n_0
);
T1_31_i_12 : LUT3
  generic map(
   INIT => X"b8"
  )
 port map (
   I0 => f_reg_n_0_28,
   I1 => ROTR11_out_15,
   I2 => g_reg_n_0_28,
   O => T1_31_i_12_n_0
);
T1_31_i_128 : LUT6
  generic map(
   INIT => X"05f5030305f5f3f3"
  )
 port map (
   I0 => T1_31_i_216_n_0,
   I1 => T1_31_i_217_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_31_i_218_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_31_i_219_n_0,
   O => T1_31_i_128_n_0
);
T1_31_i_129 : LUT6
  generic map(
   INIT => X"3030505f3f3f505f"
  )
 port map (
   I0 => T1_31_i_220_n_0,
   I1 => T1_31_i_221_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_31_i_222_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_31_i_223_n_0,
   O => T1_31_i_129_n_0
);
T1_31_i_130 : LUT6
  generic map(
   INIT => X"5050303f5f5f303f"
  )
 port map (
   I0 => T1_31_i_224_n_0,
   I1 => T1_31_i_225_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_31_i_226_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_31_i_227_n_0,
   O => T1_31_i_130_n_0
);
T1_31_i_131 : LUT6
  generic map(
   INIT => X"5050303f5f5f303f"
  )
 port map (
   I0 => T1_31_i_228_n_0,
   I1 => T1_31_i_229_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_31_i_230_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_31_i_231_n_0,
   O => T1_31_i_131_n_0
);
T1_31_i_132 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_63_26,
   I1 => W_reg_62_26,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_61_26,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_60_26,
   O => T1_31_i_132_n_0
);
T1_31_i_133 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_59_26,
   I1 => W_reg_58_26,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_57_26,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_56_26,
   O => T1_31_i_133_n_0
);
T1_31_i_134 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_55_26,
   I1 => W_reg_54_26,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_53_26,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_52_26,
   O => T1_31_i_134_n_0
);
T1_31_i_135 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_51_26,
   I1 => W_reg_50_26,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_49_26,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_48_26,
   O => T1_31_i_135_n_0
);
T1_31_i_138 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_27_26,
   I1 => W_reg_26_26,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_25_26,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_24_26,
   O => T1_31_i_138_n_0
);
T1_31_i_139 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_31_26,
   I1 => W_reg_30_26,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_29_26,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_28_26,
   O => T1_31_i_139_n_0
);
T1_31_i_14 : LUT3
  generic map(
   INIT => X"b8"
  )
 port map (
   I0 => f_reg_n_0_27,
   I1 => ROTR11_out_16,
   I2 => g_reg_n_0_27,
   O => T1_31_i_14_n_0
);
T1_31_i_140 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_19_26,
   I1 => W_reg_18_26,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_17_26,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_16_26,
   O => T1_31_i_140_n_0
);
T1_31_i_141 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_23_26,
   I1 => W_reg_22_26,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_21_26,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_20_26,
   O => T1_31_i_141_n_0
);
T1_31_i_142 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_15_26,
   I1 => W_reg_14_26,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_13_26,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_12_26,
   O => T1_31_i_142_n_0
);
T1_31_i_143 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_11_26,
   I1 => W_reg_10_26,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_9_26,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_8_26,
   O => T1_31_i_143_n_0
);
T1_31_i_144 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_7_26,
   I1 => W_reg_6_26,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_5_26,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_4_26,
   O => T1_31_i_144_n_0
);
T1_31_i_145 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_3_26,
   I1 => W_reg_2_26,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_1_26,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_0_26,
   O => T1_31_i_145_n_0
);
T1_31_i_146 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_59_25,
   I1 => W_reg_58_25,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_57_25,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_56_25,
   O => T1_31_i_146_n_0
);
T1_31_i_147 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_63_25,
   I1 => W_reg_62_25,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_61_25,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_60_25,
   O => T1_31_i_147_n_0
);
T1_31_i_148 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_55_25,
   I1 => W_reg_54_25,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_53_25,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_52_25,
   O => T1_31_i_148_n_0
);
T1_31_i_149 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_51_25,
   I1 => W_reg_50_25,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_49_25,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_48_25,
   O => T1_31_i_149_n_0
);
T1_31_i_15 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => ROTR11_out_19,
   I1 => ROTR11_out_6,
   I2 => ROTR11_out_1,
   I3 => T1_reg_31_i_10_n_4,
   O => T1_31_i_15_n_0
);
T1_31_i_152 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_27_25,
   I1 => W_reg_26_25,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_25_25,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_24_25,
   O => T1_31_i_152_n_0
);
T1_31_i_153 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_31_25,
   I1 => W_reg_30_25,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_29_25,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_28_25,
   O => T1_31_i_153_n_0
);
T1_31_i_154 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_19_25,
   I1 => W_reg_18_25,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_17_25,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_16_25,
   O => T1_31_i_154_n_0
);
T1_31_i_155 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_23_25,
   I1 => W_reg_22_25,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_21_25,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_20_25,
   O => T1_31_i_155_n_0
);
T1_31_i_156 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_15_25,
   I1 => W_reg_14_25,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_13_25,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_12_25,
   O => T1_31_i_156_n_0
);
T1_31_i_157 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_11_25,
   I1 => W_reg_10_25,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_9_25,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_8_25,
   O => T1_31_i_157_n_0
);
T1_31_i_158 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_3_25,
   I1 => W_reg_2_25,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_1_25,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_0_25,
   O => T1_31_i_158_n_0
);
T1_31_i_159 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_7_25,
   I1 => W_reg_6_25,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_5_25,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_4_25,
   O => T1_31_i_159_n_0
);
T1_31_i_16 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => ROTR11_out_2,
   I1 => ROTR11_out_20,
   I2 => ROTR11_out_7,
   I3 => T1_reg_31_i_10_n_5,
   I4 => T1_31_i_17_n_0,
   O => T1_31_i_16_n_0
);
T1_31_i_160 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_63_24,
   I1 => W_reg_62_24,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_61_24,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_60_24,
   O => T1_31_i_160_n_0
);
T1_31_i_161 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_59_24,
   I1 => W_reg_58_24,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_57_24,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_56_24,
   O => T1_31_i_161_n_0
);
T1_31_i_162 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_55_24,
   I1 => W_reg_54_24,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_53_24,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_52_24,
   O => T1_31_i_162_n_0
);
T1_31_i_163 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_51_24,
   I1 => W_reg_50_24,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_49_24,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_48_24,
   O => T1_31_i_163_n_0
);
T1_31_i_164 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_47_24,
   I1 => W_reg_46_24,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_45_24,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_44_24,
   O => T1_31_i_164_n_0
);
T1_31_i_165 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_43_24,
   I1 => W_reg_42_24,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_41_24,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_40_24,
   O => T1_31_i_165_n_0
);
T1_31_i_166 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_35_24,
   I1 => W_reg_34_24,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_33_24,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_32_24,
   O => T1_31_i_166_n_0
);
T1_31_i_167 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_39_24,
   I1 => W_reg_38_24,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_37_24,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_36_24,
   O => T1_31_i_167_n_0
);
T1_31_i_168 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_31_24,
   I1 => W_reg_30_24,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_29_24,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_28_24,
   O => T1_31_i_168_n_0
);
T1_31_i_169 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_27_24,
   I1 => W_reg_26_24,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_25_24,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_24_24,
   O => T1_31_i_169_n_0
);
T1_31_i_17 : LUT3
  generic map(
   INIT => X"b8"
  )
 port map (
   I0 => f_reg_n_0_30,
   I1 => ROTR11_out_13,
   I2 => g_reg_n_0_30,
   O => T1_31_i_17_n_0
);
T1_31_i_170 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_19_24,
   I1 => W_reg_18_24,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_17_24,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_16_24,
   O => T1_31_i_170_n_0
);
T1_31_i_171 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_23_24,
   I1 => W_reg_22_24,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_21_24,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_20_24,
   O => T1_31_i_171_n_0
);
T1_31_i_172 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_15_24,
   I1 => W_reg_14_24,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_13_24,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_12_24,
   O => T1_31_i_172_n_0
);
T1_31_i_173 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_11_24,
   I1 => W_reg_10_24,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_9_24,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_8_24,
   O => T1_31_i_173_n_0
);
T1_31_i_174 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_3_24,
   I1 => W_reg_2_24,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_1_24,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_0_24,
   O => T1_31_i_174_n_0
);
T1_31_i_175 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_7_24,
   I1 => W_reg_6_24,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_5_24,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_4_24,
   O => T1_31_i_175_n_0
);
T1_31_i_176 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_63_23,
   I1 => W_reg_62_23,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_61_23,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_60_23,
   O => T1_31_i_176_n_0
);
T1_31_i_177 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_59_23,
   I1 => W_reg_58_23,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_57_23,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_56_23,
   O => T1_31_i_177_n_0
);
T1_31_i_178 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_55_23,
   I1 => W_reg_54_23,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_53_23,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_52_23,
   O => T1_31_i_178_n_0
);
T1_31_i_179 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_51_23,
   I1 => W_reg_50_23,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_49_23,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_48_23,
   O => T1_31_i_179_n_0
);
T1_31_i_18 : LUT3
  generic map(
   INIT => X"e8"
  )
 port map (
   I0 => g0_b29_n_0,
   I1 => T1_31_i_33_n_0,
   I2 => h_29,
   O => T1_31_i_18_n_0
);
T1_31_i_180 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_47_23,
   I1 => W_reg_46_23,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_45_23,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_44_23,
   O => T1_31_i_180_n_0
);
T1_31_i_181 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_43_23,
   I1 => W_reg_42_23,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_41_23,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_40_23,
   O => T1_31_i_181_n_0
);
T1_31_i_182 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_39_23,
   I1 => W_reg_38_23,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_37_23,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_36_23,
   O => T1_31_i_182_n_0
);
T1_31_i_183 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_35_23,
   I1 => W_reg_34_23,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_33_23,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_32_23,
   O => T1_31_i_183_n_0
);
T1_31_i_184 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_27_23,
   I1 => W_reg_26_23,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_25_23,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_24_23,
   O => T1_31_i_184_n_0
);
T1_31_i_185 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_31_23,
   I1 => W_reg_30_23,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_29_23,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_28_23,
   O => T1_31_i_185_n_0
);
T1_31_i_186 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_23_23,
   I1 => W_reg_22_23,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_21_23,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_20_23,
   O => T1_31_i_186_n_0
);
T1_31_i_187 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_19_23,
   I1 => W_reg_18_23,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_17_23,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_16_23,
   O => T1_31_i_187_n_0
);
T1_31_i_188 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_15_23,
   I1 => W_reg_14_23,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_13_23,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_12_23,
   O => T1_31_i_188_n_0
);
T1_31_i_189 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_11_23,
   I1 => W_reg_10_23,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_9_23,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_8_23,
   O => T1_31_i_189_n_0
);
T1_31_i_19 : LUT3
  generic map(
   INIT => X"e8"
  )
 port map (
   I0 => g0_b28_n_0,
   I1 => T1_31_i_34_n_0,
   I2 => h_28,
   O => T1_31_i_19_n_0
);
T1_31_i_190 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_3_23,
   I1 => W_reg_2_23,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_1_23,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_0_23,
   O => T1_31_i_190_n_0
);
T1_31_i_191 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_7_23,
   I1 => W_reg_6_23,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_5_23,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_4_23,
   O => T1_31_i_191_n_0
);
T1_31_i_192 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_35_28,
   I1 => W_reg_34_28,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_33_28,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_32_28,
   O => T1_31_i_192_n_0
);
T1_31_i_193 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_39_28,
   I1 => W_reg_38_28,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_37_28,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_36_28,
   O => T1_31_i_193_n_0
);
T1_31_i_194 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_43_28,
   I1 => W_reg_42_28,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_41_28,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_40_28,
   O => T1_31_i_194_n_0
);
T1_31_i_195 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_47_28,
   I1 => W_reg_46_28,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_45_28,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_44_28,
   O => T1_31_i_195_n_0
);
T1_31_i_196 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_35_27,
   I1 => W_reg_34_27,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_33_27,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_32_27,
   O => T1_31_i_196_n_0
);
T1_31_i_197 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_39_27,
   I1 => W_reg_38_27,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_37_27,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_36_27,
   O => T1_31_i_197_n_0
);
T1_31_i_198 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_43_27,
   I1 => W_reg_42_27,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_41_27,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_40_27,
   O => T1_31_i_198_n_0
);
T1_31_i_199 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_47_27,
   I1 => W_reg_46_27,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_45_27,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_44_27,
   O => T1_31_i_199_n_0
);
T1_31_i_20 : LUT3
  generic map(
   INIT => X"e8"
  )
 port map (
   I0 => g0_b27_n_0,
   I1 => T1_31_i_35_n_0,
   I2 => h_27,
   O => T1_31_i_20_n_0
);
T1_31_i_200 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_51_30,
   I1 => W_reg_50_30,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_49_30,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_48_30,
   O => T1_31_i_200_n_0
);
T1_31_i_201 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_55_30,
   I1 => W_reg_54_30,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_53_30,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_52_30,
   O => T1_31_i_201_n_0
);
T1_31_i_202 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_59_30,
   I1 => W_reg_58_30,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_57_30,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_56_30,
   O => T1_31_i_202_n_0
);
T1_31_i_203 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_63_30,
   I1 => W_reg_62_30,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_61_30,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_60_30,
   O => T1_31_i_203_n_0
);
T1_31_i_204 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_35_30,
   I1 => W_reg_34_30,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_33_30,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_32_30,
   O => T1_31_i_204_n_0
);
T1_31_i_205 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_39_30,
   I1 => W_reg_38_30,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_37_30,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_36_30,
   O => T1_31_i_205_n_0
);
T1_31_i_206 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_43_30,
   I1 => W_reg_42_30,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_41_30,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_40_30,
   O => T1_31_i_206_n_0
);
T1_31_i_207 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_47_30,
   I1 => W_reg_46_30,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_45_30,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_44_30,
   O => T1_31_i_207_n_0
);
T1_31_i_208 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_19_30,
   I1 => W_reg_18_30,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_17_30,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_16_30,
   O => T1_31_i_208_n_0
);
T1_31_i_209 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_23_30,
   I1 => W_reg_22_30,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_21_30,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_20_30,
   O => T1_31_i_209_n_0
);
T1_31_i_21 : LUT6
  generic map(
   INIT => X"e81717e817e8e817"
  )
 port map (
   I0 => h_30,
   I1 => T1_31_i_36_n_0,
   I2 => g0_b30_n_0,
   I3 => g0_b31_n_0,
   I4 => h_31,
   I5 => T1_reg_31_i_37_n_0,
   O => T1_31_i_21_n_0
);
T1_31_i_210 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_27_30,
   I1 => W_reg_26_30,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_25_30,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_24_30,
   O => T1_31_i_210_n_0
);
T1_31_i_211 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_31_30,
   I1 => W_reg_30_30,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_29_30,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_28_30,
   O => T1_31_i_211_n_0
);
T1_31_i_212 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_3_30,
   I1 => W_reg_2_30,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_1_30,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_0_30,
   O => T1_31_i_212_n_0
);
T1_31_i_213 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_7_30,
   I1 => W_reg_6_30,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_5_30,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_4_30,
   O => T1_31_i_213_n_0
);
T1_31_i_214 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_11_30,
   I1 => W_reg_10_30,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_9_30,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_8_30,
   O => T1_31_i_214_n_0
);
T1_31_i_215 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_15_30,
   I1 => W_reg_14_30,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_13_30,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_12_30,
   O => T1_31_i_215_n_0
);
T1_31_i_216 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_7_31,
   I1 => W_reg_6_31,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_5_31,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_4_31,
   O => T1_31_i_216_n_0
);
T1_31_i_217 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_3_31,
   I1 => W_reg_2_31,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_1_31,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_0_31,
   O => T1_31_i_217_n_0
);
T1_31_i_218 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_15_31,
   I1 => W_reg_14_31,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_13_31,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_12_31,
   O => T1_31_i_218_n_0
);
T1_31_i_219 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_11_31,
   I1 => W_reg_10_31,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_9_31,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_8_31,
   O => T1_31_i_219_n_0
);
T1_31_i_22 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => T1_31_i_18_n_0,
   I1 => g0_b30_n_0,
   I2 => T1_31_i_36_n_0,
   I3 => h_30,
   O => T1_31_i_22_n_0
);
T1_31_i_220 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_27_31,
   I1 => W_reg_26_31,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_25_31,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_24_31,
   O => T1_31_i_220_n_0
);
T1_31_i_221 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_31_31,
   I1 => W_reg_30_31,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_29_31,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_28_31,
   O => T1_31_i_221_n_0
);
T1_31_i_222 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_19_31,
   I1 => W_reg_18_31,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_17_31,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_16_31,
   O => T1_31_i_222_n_0
);
T1_31_i_223 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_23_31,
   I1 => W_reg_22_31,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_21_31,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_20_31,
   O => T1_31_i_223_n_0
);
T1_31_i_224 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_47_31,
   I1 => W_reg_46_31,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_45_31,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_44_31,
   O => T1_31_i_224_n_0
);
T1_31_i_225 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_43_31,
   I1 => W_reg_42_31,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_41_31,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_40_31,
   O => T1_31_i_225_n_0
);
T1_31_i_226 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_35_31,
   I1 => W_reg_34_31,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_33_31,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_32_31,
   O => T1_31_i_226_n_0
);
T1_31_i_227 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_39_31,
   I1 => W_reg_38_31,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_37_31,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_36_31,
   O => T1_31_i_227_n_0
);
T1_31_i_228 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_63_31,
   I1 => W_reg_62_31,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_61_31,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_60_31,
   O => T1_31_i_228_n_0
);
T1_31_i_229 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_59_31,
   I1 => W_reg_58_31,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_57_31,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_56_31,
   O => T1_31_i_229_n_0
);
T1_31_i_23 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => g0_b29_n_0,
   I1 => T1_31_i_33_n_0,
   I2 => h_29,
   I3 => T1_31_i_19_n_0,
   O => T1_31_i_23_n_0
);
T1_31_i_230 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_51_31,
   I1 => W_reg_50_31,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_49_31,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_48_31,
   O => T1_31_i_230_n_0
);
T1_31_i_231 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_55_31,
   I1 => W_reg_54_31,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_53_31,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_52_31,
   O => T1_31_i_231_n_0
);
T1_31_i_232 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_35_26,
   I1 => W_reg_34_26,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_33_26,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_32_26,
   O => T1_31_i_232_n_0
);
T1_31_i_233 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_39_26,
   I1 => W_reg_38_26,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_37_26,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_36_26,
   O => T1_31_i_233_n_0
);
T1_31_i_234 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_43_26,
   I1 => W_reg_42_26,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_41_26,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_40_26,
   O => T1_31_i_234_n_0
);
T1_31_i_235 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_47_26,
   I1 => W_reg_46_26,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_45_26,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_44_26,
   O => T1_31_i_235_n_0
);
T1_31_i_236 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_35_25,
   I1 => W_reg_34_25,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_33_25,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_32_25,
   O => T1_31_i_236_n_0
);
T1_31_i_237 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_39_25,
   I1 => W_reg_38_25,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_37_25,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_36_25,
   O => T1_31_i_237_n_0
);
T1_31_i_238 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_43_25,
   I1 => W_reg_42_25,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_41_25,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_40_25,
   O => T1_31_i_238_n_0
);
T1_31_i_239 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_47_25,
   I1 => W_reg_46_25,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_45_25,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_44_25,
   O => T1_31_i_239_n_0
);
T1_31_i_24 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => g0_b28_n_0,
   I1 => T1_31_i_34_n_0,
   I2 => h_28,
   I3 => T1_31_i_20_n_0,
   O => T1_31_i_24_n_0
);
T1_31_i_25 : LUT3
  generic map(
   INIT => X"e8"
  )
 port map (
   I0 => g0_b26_n_0,
   I1 => T1_31_i_38_n_0,
   I2 => h_26,
   O => T1_31_i_25_n_0
);
T1_31_i_26 : LUT3
  generic map(
   INIT => X"e8"
  )
 port map (
   I0 => g0_b25_n_0,
   I1 => T1_31_i_39_n_0,
   I2 => h_25,
   O => T1_31_i_26_n_0
);
T1_31_i_27 : LUT3
  generic map(
   INIT => X"e8"
  )
 port map (
   I0 => g0_b24_n_0,
   I1 => T1_31_i_40_n_0,
   I2 => h_24,
   O => T1_31_i_27_n_0
);
T1_31_i_28 : LUT3
  generic map(
   INIT => X"e8"
  )
 port map (
   I0 => g0_b23_n_0,
   I1 => T1_31_i_41_n_0,
   I2 => h_23,
   O => T1_31_i_28_n_0
);
T1_31_i_29 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => g0_b27_n_0,
   I1 => T1_31_i_35_n_0,
   I2 => h_27,
   I3 => T1_31_i_25_n_0,
   O => T1_31_i_29_n_0
);
T1_31_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => ROTR11_out_3,
   I1 => ROTR11_out_21,
   I2 => ROTR11_out_8,
   I3 => T1_reg_31_i_10_n_6,
   I4 => T1_31_i_11_n_0,
   O => T1_31_i_3_n_0
);
T1_31_i_30 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => g0_b26_n_0,
   I1 => T1_31_i_38_n_0,
   I2 => h_26,
   I3 => T1_31_i_26_n_0,
   O => T1_31_i_30_n_0
);
T1_31_i_31 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => g0_b25_n_0,
   I1 => T1_31_i_39_n_0,
   I2 => h_25,
   I3 => T1_31_i_27_n_0,
   O => T1_31_i_31_n_0
);
T1_31_i_32 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => g0_b24_n_0,
   I1 => T1_31_i_40_n_0,
   I2 => h_24,
   I3 => T1_31_i_28_n_0,
   O => T1_31_i_32_n_0
);
T1_31_i_33 : LUT6
  generic map(
   INIT => X"505f505f30303f3f"
  )
 port map (
   I0 => T1_31_i_42_n_0,
   I1 => T1_31_i_43_n_0,
   I2 => HASH_02_COUNTER_5,
   I3 => T1_31_i_44_n_0,
   I4 => T1_31_i_45_n_0,
   I5 => HASH_02_COUNTER_4,
   O => T1_31_i_33_n_0
);
T1_31_i_34 : LUT6
  generic map(
   INIT => X"505f505fc0c0cfcf"
  )
 port map (
   I0 => T1_31_i_46_n_0,
   I1 => T1_reg_31_i_47_n_0,
   I2 => HASH_02_COUNTER_5,
   I3 => T1_31_i_48_n_0,
   I4 => T1_31_i_49_n_0,
   I5 => HASH_02_COUNTER_4,
   O => T1_31_i_34_n_0
);
T1_31_i_35 : LUT6
  generic map(
   INIT => X"505f505fc0c0cfcf"
  )
 port map (
   I0 => T1_31_i_50_n_0,
   I1 => T1_reg_31_i_51_n_0,
   I2 => HASH_02_COUNTER_5,
   I3 => T1_31_i_52_n_0,
   I4 => T1_31_i_53_n_0,
   I5 => HASH_02_COUNTER_4,
   O => T1_31_i_35_n_0
);
T1_31_i_36 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => T1_reg_31_i_54_n_0,
   I1 => T1_reg_31_i_55_n_0,
   I2 => HASH_02_COUNTER_5,
   I3 => T1_reg_31_i_56_n_0,
   I4 => HASH_02_COUNTER_4,
   I5 => T1_reg_31_i_57_n_0,
   O => T1_31_i_36_n_0
);
T1_31_i_38 : LUT6
  generic map(
   INIT => X"505f505fc0c0cfcf"
  )
 port map (
   I0 => T1_31_i_60_n_0,
   I1 => T1_reg_31_i_61_n_0,
   I2 => HASH_02_COUNTER_5,
   I3 => T1_31_i_62_n_0,
   I4 => T1_31_i_63_n_0,
   I5 => HASH_02_COUNTER_4,
   O => T1_31_i_38_n_0
);
T1_31_i_39 : LUT6
  generic map(
   INIT => X"505f505fc0c0cfcf"
  )
 port map (
   I0 => T1_31_i_64_n_0,
   I1 => T1_reg_31_i_65_n_0,
   I2 => HASH_02_COUNTER_5,
   I3 => T1_31_i_66_n_0,
   I4 => T1_31_i_67_n_0,
   I5 => HASH_02_COUNTER_4,
   O => T1_31_i_39_n_0
);
T1_31_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => ROTR11_out_4,
   I1 => ROTR11_out_22,
   I2 => ROTR11_out_9,
   I3 => T1_reg_31_i_10_n_7,
   I4 => T1_31_i_12_n_0,
   O => T1_31_i_4_n_0
);
T1_31_i_40 : LUT6
  generic map(
   INIT => X"505f505f30303f3f"
  )
 port map (
   I0 => T1_31_i_68_n_0,
   I1 => T1_31_i_69_n_0,
   I2 => HASH_02_COUNTER_5,
   I3 => T1_31_i_70_n_0,
   I4 => T1_31_i_71_n_0,
   I5 => HASH_02_COUNTER_4,
   O => T1_31_i_40_n_0
);
T1_31_i_41 : LUT6
  generic map(
   INIT => X"505f505f30303f3f"
  )
 port map (
   I0 => T1_31_i_72_n_0,
   I1 => T1_31_i_73_n_0,
   I2 => HASH_02_COUNTER_5,
   I3 => T1_31_i_74_n_0,
   I4 => T1_31_i_75_n_0,
   I5 => HASH_02_COUNTER_4,
   O => T1_31_i_41_n_0
);
T1_31_i_42 : LUT6
  generic map(
   INIT => X"5050303f5f5f303f"
  )
 port map (
   I0 => T1_31_i_76_n_0,
   I1 => T1_31_i_77_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_31_i_78_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_31_i_79_n_0,
   O => T1_31_i_42_n_0
);
T1_31_i_43 : LUT6
  generic map(
   INIT => X"3030505f3f3f505f"
  )
 port map (
   I0 => T1_31_i_80_n_0,
   I1 => T1_31_i_81_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_31_i_82_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_31_i_83_n_0,
   O => T1_31_i_43_n_0
);
T1_31_i_44 : LUT6
  generic map(
   INIT => X"505f3030505f3f3f"
  )
 port map (
   I0 => T1_31_i_84_n_0,
   I1 => T1_31_i_85_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_31_i_86_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_31_i_87_n_0,
   O => T1_31_i_44_n_0
);
T1_31_i_45 : LUT6
  generic map(
   INIT => X"505f3030505f3f3f"
  )
 port map (
   I0 => T1_31_i_88_n_0,
   I1 => T1_31_i_89_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_31_i_90_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_31_i_91_n_0,
   O => T1_31_i_45_n_0
);
T1_31_i_46 : LUT6
  generic map(
   INIT => X"3030505f3f3f505f"
  )
 port map (
   I0 => T1_31_i_92_n_0,
   I1 => T1_31_i_93_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_31_i_94_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_31_i_95_n_0,
   O => T1_31_i_46_n_0
);
T1_31_i_48 : LUT6
  generic map(
   INIT => X"303f5050303f5f5f"
  )
 port map (
   I0 => T1_31_i_98_n_0,
   I1 => T1_31_i_99_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_31_i_100_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_31_i_101_n_0,
   O => T1_31_i_48_n_0
);
T1_31_i_49 : LUT6
  generic map(
   INIT => X"5050303f5f5f303f"
  )
 port map (
   I0 => T1_31_i_102_n_0,
   I1 => T1_31_i_103_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_31_i_104_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_31_i_105_n_0,
   O => T1_31_i_49_n_0
);
T1_31_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => ROTR11_out_5,
   I1 => ROTR11_out_23,
   I2 => ROTR11_out_10,
   I3 => T1_reg_31_i_13_n_4,
   I4 => T1_31_i_14_n_0,
   O => T1_31_i_5_n_0
);
T1_31_i_50 : LUT6
  generic map(
   INIT => X"303f5050303f5f5f"
  )
 port map (
   I0 => T1_31_i_106_n_0,
   I1 => T1_31_i_107_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_31_i_108_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_31_i_109_n_0,
   O => T1_31_i_50_n_0
);
T1_31_i_52 : LUT6
  generic map(
   INIT => X"303f5050303f5f5f"
  )
 port map (
   I0 => T1_31_i_112_n_0,
   I1 => T1_31_i_113_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_31_i_114_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_31_i_115_n_0,
   O => T1_31_i_52_n_0
);
T1_31_i_53 : LUT6
  generic map(
   INIT => X"303f5050303f5f5f"
  )
 port map (
   I0 => T1_31_i_116_n_0,
   I1 => T1_31_i_117_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_31_i_118_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_31_i_119_n_0,
   O => T1_31_i_53_n_0
);
T1_31_i_6 : LUT5
  generic map(
   INIT => X"b84747b8"
  )
 port map (
   I0 => f_reg_n_0_31,
   I1 => ROTR11_out_12,
   I2 => g_reg_n_0_31,
   I3 => T1_31_i_15_n_0,
   I4 => T1_31_i_16_n_0,
   O => T1_31_i_6_n_0
);
T1_31_i_60 : LUT6
  generic map(
   INIT => X"505f3030505f3f3f"
  )
 port map (
   I0 => T1_31_i_132_n_0,
   I1 => T1_31_i_133_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_31_i_134_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_31_i_135_n_0,
   O => T1_31_i_60_n_0
);
T1_31_i_62 : LUT6
  generic map(
   INIT => X"3030505f3f3f505f"
  )
 port map (
   I0 => T1_31_i_138_n_0,
   I1 => T1_31_i_139_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_31_i_140_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_31_i_141_n_0,
   O => T1_31_i_62_n_0
);
T1_31_i_63 : LUT6
  generic map(
   INIT => X"505f3030505f3f3f"
  )
 port map (
   I0 => T1_31_i_142_n_0,
   I1 => T1_31_i_143_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_31_i_144_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_31_i_145_n_0,
   O => T1_31_i_63_n_0
);
T1_31_i_64 : LUT6
  generic map(
   INIT => X"303f5050303f5f5f"
  )
 port map (
   I0 => T1_31_i_146_n_0,
   I1 => T1_31_i_147_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_31_i_148_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_31_i_149_n_0,
   O => T1_31_i_64_n_0
);
T1_31_i_66 : LUT6
  generic map(
   INIT => X"3030505f3f3f505f"
  )
 port map (
   I0 => T1_31_i_152_n_0,
   I1 => T1_31_i_153_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_31_i_154_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_31_i_155_n_0,
   O => T1_31_i_66_n_0
);
T1_31_i_67 : LUT6
  generic map(
   INIT => X"5050303f5f5f303f"
  )
 port map (
   I0 => T1_31_i_156_n_0,
   I1 => T1_31_i_157_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_31_i_158_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_31_i_159_n_0,
   O => T1_31_i_67_n_0
);
T1_31_i_68 : LUT6
  generic map(
   INIT => X"505f3030505f3f3f"
  )
 port map (
   I0 => T1_31_i_160_n_0,
   I1 => T1_31_i_161_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_31_i_162_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_31_i_163_n_0,
   O => T1_31_i_68_n_0
);
T1_31_i_69 : LUT6
  generic map(
   INIT => X"5050303f5f5f303f"
  )
 port map (
   I0 => T1_31_i_164_n_0,
   I1 => T1_31_i_165_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_31_i_166_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_31_i_167_n_0,
   O => T1_31_i_69_n_0
);
T1_31_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => T1_31_i_3_n_0,
   I1 => ROTR11_out_2,
   I2 => ROTR11_out_20,
   I3 => ROTR11_out_7,
   I4 => T1_reg_31_i_10_n_5,
   I5 => T1_31_i_17_n_0,
   O => T1_31_i_7_n_0
);
T1_31_i_70 : LUT6
  generic map(
   INIT => X"5050303f5f5f303f"
  )
 port map (
   I0 => T1_31_i_168_n_0,
   I1 => T1_31_i_169_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_31_i_170_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_31_i_171_n_0,
   O => T1_31_i_70_n_0
);
T1_31_i_71 : LUT6
  generic map(
   INIT => X"5050303f5f5f303f"
  )
 port map (
   I0 => T1_31_i_172_n_0,
   I1 => T1_31_i_173_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_31_i_174_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_31_i_175_n_0,
   O => T1_31_i_71_n_0
);
T1_31_i_72 : LUT6
  generic map(
   INIT => X"505f3030505f3f3f"
  )
 port map (
   I0 => T1_31_i_176_n_0,
   I1 => T1_31_i_177_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_31_i_178_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_31_i_179_n_0,
   O => T1_31_i_72_n_0
);
T1_31_i_73 : LUT6
  generic map(
   INIT => X"505f3030505f3f3f"
  )
 port map (
   I0 => T1_31_i_180_n_0,
   I1 => T1_31_i_181_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_31_i_182_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_31_i_183_n_0,
   O => T1_31_i_73_n_0
);
T1_31_i_74 : LUT6
  generic map(
   INIT => X"303f5050303f5f5f"
  )
 port map (
   I0 => T1_31_i_184_n_0,
   I1 => T1_31_i_185_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_31_i_186_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_31_i_187_n_0,
   O => T1_31_i_74_n_0
);
T1_31_i_75 : LUT6
  generic map(
   INIT => X"5050303f5f5f303f"
  )
 port map (
   I0 => T1_31_i_188_n_0,
   I1 => T1_31_i_189_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_31_i_190_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_31_i_191_n_0,
   O => T1_31_i_75_n_0
);
T1_31_i_76 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_63_29,
   I1 => W_reg_62_29,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_61_29,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_60_29,
   O => T1_31_i_76_n_0
);
T1_31_i_77 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_59_29,
   I1 => W_reg_58_29,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_57_29,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_56_29,
   O => T1_31_i_77_n_0
);
T1_31_i_78 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_51_29,
   I1 => W_reg_50_29,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_49_29,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_48_29,
   O => T1_31_i_78_n_0
);
T1_31_i_79 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_55_29,
   I1 => W_reg_54_29,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_53_29,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_52_29,
   O => T1_31_i_79_n_0
);
T1_31_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => T1_31_i_4_n_0,
   I1 => T1_reg_31_i_10_n_6,
   I2 => T1_31_i_11_n_0,
   I3 => ROTR11_out_3,
   I4 => ROTR11_out_21,
   I5 => ROTR11_out_8,
   O => T1_31_i_8_n_0
);
T1_31_i_80 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_43_29,
   I1 => W_reg_42_29,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_41_29,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_40_29,
   O => T1_31_i_80_n_0
);
T1_31_i_81 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_47_29,
   I1 => W_reg_46_29,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_45_29,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_44_29,
   O => T1_31_i_81_n_0
);
T1_31_i_82 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_35_29,
   I1 => W_reg_34_29,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_33_29,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_32_29,
   O => T1_31_i_82_n_0
);
T1_31_i_83 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_39_29,
   I1 => W_reg_38_29,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_37_29,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_36_29,
   O => T1_31_i_83_n_0
);
T1_31_i_84 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_31_29,
   I1 => W_reg_30_29,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_29_29,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_28_29,
   O => T1_31_i_84_n_0
);
T1_31_i_85 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_27_29,
   I1 => W_reg_26_29,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_25_29,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_24_29,
   O => T1_31_i_85_n_0
);
T1_31_i_86 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_23_29,
   I1 => W_reg_22_29,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_21_29,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_20_29,
   O => T1_31_i_86_n_0
);
T1_31_i_87 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_19_29,
   I1 => W_reg_18_29,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_17_29,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_16_29,
   O => T1_31_i_87_n_0
);
T1_31_i_88 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_15_29,
   I1 => W_reg_14_29,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_13_29,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_12_29,
   O => T1_31_i_88_n_0
);
T1_31_i_89 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_11_29,
   I1 => W_reg_10_29,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_9_29,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_8_29,
   O => T1_31_i_89_n_0
);
T1_31_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => T1_31_i_5_n_0,
   I1 => ROTR11_out_4,
   I2 => ROTR11_out_22,
   I3 => ROTR11_out_9,
   I4 => T1_reg_31_i_10_n_7,
   I5 => T1_31_i_12_n_0,
   O => T1_31_i_9_n_0
);
T1_31_i_90 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_7_29,
   I1 => W_reg_6_29,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_5_29,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_4_29,
   O => T1_31_i_90_n_0
);
T1_31_i_91 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_3_29,
   I1 => W_reg_2_29,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_1_29,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_0_29,
   O => T1_31_i_91_n_0
);
T1_31_i_92 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_59_28,
   I1 => W_reg_58_28,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_57_28,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_56_28,
   O => T1_31_i_92_n_0
);
T1_31_i_93 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_63_28,
   I1 => W_reg_62_28,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_61_28,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_60_28,
   O => T1_31_i_93_n_0
);
T1_31_i_94 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_51_28,
   I1 => W_reg_50_28,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_49_28,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_48_28,
   O => T1_31_i_94_n_0
);
T1_31_i_95 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_55_28,
   I1 => W_reg_54_28,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_53_28,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_52_28,
   O => T1_31_i_95_n_0
);
T1_31_i_98 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_27_28,
   I1 => W_reg_26_28,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_25_28,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_24_28,
   O => T1_31_i_98_n_0
);
T1_31_i_99 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_31_28,
   I1 => W_reg_30_28,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_29_28,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_28_28,
   O => T1_31_i_99_n_0
);
T1_3_i_10 : LUT3
  generic map(
   INIT => X"b8"
  )
 port map (
   I0 => f_reg_n_0_1,
   I1 => ROTR11_out_10,
   I2 => g_reg_n_0_1,
   O => T1_3_i_10_n_0
);
T1_3_i_11 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => ROTR11_out_5,
   I1 => ROTR11_out_32,
   I2 => ROTR11_out_18,
   O => T1_3_i_11_n_0
);
T1_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => ROTR11_out_3,
   I1 => ROTR11_out_30,
   I2 => ROTR11_out_16,
   I3 => T1_reg_7_i_13_n_5,
   I4 => T1_3_i_9_n_0,
   O => T1_3_i_2_n_0
);
T1_3_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => ROTR11_out_4,
   I1 => ROTR11_out_31,
   I2 => ROTR11_out_17,
   I3 => T1_reg_7_i_13_n_6,
   I4 => T1_3_i_10_n_0,
   O => T1_3_i_3_n_0
);
T1_3_i_4 : LUT5
  generic map(
   INIT => X"ffb8b800"
  )
 port map (
   I0 => f_reg_n_0_0,
   I1 => ROTR11_out_11,
   I2 => g_reg_n_0_0,
   I3 => T1_reg_7_i_13_n_7,
   I4 => T1_3_i_11_n_0,
   O => T1_3_i_4_n_0
);
T1_3_i_5 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => T1_3_i_2_n_0,
   I1 => T1_reg_7_i_13_n_4,
   I2 => T1_7_i_14_n_0,
   I3 => ROTR11_out_29,
   I4 => ROTR11_out_15,
   I5 => ROTR11_out_2,
   O => T1_3_i_5_n_0
);
T1_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => T1_3_i_3_n_0,
   I1 => T1_reg_7_i_13_n_5,
   I2 => T1_3_i_9_n_0,
   I3 => ROTR11_out_3,
   I4 => ROTR11_out_30,
   I5 => ROTR11_out_16,
   O => T1_3_i_6_n_0
);
T1_3_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => T1_3_i_4_n_0,
   I1 => T1_reg_7_i_13_n_6,
   I2 => T1_3_i_10_n_0,
   I3 => ROTR11_out_4,
   I4 => ROTR11_out_31,
   I5 => ROTR11_out_17,
   O => T1_3_i_7_n_0
);
T1_3_i_8 : LUT5
  generic map(
   INIT => X"b84747b8"
  )
 port map (
   I0 => f_reg_n_0_0,
   I1 => ROTR11_out_11,
   I2 => g_reg_n_0_0,
   I3 => T1_reg_7_i_13_n_7,
   I4 => T1_3_i_11_n_0,
   O => T1_3_i_8_n_0
);
T1_3_i_9 : LUT3
  generic map(
   INIT => X"b8"
  )
 port map (
   I0 => f_reg_n_0_2,
   I1 => ROTR11_out_9,
   I2 => g_reg_n_0_2,
   O => T1_3_i_9_n_0
);
T1_7_i_10 : LUT3
  generic map(
   INIT => X"b8"
  )
 port map (
   I0 => f_reg_n_0_6,
   I1 => ROTR11_out_5,
   I2 => g_reg_n_0_6,
   O => T1_7_i_10_n_0
);
T1_7_i_11 : LUT3
  generic map(
   INIT => X"b8"
  )
 port map (
   I0 => f_reg_n_0_5,
   I1 => ROTR11_out_6,
   I2 => g_reg_n_0_5,
   O => T1_7_i_11_n_0
);
T1_7_i_12 : LUT3
  generic map(
   INIT => X"b8"
  )
 port map (
   I0 => f_reg_n_0_4,
   I1 => ROTR11_out_7,
   I2 => g_reg_n_0_4,
   O => T1_7_i_12_n_0
);
T1_7_i_14 : LUT3
  generic map(
   INIT => X"b8"
  )
 port map (
   I0 => f_reg_n_0_3,
   I1 => ROTR11_out_8,
   I2 => g_reg_n_0_3,
   O => T1_7_i_14_n_0
);
T1_7_i_15 : LUT3
  generic map(
   INIT => X"e8"
  )
 port map (
   I0 => g0_b2_n_0,
   I1 => T1_7_i_22_n_0,
   I2 => h_2,
   O => T1_7_i_15_n_0
);
T1_7_i_16 : LUT3
  generic map(
   INIT => X"e8"
  )
 port map (
   I0 => g0_b1_n_0,
   I1 => T1_7_i_23_n_0,
   I2 => h_1,
   O => T1_7_i_16_n_0
);
T1_7_i_17 : LUT3
  generic map(
   INIT => X"e8"
  )
 port map (
   I0 => g0_b0_n_0,
   I1 => T1_7_i_24_n_0,
   I2 => h_0,
   O => T1_7_i_17_n_0
);
T1_7_i_18 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => g0_b3_n_0,
   I1 => T1_11_i_26_n_0,
   I2 => h_3,
   I3 => T1_7_i_15_n_0,
   O => T1_7_i_18_n_0
);
T1_7_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => g0_b2_n_0,
   I1 => T1_7_i_22_n_0,
   I2 => h_2,
   I3 => T1_7_i_16_n_0,
   O => T1_7_i_19_n_0
);
T1_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => ROTR11_out_12,
   I1 => ROTR11_out_26,
   I2 => ROTR11_out_31,
   I3 => T1_reg_11_i_13_n_5,
   I4 => T1_7_i_10_n_0,
   O => T1_7_i_2_n_0
);
T1_7_i_20 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => g0_b1_n_0,
   I1 => T1_7_i_23_n_0,
   I2 => h_1,
   I3 => T1_7_i_17_n_0,
   O => T1_7_i_20_n_0
);
T1_7_i_21 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => g0_b0_n_0,
   I1 => T1_7_i_24_n_0,
   I2 => h_0,
   O => T1_7_i_21_n_0
);
T1_7_i_22 : LUT6
  generic map(
   INIT => X"303f303f50505f5f"
  )
 port map (
   I0 => T1_7_i_25_n_0,
   I1 => T1_7_i_26_n_0,
   I2 => HASH_02_COUNTER_5,
   I3 => T1_7_i_27_n_0,
   I4 => T1_7_i_28_n_0,
   I5 => HASH_02_COUNTER_4,
   O => T1_7_i_22_n_0
);
T1_7_i_23 : LUT6
  generic map(
   INIT => X"505f505f30303f3f"
  )
 port map (
   I0 => T1_7_i_29_n_0,
   I1 => T1_7_i_30_n_0,
   I2 => HASH_02_COUNTER_5,
   I3 => T1_7_i_31_n_0,
   I4 => T1_7_i_32_n_0,
   I5 => HASH_02_COUNTER_4,
   O => T1_7_i_23_n_0
);
T1_7_i_24 : LUT6
  generic map(
   INIT => X"303f303f50505f5f"
  )
 port map (
   I0 => T1_7_i_33_n_0,
   I1 => T1_7_i_34_n_0,
   I2 => HASH_02_COUNTER_5,
   I3 => T1_7_i_35_n_0,
   I4 => T1_7_i_36_n_0,
   I5 => HASH_02_COUNTER_4,
   O => T1_7_i_24_n_0
);
T1_7_i_25 : LUT6
  generic map(
   INIT => X"5050303f5f5f303f"
  )
 port map (
   I0 => T1_7_i_37_n_0,
   I1 => T1_7_i_38_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_7_i_39_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_7_i_40_n_0,
   O => T1_7_i_25_n_0
);
T1_7_i_26 : LUT6
  generic map(
   INIT => X"303f5050303f5f5f"
  )
 port map (
   I0 => T1_7_i_41_n_0,
   I1 => T1_7_i_42_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_7_i_43_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_7_i_44_n_0,
   O => T1_7_i_26_n_0
);
T1_7_i_27 : LUT6
  generic map(
   INIT => X"3030505f3f3f505f"
  )
 port map (
   I0 => T1_7_i_45_n_0,
   I1 => T1_7_i_46_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_7_i_47_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_7_i_48_n_0,
   O => T1_7_i_27_n_0
);
T1_7_i_28 : LUT6
  generic map(
   INIT => X"505f3030505f3f3f"
  )
 port map (
   I0 => T1_7_i_49_n_0,
   I1 => T1_7_i_50_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_7_i_51_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_7_i_52_n_0,
   O => T1_7_i_28_n_0
);
T1_7_i_29 : LUT6
  generic map(
   INIT => X"303f5050303f5f5f"
  )
 port map (
   I0 => T1_7_i_53_n_0,
   I1 => T1_7_i_54_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_7_i_55_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_7_i_56_n_0,
   O => T1_7_i_29_n_0
);
T1_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => ROTR11_out_32,
   I1 => ROTR11_out_27,
   I2 => ROTR11_out_13,
   I3 => T1_reg_11_i_13_n_6,
   I4 => T1_7_i_11_n_0,
   O => T1_7_i_3_n_0
);
T1_7_i_30 : LUT6
  generic map(
   INIT => X"5050303f5f5f303f"
  )
 port map (
   I0 => T1_7_i_57_n_0,
   I1 => T1_7_i_58_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_7_i_59_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_7_i_60_n_0,
   O => T1_7_i_30_n_0
);
T1_7_i_31 : LUT6
  generic map(
   INIT => X"5050303f5f5f303f"
  )
 port map (
   I0 => T1_7_i_61_n_0,
   I1 => T1_7_i_62_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_7_i_63_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_7_i_64_n_0,
   O => T1_7_i_31_n_0
);
T1_7_i_32 : LUT6
  generic map(
   INIT => X"5050303f5f5f303f"
  )
 port map (
   I0 => T1_7_i_65_n_0,
   I1 => T1_7_i_66_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_7_i_67_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_7_i_68_n_0,
   O => T1_7_i_32_n_0
);
T1_7_i_33 : LUT6
  generic map(
   INIT => X"5050303f5f5f303f"
  )
 port map (
   I0 => T1_7_i_69_n_0,
   I1 => T1_7_i_70_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_7_i_71_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_7_i_72_n_0,
   O => T1_7_i_33_n_0
);
T1_7_i_34 : LUT6
  generic map(
   INIT => X"303f5050303f5f5f"
  )
 port map (
   I0 => T1_7_i_73_n_0,
   I1 => T1_7_i_74_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_7_i_75_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_7_i_76_n_0,
   O => T1_7_i_34_n_0
);
T1_7_i_35 : LUT6
  generic map(
   INIT => X"3030505f3f3f505f"
  )
 port map (
   I0 => T1_7_i_77_n_0,
   I1 => T1_7_i_78_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_7_i_79_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_7_i_80_n_0,
   O => T1_7_i_35_n_0
);
T1_7_i_36 : LUT6
  generic map(
   INIT => X"303f5050303f5f5f"
  )
 port map (
   I0 => T1_7_i_81_n_0,
   I1 => T1_7_i_82_n_0,
   I2 => HASH_02_COUNTER_3,
   I3 => T1_7_i_83_n_0,
   I4 => HASH_02_COUNTER_2,
   I5 => T1_7_i_84_n_0,
   O => T1_7_i_36_n_0
);
T1_7_i_37 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_47_2,
   I1 => W_reg_46_2,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_45_2,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_44_2,
   O => T1_7_i_37_n_0
);
T1_7_i_38 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_43_2,
   I1 => W_reg_42_2,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_41_2,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_40_2,
   O => T1_7_i_38_n_0
);
T1_7_i_39 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_35_2,
   I1 => W_reg_34_2,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_33_2,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_32_2,
   O => T1_7_i_39_n_0
);
T1_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => ROTR11_out_1,
   I1 => ROTR11_out_28,
   I2 => ROTR11_out_14,
   I3 => T1_reg_11_i_13_n_7,
   I4 => T1_7_i_12_n_0,
   O => T1_7_i_4_n_0
);
T1_7_i_40 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_39_2,
   I1 => W_reg_38_2,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_37_2,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_36_2,
   O => T1_7_i_40_n_0
);
T1_7_i_41 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_59_2,
   I1 => W_reg_58_2,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_57_2,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_56_2,
   O => T1_7_i_41_n_0
);
T1_7_i_42 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_63_2,
   I1 => W_reg_62_2,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_61_2,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_60_2,
   O => T1_7_i_42_n_0
);
T1_7_i_43 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_55_2,
   I1 => W_reg_54_2,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_53_2,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_52_2,
   O => T1_7_i_43_n_0
);
T1_7_i_44 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_51_2,
   I1 => W_reg_50_2,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_49_2,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_48_2,
   O => T1_7_i_44_n_0
);
T1_7_i_45 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_27_2,
   I1 => W_reg_26_2,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_25_2,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_24_2,
   O => T1_7_i_45_n_0
);
T1_7_i_46 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_31_2,
   I1 => W_reg_30_2,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_29_2,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_28_2,
   O => T1_7_i_46_n_0
);
T1_7_i_47 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_19_2,
   I1 => W_reg_18_2,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_17_2,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_16_2,
   O => T1_7_i_47_n_0
);
T1_7_i_48 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_23_2,
   I1 => W_reg_22_2,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_21_2,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_20_2,
   O => T1_7_i_48_n_0
);
T1_7_i_49 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_15_2,
   I1 => W_reg_14_2,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_13_2,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_12_2,
   O => T1_7_i_49_n_0
);
T1_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => ROTR11_out_29,
   I1 => ROTR11_out_15,
   I2 => ROTR11_out_2,
   I3 => T1_reg_7_i_13_n_4,
   I4 => T1_7_i_14_n_0,
   O => T1_7_i_5_n_0
);
T1_7_i_50 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_11_2,
   I1 => W_reg_10_2,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_9_2,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_8_2,
   O => T1_7_i_50_n_0
);
T1_7_i_51 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_7_2,
   I1 => W_reg_6_2,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_5_2,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_4_2,
   O => T1_7_i_51_n_0
);
T1_7_i_52 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_3_2,
   I1 => W_reg_2_2,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_1_2,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_0_2,
   O => T1_7_i_52_n_0
);
T1_7_i_53 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_59_1,
   I1 => W_reg_58_1,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_57_1,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_56_1,
   O => T1_7_i_53_n_0
);
T1_7_i_54 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_63_1,
   I1 => W_reg_62_1,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_61_1,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_60_1,
   O => T1_7_i_54_n_0
);
T1_7_i_55 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_55_1,
   I1 => W_reg_54_1,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_53_1,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_52_1,
   O => T1_7_i_55_n_0
);
T1_7_i_56 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_51_1,
   I1 => W_reg_50_1,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_49_1,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_48_1,
   O => T1_7_i_56_n_0
);
T1_7_i_57 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_47_1,
   I1 => W_reg_46_1,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_45_1,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_44_1,
   O => T1_7_i_57_n_0
);
T1_7_i_58 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_43_1,
   I1 => W_reg_42_1,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_41_1,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_40_1,
   O => T1_7_i_58_n_0
);
T1_7_i_59 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_35_1,
   I1 => W_reg_34_1,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_33_1,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_32_1,
   O => T1_7_i_59_n_0
);
T1_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => T1_7_i_2_n_0,
   I1 => T1_reg_11_i_13_n_4,
   I2 => T1_11_i_14_n_0,
   I3 => ROTR11_out_25,
   I4 => ROTR11_out_11,
   I5 => ROTR11_out_30,
   O => T1_7_i_6_n_0
);
T1_7_i_60 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_39_1,
   I1 => W_reg_38_1,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_37_1,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_36_1,
   O => T1_7_i_60_n_0
);
T1_7_i_61 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_31_1,
   I1 => W_reg_30_1,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_29_1,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_28_1,
   O => T1_7_i_61_n_0
);
T1_7_i_62 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_27_1,
   I1 => W_reg_26_1,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_25_1,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_24_1,
   O => T1_7_i_62_n_0
);
T1_7_i_63 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_19_1,
   I1 => W_reg_18_1,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_17_1,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_16_1,
   O => T1_7_i_63_n_0
);
T1_7_i_64 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_23_1,
   I1 => W_reg_22_1,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_21_1,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_20_1,
   O => T1_7_i_64_n_0
);
T1_7_i_65 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_15_1,
   I1 => W_reg_14_1,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_13_1,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_12_1,
   O => T1_7_i_65_n_0
);
T1_7_i_66 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_11_1,
   I1 => W_reg_10_1,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_9_1,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_8_1,
   O => T1_7_i_66_n_0
);
T1_7_i_67 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_3_1,
   I1 => W_reg_2_1,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_1_1,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_0_1,
   O => T1_7_i_67_n_0
);
T1_7_i_68 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_7_1,
   I1 => W_reg_6_1,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_5_1,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_4_1,
   O => T1_7_i_68_n_0
);
T1_7_i_69 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_47_0,
   I1 => W_reg_46_0,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_45_0,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_44_0,
   O => T1_7_i_69_n_0
);
T1_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => T1_7_i_3_n_0,
   I1 => T1_reg_11_i_13_n_5,
   I2 => T1_7_i_10_n_0,
   I3 => ROTR11_out_12,
   I4 => ROTR11_out_26,
   I5 => ROTR11_out_31,
   O => T1_7_i_7_n_0
);
T1_7_i_70 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_43_0,
   I1 => W_reg_42_0,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_41_0,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_40_0,
   O => T1_7_i_70_n_0
);
T1_7_i_71 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_35_0,
   I1 => W_reg_34_0,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_33_0,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_32_0,
   O => T1_7_i_71_n_0
);
T1_7_i_72 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_39_0,
   I1 => W_reg_38_0,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_37_0,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_36_0,
   O => T1_7_i_72_n_0
);
T1_7_i_73 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_59_0,
   I1 => W_reg_58_0,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_57_0,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_56_0,
   O => T1_7_i_73_n_0
);
T1_7_i_74 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_63_0,
   I1 => W_reg_62_0,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_61_0,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_60_0,
   O => T1_7_i_74_n_0
);
T1_7_i_75 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_55_0,
   I1 => W_reg_54_0,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_53_0,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_52_0,
   O => T1_7_i_75_n_0
);
T1_7_i_76 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_51_0,
   I1 => W_reg_50_0,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_49_0,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_48_0,
   O => T1_7_i_76_n_0
);
T1_7_i_77 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_27_0,
   I1 => W_reg_26_0,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_25_0,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_24_0,
   O => T1_7_i_77_n_0
);
T1_7_i_78 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_31_0,
   I1 => W_reg_30_0,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_29_0,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_28_0,
   O => T1_7_i_78_n_0
);
T1_7_i_79 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_19_0,
   I1 => W_reg_18_0,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_17_0,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_16_0,
   O => T1_7_i_79_n_0
);
T1_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => T1_7_i_4_n_0,
   I1 => ROTR11_out_32,
   I2 => ROTR11_out_27,
   I3 => ROTR11_out_13,
   I4 => T1_reg_11_i_13_n_6,
   I5 => T1_7_i_11_n_0,
   O => T1_7_i_8_n_0
);
T1_7_i_80 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_23_0,
   I1 => W_reg_22_0,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_21_0,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_20_0,
   O => T1_7_i_80_n_0
);
T1_7_i_81 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_11_0,
   I1 => W_reg_10_0,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_9_0,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_8_0,
   O => T1_7_i_81_n_0
);
T1_7_i_82 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_15_0,
   I1 => W_reg_14_0,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_13_0,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_12_0,
   O => T1_7_i_82_n_0
);
T1_7_i_83 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_7_0,
   I1 => W_reg_6_0,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_5_0,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_4_0,
   O => T1_7_i_83_n_0
);
T1_7_i_84 : LUT6
  generic map(
   INIT => X"afa0cfcfafa0c0c0"
  )
 port map (
   I0 => W_reg_3_0,
   I1 => W_reg_2_0,
   I2 => HASH_02_COUNTER_1,
   I3 => W_reg_1_0,
   I4 => HASH_02_COUNTER_0,
   I5 => W_reg_0_0,
   O => T1_7_i_84_n_0
);
T1_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => T1_7_i_5_n_0,
   I1 => ROTR11_out_1,
   I2 => ROTR11_out_28,
   I3 => ROTR11_out_14,
   I4 => T1_reg_11_i_13_n_7,
   I5 => T1_7_i_12_n_0,
   O => T1_7_i_9_n_0
);
T1_reg_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T100_in_0,
   R => '0',
   Q => T1_0_0
);
T1_reg_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T100_in_10,
   R => '0',
   Q => T1_0_10
);
T1_reg_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T100_in_11,
   R => '0',
   Q => T1_0_11
);
T1_reg_11_i_1 : CARRY4
 port map (
   CI => T1_reg_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => T1_11_i_5_n_0,
   DI(1) => T1_11_i_4_n_0,
   DI(2) => T1_11_i_3_n_0,
   DI(3) => T1_11_i_2_n_0,
   S(0) => T1_11_i_9_n_0,
   S(1) => T1_11_i_8_n_0,
   S(2) => T1_11_i_7_n_0,
   S(3) => T1_11_i_6_n_0,
   CO(0) => T1_reg_11_i_1_n_3,
   CO(1) => T1_reg_11_i_1_n_2,
   CO(2) => T1_reg_11_i_1_n_1,
   CO(3) => T1_reg_11_i_1_n_0,
   O(0) => T100_in_8,
   O(1) => T100_in_9,
   O(2) => T100_in_10,
   O(3) => T100_in_11
);
T1_reg_11_i_13 : CARRY4
 port map (
   CI => T1_reg_7_i_13_n_0,
   CYINIT => '0',
   DI(0) => T1_11_i_18_n_0,
   DI(1) => T1_11_i_17_n_0,
   DI(2) => T1_11_i_16_n_0,
   DI(3) => T1_11_i_15_n_0,
   S(0) => T1_11_i_22_n_0,
   S(1) => T1_11_i_21_n_0,
   S(2) => T1_11_i_20_n_0,
   S(3) => T1_11_i_19_n_0,
   CO(0) => T1_reg_11_i_13_n_3,
   CO(1) => T1_reg_11_i_13_n_2,
   CO(2) => T1_reg_11_i_13_n_1,
   CO(3) => T1_reg_11_i_13_n_0,
   O(0) => T1_reg_11_i_13_n_7,
   O(1) => T1_reg_11_i_13_n_6,
   O(2) => T1_reg_11_i_13_n_5,
   O(3) => T1_reg_11_i_13_n_4
);
T1_reg_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T100_in_12,
   R => '0',
   Q => T1_0_12
);
T1_reg_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T100_in_13,
   R => '0',
   Q => T1_0_13
);
T1_reg_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T100_in_14,
   R => '0',
   Q => T1_0_14
);
T1_reg_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T100_in_15,
   R => '0',
   Q => T1_0_15
);
T1_reg_15_i_1 : CARRY4
 port map (
   CI => T1_reg_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => T1_15_i_5_n_0,
   DI(1) => T1_15_i_4_n_0,
   DI(2) => T1_15_i_3_n_0,
   DI(3) => T1_15_i_2_n_0,
   S(0) => T1_15_i_9_n_0,
   S(1) => T1_15_i_8_n_0,
   S(2) => T1_15_i_7_n_0,
   S(3) => T1_15_i_6_n_0,
   CO(0) => T1_reg_15_i_1_n_3,
   CO(1) => T1_reg_15_i_1_n_2,
   CO(2) => T1_reg_15_i_1_n_1,
   CO(3) => T1_reg_15_i_1_n_0,
   O(0) => T100_in_12,
   O(1) => T100_in_13,
   O(2) => T100_in_14,
   O(3) => T100_in_15
);
T1_reg_15_i_13 : CARRY4
 port map (
   CI => T1_reg_11_i_13_n_0,
   CYINIT => '0',
   DI(0) => T1_15_i_18_n_0,
   DI(1) => T1_15_i_17_n_0,
   DI(2) => T1_15_i_16_n_0,
   DI(3) => T1_15_i_15_n_0,
   S(0) => T1_15_i_22_n_0,
   S(1) => T1_15_i_21_n_0,
   S(2) => T1_15_i_20_n_0,
   S(3) => T1_15_i_19_n_0,
   CO(0) => T1_reg_15_i_13_n_3,
   CO(1) => T1_reg_15_i_13_n_2,
   CO(2) => T1_reg_15_i_13_n_1,
   CO(3) => T1_reg_15_i_13_n_0,
   O(0) => T1_reg_15_i_13_n_7,
   O(1) => T1_reg_15_i_13_n_6,
   O(2) => T1_reg_15_i_13_n_5,
   O(3) => T1_reg_15_i_13_n_4
);
T1_reg_15_i_29 : MUXF8
 port map (
   I0 => T1_reg_15_i_51_n_0,
   I1 => T1_reg_15_i_52_n_0,
   S => HASH_02_COUNTER_3,
   O => T1_reg_15_i_29_n_0
);
T1_reg_15_i_33 : MUXF8
 port map (
   I0 => T1_reg_15_i_65_n_0,
   I1 => T1_reg_15_i_66_n_0,
   S => HASH_02_COUNTER_3,
   O => T1_reg_15_i_33_n_0
);
T1_reg_15_i_37 : MUXF8
 port map (
   I0 => T1_reg_15_i_79_n_0,
   I1 => T1_reg_15_i_80_n_0,
   S => HASH_02_COUNTER_3,
   O => T1_reg_15_i_37_n_0
);
T1_reg_15_i_51 : MUXF7
 port map (
   I0 => T1_15_i_101_n_0,
   I1 => T1_15_i_102_n_0,
   S => HASH_02_COUNTER_2,
   O => T1_reg_15_i_51_n_0
);
T1_reg_15_i_52 : MUXF7
 port map (
   I0 => T1_15_i_103_n_0,
   I1 => T1_15_i_104_n_0,
   S => HASH_02_COUNTER_2,
   O => T1_reg_15_i_52_n_0
);
T1_reg_15_i_65 : MUXF7
 port map (
   I0 => T1_15_i_105_n_0,
   I1 => T1_15_i_106_n_0,
   S => HASH_02_COUNTER_2,
   O => T1_reg_15_i_65_n_0
);
T1_reg_15_i_66 : MUXF7
 port map (
   I0 => T1_15_i_107_n_0,
   I1 => T1_15_i_108_n_0,
   S => HASH_02_COUNTER_2,
   O => T1_reg_15_i_66_n_0
);
T1_reg_15_i_79 : MUXF7
 port map (
   I0 => T1_15_i_109_n_0,
   I1 => T1_15_i_110_n_0,
   S => HASH_02_COUNTER_2,
   O => T1_reg_15_i_79_n_0
);
T1_reg_15_i_80 : MUXF7
 port map (
   I0 => T1_15_i_111_n_0,
   I1 => T1_15_i_112_n_0,
   S => HASH_02_COUNTER_2,
   O => T1_reg_15_i_80_n_0
);
T1_reg_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T100_in_16,
   R => '0',
   Q => T1_0_16
);
T1_reg_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T100_in_17,
   R => '0',
   Q => T1_0_17
);
T1_reg_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T100_in_18,
   R => '0',
   Q => T1_0_18
);
T1_reg_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T100_in_19,
   R => '0',
   Q => T1_0_19
);
T1_reg_19_i_1 : CARRY4
 port map (
   CI => T1_reg_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => T1_19_i_5_n_0,
   DI(1) => T1_19_i_4_n_0,
   DI(2) => T1_19_i_3_n_0,
   DI(3) => T1_19_i_2_n_0,
   S(0) => T1_19_i_9_n_0,
   S(1) => T1_19_i_8_n_0,
   S(2) => T1_19_i_7_n_0,
   S(3) => T1_19_i_6_n_0,
   CO(0) => T1_reg_19_i_1_n_3,
   CO(1) => T1_reg_19_i_1_n_2,
   CO(2) => T1_reg_19_i_1_n_1,
   CO(3) => T1_reg_19_i_1_n_0,
   O(0) => T100_in_16,
   O(1) => T100_in_17,
   O(2) => T100_in_18,
   O(3) => T100_in_19
);
T1_reg_19_i_100 : MUXF7
 port map (
   I0 => T1_19_i_107_n_0,
   I1 => T1_19_i_108_n_0,
   S => HASH_02_COUNTER_2,
   O => T1_reg_19_i_100_n_0
);
T1_reg_19_i_13 : CARRY4
 port map (
   CI => T1_reg_15_i_13_n_0,
   CYINIT => '0',
   DI(0) => T1_19_i_18_n_0,
   DI(1) => T1_19_i_17_n_0,
   DI(2) => T1_19_i_16_n_0,
   DI(3) => T1_19_i_15_n_0,
   S(0) => T1_19_i_22_n_0,
   S(1) => T1_19_i_21_n_0,
   S(2) => T1_19_i_20_n_0,
   S(3) => T1_19_i_19_n_0,
   CO(0) => T1_reg_19_i_13_n_3,
   CO(1) => T1_reg_19_i_13_n_2,
   CO(2) => T1_reg_19_i_13_n_1,
   CO(3) => T1_reg_19_i_13_n_0,
   O(0) => T1_reg_19_i_13_n_7,
   O(1) => T1_reg_19_i_13_n_6,
   O(2) => T1_reg_19_i_13_n_5,
   O(3) => T1_reg_19_i_13_n_4
);
T1_reg_19_i_41 : MUXF8
 port map (
   I0 => T1_reg_19_i_99_n_0,
   I1 => T1_reg_19_i_100_n_0,
   S => HASH_02_COUNTER_3,
   O => T1_reg_19_i_41_n_0
);
T1_reg_19_i_99 : MUXF7
 port map (
   I0 => T1_19_i_105_n_0,
   I1 => T1_19_i_106_n_0,
   S => HASH_02_COUNTER_2,
   O => T1_reg_19_i_99_n_0
);
T1_reg_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T100_in_1,
   R => '0',
   Q => T1_0_1
);
T1_reg_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T100_in_20,
   R => '0',
   Q => T1_0_20
);
T1_reg_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T100_in_21,
   R => '0',
   Q => T1_0_21
);
T1_reg_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T100_in_22,
   R => '0',
   Q => T1_0_22
);
T1_reg_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T100_in_23,
   R => '0',
   Q => T1_0_23
);
T1_reg_23_i_1 : CARRY4
 port map (
   CI => T1_reg_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => T1_23_i_5_n_0,
   DI(1) => T1_23_i_4_n_0,
   DI(2) => T1_23_i_3_n_0,
   DI(3) => T1_23_i_2_n_0,
   S(0) => T1_23_i_9_n_0,
   S(1) => T1_23_i_8_n_0,
   S(2) => T1_23_i_7_n_0,
   S(3) => T1_23_i_6_n_0,
   CO(0) => T1_reg_23_i_1_n_3,
   CO(1) => T1_reg_23_i_1_n_2,
   CO(2) => T1_reg_23_i_1_n_1,
   CO(3) => T1_reg_23_i_1_n_0,
   O(0) => T100_in_20,
   O(1) => T100_in_21,
   O(2) => T100_in_22,
   O(3) => T100_in_23
);
T1_reg_23_i_13 : CARRY4
 port map (
   CI => T1_reg_19_i_13_n_0,
   CYINIT => '0',
   DI(0) => T1_23_i_18_n_0,
   DI(1) => T1_23_i_17_n_0,
   DI(2) => T1_23_i_16_n_0,
   DI(3) => T1_23_i_15_n_0,
   S(0) => T1_23_i_22_n_0,
   S(1) => T1_23_i_21_n_0,
   S(2) => T1_23_i_20_n_0,
   S(3) => T1_23_i_19_n_0,
   CO(0) => T1_reg_23_i_13_n_3,
   CO(1) => T1_reg_23_i_13_n_2,
   CO(2) => T1_reg_23_i_13_n_1,
   CO(3) => T1_reg_23_i_13_n_0,
   O(0) => T1_reg_23_i_13_n_7,
   O(1) => T1_reg_23_i_13_n_6,
   O(2) => T1_reg_23_i_13_n_5,
   O(3) => T1_reg_23_i_13_n_4
);
T1_reg_23_i_40 : MUXF8
 port map (
   I0 => T1_reg_23_i_95_n_0,
   I1 => T1_reg_23_i_96_n_0,
   S => HASH_02_COUNTER_3,
   O => T1_reg_23_i_40_n_0
);
T1_reg_23_i_95 : MUXF7
 port map (
   I0 => T1_23_i_105_n_0,
   I1 => T1_23_i_106_n_0,
   S => HASH_02_COUNTER_2,
   O => T1_reg_23_i_95_n_0
);
T1_reg_23_i_96 : MUXF7
 port map (
   I0 => T1_23_i_107_n_0,
   I1 => T1_23_i_108_n_0,
   S => HASH_02_COUNTER_2,
   O => T1_reg_23_i_96_n_0
);
T1_reg_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T100_in_24,
   R => '0',
   Q => T1_0_24
);
T1_reg_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T100_in_25,
   R => '0',
   Q => T1_0_25
);
T1_reg_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T100_in_26,
   R => '0',
   Q => T1_0_26
);
T1_reg_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T100_in_27,
   R => '0',
   Q => T1_0_27
);
T1_reg_27_i_1 : CARRY4
 port map (
   CI => T1_reg_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => T1_27_i_5_n_0,
   DI(1) => T1_27_i_4_n_0,
   DI(2) => T1_27_i_3_n_0,
   DI(3) => T1_27_i_2_n_0,
   S(0) => T1_27_i_9_n_0,
   S(1) => T1_27_i_8_n_0,
   S(2) => T1_27_i_7_n_0,
   S(3) => T1_27_i_6_n_0,
   CO(0) => T1_reg_27_i_1_n_3,
   CO(1) => T1_reg_27_i_1_n_2,
   CO(2) => T1_reg_27_i_1_n_1,
   CO(3) => T1_reg_27_i_1_n_0,
   O(0) => T100_in_24,
   O(1) => T100_in_25,
   O(2) => T100_in_26,
   O(3) => T100_in_27
);
T1_reg_27_i_13 : CARRY4
 port map (
   CI => T1_reg_23_i_13_n_0,
   CYINIT => '0',
   DI(0) => T1_27_i_18_n_0,
   DI(1) => T1_27_i_17_n_0,
   DI(2) => T1_27_i_16_n_0,
   DI(3) => T1_27_i_15_n_0,
   S(0) => T1_27_i_22_n_0,
   S(1) => T1_27_i_21_n_0,
   S(2) => T1_27_i_20_n_0,
   S(3) => T1_27_i_19_n_0,
   CO(0) => T1_reg_27_i_13_n_3,
   CO(1) => T1_reg_27_i_13_n_2,
   CO(2) => T1_reg_27_i_13_n_1,
   CO(3) => T1_reg_27_i_13_n_0,
   O(0) => T1_reg_27_i_13_n_7,
   O(1) => T1_reg_27_i_13_n_6,
   O(2) => T1_reg_27_i_13_n_5,
   O(3) => T1_reg_27_i_13_n_4
);
T1_reg_27_i_28 : MUXF8
 port map (
   I0 => T1_reg_27_i_47_n_0,
   I1 => T1_reg_27_i_48_n_0,
   S => HASH_02_COUNTER_3,
   O => T1_reg_27_i_28_n_0
);
T1_reg_27_i_47 : MUXF7
 port map (
   I0 => T1_27_i_105_n_0,
   I1 => T1_27_i_106_n_0,
   S => HASH_02_COUNTER_2,
   O => T1_reg_27_i_47_n_0
);
T1_reg_27_i_48 : MUXF7
 port map (
   I0 => T1_27_i_107_n_0,
   I1 => T1_27_i_108_n_0,
   S => HASH_02_COUNTER_2,
   O => T1_reg_27_i_48_n_0
);
T1_reg_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T100_in_28,
   R => '0',
   Q => T1_0_28
);
T1_reg_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T100_in_29,
   R => '0',
   Q => T1_0_29
);
T1_reg_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T100_in_2,
   R => '0',
   Q => T1_0_2
);
T1_reg_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T100_in_30,
   R => '0',
   Q => T1_0_30
);
T1_reg_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T100_in_31,
   R => '0',
   Q => T1_0_31
);
T1_reg_31_i_10 : CARRY4
 port map (
   CI => T1_reg_31_i_13_n_0,
   CYINIT => '0',
   DI(0) => T1_31_i_20_n_0,
   DI(1) => T1_31_i_19_n_0,
   DI(2) => T1_31_i_18_n_0,
   DI(3) => '0',
   S(0) => T1_31_i_24_n_0,
   S(1) => T1_31_i_23_n_0,
   S(2) => T1_31_i_22_n_0,
   S(3) => T1_31_i_21_n_0,
   CO(0) => T1_reg_31_i_10_n_3,
   CO(1) => T1_reg_31_i_10_n_2,
   CO(2) => T1_reg_31_i_10_n_1,
   CO(3) => NLW_T1_reg_31_i_10_CO_UNCONNECTED_3,
   O(0) => T1_reg_31_i_10_n_7,
   O(1) => T1_reg_31_i_10_n_6,
   O(2) => T1_reg_31_i_10_n_5,
   O(3) => T1_reg_31_i_10_n_4
);
T1_reg_31_i_110 : MUXF7
 port map (
   I0 => T1_31_i_196_n_0,
   I1 => T1_31_i_197_n_0,
   S => HASH_02_COUNTER_2,
   O => T1_reg_31_i_110_n_0
);
T1_reg_31_i_111 : MUXF7
 port map (
   I0 => T1_31_i_198_n_0,
   I1 => T1_31_i_199_n_0,
   S => HASH_02_COUNTER_2,
   O => T1_reg_31_i_111_n_0
);
T1_reg_31_i_120 : MUXF7
 port map (
   I0 => T1_31_i_200_n_0,
   I1 => T1_31_i_201_n_0,
   S => HASH_02_COUNTER_2,
   O => T1_reg_31_i_120_n_0
);
T1_reg_31_i_121 : MUXF7
 port map (
   I0 => T1_31_i_202_n_0,
   I1 => T1_31_i_203_n_0,
   S => HASH_02_COUNTER_2,
   O => T1_reg_31_i_121_n_0
);
T1_reg_31_i_122 : MUXF7
 port map (
   I0 => T1_31_i_204_n_0,
   I1 => T1_31_i_205_n_0,
   S => HASH_02_COUNTER_2,
   O => T1_reg_31_i_122_n_0
);
T1_reg_31_i_123 : MUXF7
 port map (
   I0 => T1_31_i_206_n_0,
   I1 => T1_31_i_207_n_0,
   S => HASH_02_COUNTER_2,
   O => T1_reg_31_i_123_n_0
);
T1_reg_31_i_124 : MUXF7
 port map (
   I0 => T1_31_i_208_n_0,
   I1 => T1_31_i_209_n_0,
   S => HASH_02_COUNTER_2,
   O => T1_reg_31_i_124_n_0
);
T1_reg_31_i_125 : MUXF7
 port map (
   I0 => T1_31_i_210_n_0,
   I1 => T1_31_i_211_n_0,
   S => HASH_02_COUNTER_2,
   O => T1_reg_31_i_125_n_0
);
T1_reg_31_i_126 : MUXF7
 port map (
   I0 => T1_31_i_212_n_0,
   I1 => T1_31_i_213_n_0,
   S => HASH_02_COUNTER_2,
   O => T1_reg_31_i_126_n_0
);
T1_reg_31_i_127 : MUXF7
 port map (
   I0 => T1_31_i_214_n_0,
   I1 => T1_31_i_215_n_0,
   S => HASH_02_COUNTER_2,
   O => T1_reg_31_i_127_n_0
);
T1_reg_31_i_13 : CARRY4
 port map (
   CI => T1_reg_27_i_13_n_0,
   CYINIT => '0',
   DI(0) => T1_31_i_28_n_0,
   DI(1) => T1_31_i_27_n_0,
   DI(2) => T1_31_i_26_n_0,
   DI(3) => T1_31_i_25_n_0,
   S(0) => T1_31_i_32_n_0,
   S(1) => T1_31_i_31_n_0,
   S(2) => T1_31_i_30_n_0,
   S(3) => T1_31_i_29_n_0,
   CO(0) => T1_reg_31_i_13_n_3,
   CO(1) => T1_reg_31_i_13_n_2,
   CO(2) => T1_reg_31_i_13_n_1,
   CO(3) => T1_reg_31_i_13_n_0,
   O(0) => T1_reg_31_i_13_n_7,
   O(1) => T1_reg_31_i_13_n_6,
   O(2) => T1_reg_31_i_13_n_5,
   O(3) => T1_reg_31_i_13_n_4
);
T1_reg_31_i_136 : MUXF7
 port map (
   I0 => T1_31_i_232_n_0,
   I1 => T1_31_i_233_n_0,
   S => HASH_02_COUNTER_2,
   O => T1_reg_31_i_136_n_0
);
T1_reg_31_i_137 : MUXF7
 port map (
   I0 => T1_31_i_234_n_0,
   I1 => T1_31_i_235_n_0,
   S => HASH_02_COUNTER_2,
   O => T1_reg_31_i_137_n_0
);
T1_reg_31_i_150 : MUXF7
 port map (
   I0 => T1_31_i_236_n_0,
   I1 => T1_31_i_237_n_0,
   S => HASH_02_COUNTER_2,
   O => T1_reg_31_i_150_n_0
);
T1_reg_31_i_151 : MUXF7
 port map (
   I0 => T1_31_i_238_n_0,
   I1 => T1_31_i_239_n_0,
   S => HASH_02_COUNTER_2,
   O => T1_reg_31_i_151_n_0
);
T1_reg_31_i_2 : CARRY4
 port map (
   CI => T1_reg_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => T1_31_i_5_n_0,
   DI(1) => T1_31_i_4_n_0,
   DI(2) => T1_31_i_3_n_0,
   DI(3) => '0',
   S(0) => T1_31_i_9_n_0,
   S(1) => T1_31_i_8_n_0,
   S(2) => T1_31_i_7_n_0,
   S(3) => T1_31_i_6_n_0,
   CO(0) => T1_reg_31_i_2_n_3,
   CO(1) => T1_reg_31_i_2_n_2,
   CO(2) => T1_reg_31_i_2_n_1,
   CO(3) => NLW_T1_reg_31_i_2_CO_UNCONNECTED_3,
   O(0) => T100_in_28,
   O(1) => T100_in_29,
   O(2) => T100_in_30,
   O(3) => T100_in_31
);
T1_reg_31_i_37 : MUXF8
 port map (
   I0 => T1_reg_31_i_58_n_0,
   I1 => T1_reg_31_i_59_n_0,
   S => HASH_02_COUNTER_5,
   O => T1_reg_31_i_37_n_0
);
T1_reg_31_i_47 : MUXF8
 port map (
   I0 => T1_reg_31_i_96_n_0,
   I1 => T1_reg_31_i_97_n_0,
   S => HASH_02_COUNTER_3,
   O => T1_reg_31_i_47_n_0
);
T1_reg_31_i_51 : MUXF8
 port map (
   I0 => T1_reg_31_i_110_n_0,
   I1 => T1_reg_31_i_111_n_0,
   S => HASH_02_COUNTER_3,
   O => T1_reg_31_i_51_n_0
);
T1_reg_31_i_54 : MUXF8
 port map (
   I0 => T1_reg_31_i_120_n_0,
   I1 => T1_reg_31_i_121_n_0,
   S => HASH_02_COUNTER_3,
   O => T1_reg_31_i_54_n_0
);
T1_reg_31_i_55 : MUXF8
 port map (
   I0 => T1_reg_31_i_122_n_0,
   I1 => T1_reg_31_i_123_n_0,
   S => HASH_02_COUNTER_3,
   O => T1_reg_31_i_55_n_0
);
T1_reg_31_i_56 : MUXF8
 port map (
   I0 => T1_reg_31_i_124_n_0,
   I1 => T1_reg_31_i_125_n_0,
   S => HASH_02_COUNTER_3,
   O => T1_reg_31_i_56_n_0
);
T1_reg_31_i_57 : MUXF8
 port map (
   I0 => T1_reg_31_i_126_n_0,
   I1 => T1_reg_31_i_127_n_0,
   S => HASH_02_COUNTER_3,
   O => T1_reg_31_i_57_n_0
);
T1_reg_31_i_58 : MUXF7
 port map (
   I0 => T1_31_i_128_n_0,
   I1 => T1_31_i_129_n_0,
   S => HASH_02_COUNTER_4,
   O => T1_reg_31_i_58_n_0
);
T1_reg_31_i_59 : MUXF7
 port map (
   I0 => T1_31_i_130_n_0,
   I1 => T1_31_i_131_n_0,
   S => HASH_02_COUNTER_4,
   O => T1_reg_31_i_59_n_0
);
T1_reg_31_i_61 : MUXF8
 port map (
   I0 => T1_reg_31_i_136_n_0,
   I1 => T1_reg_31_i_137_n_0,
   S => HASH_02_COUNTER_3,
   O => T1_reg_31_i_61_n_0
);
T1_reg_31_i_65 : MUXF8
 port map (
   I0 => T1_reg_31_i_150_n_0,
   I1 => T1_reg_31_i_151_n_0,
   S => HASH_02_COUNTER_3,
   O => T1_reg_31_i_65_n_0
);
T1_reg_31_i_96 : MUXF7
 port map (
   I0 => T1_31_i_192_n_0,
   I1 => T1_31_i_193_n_0,
   S => HASH_02_COUNTER_2,
   O => T1_reg_31_i_96_n_0
);
T1_reg_31_i_97 : MUXF7
 port map (
   I0 => T1_31_i_194_n_0,
   I1 => T1_31_i_195_n_0,
   S => HASH_02_COUNTER_2,
   O => T1_reg_31_i_97_n_0
);
T1_reg_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T100_in_3,
   R => '0',
   Q => T1_0_3
);
T1_reg_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => '0',
   DI(1) => T1_3_i_4_n_0,
   DI(2) => T1_3_i_3_n_0,
   DI(3) => T1_3_i_2_n_0,
   S(0) => T1_3_i_8_n_0,
   S(1) => T1_3_i_7_n_0,
   S(2) => T1_3_i_6_n_0,
   S(3) => T1_3_i_5_n_0,
   CO(0) => T1_reg_3_i_1_n_3,
   CO(1) => T1_reg_3_i_1_n_2,
   CO(2) => T1_reg_3_i_1_n_1,
   CO(3) => T1_reg_3_i_1_n_0,
   O(0) => T100_in_0,
   O(1) => T100_in_1,
   O(2) => T100_in_2,
   O(3) => T100_in_3
);
T1_reg_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T100_in_4,
   R => '0',
   Q => T1_0_4
);
T1_reg_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T100_in_5,
   R => '0',
   Q => T1_0_5
);
T1_reg_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T100_in_6,
   R => '0',
   Q => T1_0_6
);
T1_reg_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T100_in_7,
   R => '0',
   Q => T1_0_7
);
T1_reg_7_i_1 : CARRY4
 port map (
   CI => T1_reg_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => T1_7_i_5_n_0,
   DI(1) => T1_7_i_4_n_0,
   DI(2) => T1_7_i_3_n_0,
   DI(3) => T1_7_i_2_n_0,
   S(0) => T1_7_i_9_n_0,
   S(1) => T1_7_i_8_n_0,
   S(2) => T1_7_i_7_n_0,
   S(3) => T1_7_i_6_n_0,
   CO(0) => T1_reg_7_i_1_n_3,
   CO(1) => T1_reg_7_i_1_n_2,
   CO(2) => T1_reg_7_i_1_n_1,
   CO(3) => T1_reg_7_i_1_n_0,
   O(0) => T100_in_4,
   O(1) => T100_in_5,
   O(2) => T100_in_6,
   O(3) => T100_in_7
);
T1_reg_7_i_13 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => '0',
   DI(1) => T1_7_i_17_n_0,
   DI(2) => T1_7_i_16_n_0,
   DI(3) => T1_7_i_15_n_0,
   S(0) => T1_7_i_21_n_0,
   S(1) => T1_7_i_20_n_0,
   S(2) => T1_7_i_19_n_0,
   S(3) => T1_7_i_18_n_0,
   CO(0) => T1_reg_7_i_13_n_3,
   CO(1) => T1_reg_7_i_13_n_2,
   CO(2) => T1_reg_7_i_13_n_1,
   CO(3) => T1_reg_7_i_13_n_0,
   O(0) => T1_reg_7_i_13_n_7,
   O(1) => T1_reg_7_i_13_n_6,
   O(2) => T1_reg_7_i_13_n_5,
   O(3) => T1_reg_7_i_13_n_4
);
T1_reg_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T100_in_8,
   R => '0',
   Q => T1_0_8
);
T1_reg_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T100_in_9,
   R => '0',
   Q => T1_0_9
);
T2_11_i_2 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => ROTR2_out_21,
   I1 => ROTR2_out_12,
   I2 => ROTR2_out_32,
   O => SIGMA_UCASE_0_11
);
T2_11_i_3 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => ROTR2_out_22,
   I1 => ROTR2_out_13,
   I2 => ROTR2_out_1,
   O => SIGMA_UCASE_0_10
);
T2_11_i_4 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => ROTR2_out_23,
   I1 => ROTR2_out_14,
   I2 => ROTR2_out_2,
   O => SIGMA_UCASE_0_9
);
T2_11_i_5 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => ROTR2_out_24,
   I1 => ROTR2_out_15,
   I2 => ROTR2_out_3,
   O => SIGMA_UCASE_0_8
);
T2_11_i_6 : LUT6
  generic map(
   INIT => X"6969699669969696"
  )
 port map (
   I0 => ROTR2_out_32,
   I1 => ROTR2_out_12,
   I2 => ROTR2_out_21,
   I3 => b_reg_n_0_11,
   I4 => c_reg_n_0_11,
   I5 => ROTR2_out_2,
   O => T2_11_i_6_n_0
);
T2_11_i_7 : LUT6
  generic map(
   INIT => X"6969699669969696"
  )
 port map (
   I0 => ROTR2_out_1,
   I1 => ROTR2_out_13,
   I2 => ROTR2_out_22,
   I3 => b_reg_n_0_10,
   I4 => c_reg_n_0_10,
   I5 => ROTR2_out_3,
   O => T2_11_i_7_n_0
);
T2_11_i_8 : LUT6
  generic map(
   INIT => X"6969699669969696"
  )
 port map (
   I0 => ROTR2_out_2,
   I1 => ROTR2_out_14,
   I2 => ROTR2_out_23,
   I3 => b_reg_n_0_9,
   I4 => c_reg_n_0_9,
   I5 => ROTR2_out_4,
   O => T2_11_i_8_n_0
);
T2_11_i_9 : LUT6
  generic map(
   INIT => X"6969699669969696"
  )
 port map (
   I0 => ROTR2_out_3,
   I1 => ROTR2_out_15,
   I2 => ROTR2_out_24,
   I3 => b_reg_n_0_8,
   I4 => c_reg_n_0_8,
   I5 => ROTR2_out_5,
   O => T2_11_i_9_n_0
);
T2_15_i_2 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => ROTR2_out_17,
   I1 => ROTR2_out_28,
   I2 => ROTR2_out_8,
   O => SIGMA_UCASE_0_15
);
T2_15_i_3 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => ROTR2_out_18,
   I1 => ROTR2_out_29,
   I2 => ROTR2_out_9,
   O => SIGMA_UCASE_0_14
);
T2_15_i_4 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => ROTR2_out_19,
   I1 => ROTR2_out_30,
   I2 => ROTR2_out_10,
   O => SIGMA_UCASE_0_13
);
T2_15_i_5 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => ROTR2_out_20,
   I1 => ROTR2_out_31,
   I2 => ROTR2_out_11,
   O => SIGMA_UCASE_0_12
);
T2_15_i_6 : LUT6
  generic map(
   INIT => X"6969699669969696"
  )
 port map (
   I0 => ROTR2_out_8,
   I1 => ROTR2_out_28,
   I2 => ROTR2_out_17,
   I3 => b_reg_n_0_15,
   I4 => c_reg_n_0_15,
   I5 => ROTR2_out_30,
   O => T2_15_i_6_n_0
);
T2_15_i_7 : LUT6
  generic map(
   INIT => X"6969699669969696"
  )
 port map (
   I0 => ROTR2_out_9,
   I1 => ROTR2_out_29,
   I2 => ROTR2_out_18,
   I3 => b_reg_n_0_14,
   I4 => c_reg_n_0_14,
   I5 => ROTR2_out_31,
   O => T2_15_i_7_n_0
);
T2_15_i_8 : LUT6
  generic map(
   INIT => X"6969699669969696"
  )
 port map (
   I0 => ROTR2_out_10,
   I1 => ROTR2_out_30,
   I2 => ROTR2_out_19,
   I3 => b_reg_n_0_13,
   I4 => c_reg_n_0_13,
   I5 => ROTR2_out_32,
   O => T2_15_i_8_n_0
);
T2_15_i_9 : LUT6
  generic map(
   INIT => X"6969699669969696"
  )
 port map (
   I0 => ROTR2_out_11,
   I1 => ROTR2_out_31,
   I2 => ROTR2_out_20,
   I3 => b_reg_n_0_12,
   I4 => c_reg_n_0_12,
   I5 => ROTR2_out_1,
   O => T2_15_i_9_n_0
);
T2_19_i_2 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => ROTR2_out_13,
   I1 => ROTR2_out_24,
   I2 => ROTR2_out_4,
   O => SIGMA_UCASE_0_19
);
T2_19_i_3 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => ROTR2_out_14,
   I1 => ROTR2_out_25,
   I2 => ROTR2_out_5,
   O => SIGMA_UCASE_0_18
);
T2_19_i_4 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => ROTR2_out_15,
   I1 => ROTR2_out_26,
   I2 => ROTR2_out_6,
   O => SIGMA_UCASE_0_17
);
T2_19_i_5 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => ROTR2_out_16,
   I1 => ROTR2_out_27,
   I2 => ROTR2_out_7,
   O => SIGMA_UCASE_0_16
);
T2_19_i_6 : LUT6
  generic map(
   INIT => X"6969699669969696"
  )
 port map (
   I0 => ROTR2_out_4,
   I1 => ROTR2_out_24,
   I2 => ROTR2_out_13,
   I3 => b_reg_n_0_19,
   I4 => c_reg_n_0_19,
   I5 => ROTR2_out_26,
   O => T2_19_i_6_n_0
);
T2_19_i_7 : LUT6
  generic map(
   INIT => X"6969699669969696"
  )
 port map (
   I0 => ROTR2_out_5,
   I1 => ROTR2_out_25,
   I2 => ROTR2_out_14,
   I3 => b_reg_n_0_18,
   I4 => c_reg_n_0_18,
   I5 => ROTR2_out_27,
   O => T2_19_i_7_n_0
);
T2_19_i_8 : LUT6
  generic map(
   INIT => X"6969699669969696"
  )
 port map (
   I0 => ROTR2_out_6,
   I1 => ROTR2_out_26,
   I2 => ROTR2_out_15,
   I3 => b_reg_n_0_17,
   I4 => c_reg_n_0_17,
   I5 => ROTR2_out_28,
   O => T2_19_i_8_n_0
);
T2_19_i_9 : LUT6
  generic map(
   INIT => X"6969699669969696"
  )
 port map (
   I0 => ROTR2_out_7,
   I1 => ROTR2_out_27,
   I2 => ROTR2_out_16,
   I3 => b_reg_n_0_16,
   I4 => c_reg_n_0_16,
   I5 => ROTR2_out_29,
   O => T2_19_i_9_n_0
);
T2_23_i_2 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => ROTR2_out_9,
   I1 => ROTR2_out_32,
   I2 => ROTR2_out_20,
   O => SIGMA_UCASE_0_23
);
T2_23_i_3 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => ROTR2_out_10,
   I1 => ROTR2_out_1,
   I2 => ROTR2_out_21,
   O => SIGMA_UCASE_0_22
);
T2_23_i_4 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => ROTR2_out_11,
   I1 => ROTR2_out_2,
   I2 => ROTR2_out_22,
   O => SIGMA_UCASE_0_21
);
T2_23_i_5 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => ROTR2_out_12,
   I1 => ROTR2_out_3,
   I2 => ROTR2_out_23,
   O => SIGMA_UCASE_0_20
);
T2_23_i_6 : LUT6
  generic map(
   INIT => X"6969699669969696"
  )
 port map (
   I0 => ROTR2_out_20,
   I1 => ROTR2_out_32,
   I2 => ROTR2_out_9,
   I3 => b_reg_n_0_23,
   I4 => c_reg_n_0_23,
   I5 => ROTR2_out_22,
   O => T2_23_i_6_n_0
);
T2_23_i_7 : LUT6
  generic map(
   INIT => X"6969699669969696"
  )
 port map (
   I0 => ROTR2_out_21,
   I1 => ROTR2_out_1,
   I2 => ROTR2_out_10,
   I3 => b_reg_n_0_22,
   I4 => c_reg_n_0_22,
   I5 => ROTR2_out_23,
   O => T2_23_i_7_n_0
);
T2_23_i_8 : LUT6
  generic map(
   INIT => X"6969699669969696"
  )
 port map (
   I0 => ROTR2_out_22,
   I1 => ROTR2_out_2,
   I2 => ROTR2_out_11,
   I3 => b_reg_n_0_21,
   I4 => c_reg_n_0_21,
   I5 => ROTR2_out_24,
   O => T2_23_i_8_n_0
);
T2_23_i_9 : LUT6
  generic map(
   INIT => X"6969699669969696"
  )
 port map (
   I0 => ROTR2_out_23,
   I1 => ROTR2_out_3,
   I2 => ROTR2_out_12,
   I3 => b_reg_n_0_20,
   I4 => c_reg_n_0_20,
   I5 => ROTR2_out_25,
   O => T2_23_i_9_n_0
);
T2_27_i_2 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => ROTR2_out_5,
   I1 => ROTR2_out_28,
   I2 => ROTR2_out_16,
   O => SIGMA_UCASE_0_27
);
T2_27_i_3 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => ROTR2_out_6,
   I1 => ROTR2_out_29,
   I2 => ROTR2_out_17,
   O => SIGMA_UCASE_0_26
);
T2_27_i_4 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => ROTR2_out_7,
   I1 => ROTR2_out_30,
   I2 => ROTR2_out_18,
   O => SIGMA_UCASE_0_25
);
T2_27_i_5 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => ROTR2_out_8,
   I1 => ROTR2_out_31,
   I2 => ROTR2_out_19,
   O => SIGMA_UCASE_0_24
);
T2_27_i_6 : LUT6
  generic map(
   INIT => X"6969699669969696"
  )
 port map (
   I0 => ROTR2_out_16,
   I1 => ROTR2_out_28,
   I2 => ROTR2_out_5,
   I3 => b_reg_n_0_27,
   I4 => c_reg_n_0_27,
   I5 => ROTR2_out_18,
   O => T2_27_i_6_n_0
);
T2_27_i_7 : LUT6
  generic map(
   INIT => X"6969699669969696"
  )
 port map (
   I0 => ROTR2_out_17,
   I1 => ROTR2_out_29,
   I2 => ROTR2_out_6,
   I3 => b_reg_n_0_26,
   I4 => c_reg_n_0_26,
   I5 => ROTR2_out_19,
   O => T2_27_i_7_n_0
);
T2_27_i_8 : LUT6
  generic map(
   INIT => X"6969699669969696"
  )
 port map (
   I0 => ROTR2_out_18,
   I1 => ROTR2_out_30,
   I2 => ROTR2_out_7,
   I3 => b_reg_n_0_25,
   I4 => c_reg_n_0_25,
   I5 => ROTR2_out_20,
   O => T2_27_i_8_n_0
);
T2_27_i_9 : LUT6
  generic map(
   INIT => X"6969699669969696"
  )
 port map (
   I0 => ROTR2_out_19,
   I1 => ROTR2_out_31,
   I2 => ROTR2_out_8,
   I3 => b_reg_n_0_24,
   I4 => c_reg_n_0_24,
   I5 => ROTR2_out_21,
   O => T2_27_i_9_n_0
);
T2_31_i_2 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => ROTR2_out_2,
   I1 => ROTR2_out_25,
   I2 => ROTR2_out_13,
   O => SIGMA_UCASE_0_30
);
T2_31_i_3 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => ROTR2_out_3,
   I1 => ROTR2_out_26,
   I2 => ROTR2_out_14,
   O => SIGMA_UCASE_0_29
);
T2_31_i_4 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => ROTR2_out_4,
   I1 => ROTR2_out_27,
   I2 => ROTR2_out_15,
   O => SIGMA_UCASE_0_28
);
T2_31_i_5 : LUT6
  generic map(
   INIT => X"6969699669969696"
  )
 port map (
   I0 => ROTR2_out_12,
   I1 => ROTR2_out_24,
   I2 => ROTR2_out_1,
   I3 => b_reg_n_0_31,
   I4 => c_reg_n_0_31,
   I5 => ROTR2_out_14,
   O => T2_31_i_5_n_0
);
T2_31_i_6 : LUT6
  generic map(
   INIT => X"6969699669969696"
  )
 port map (
   I0 => ROTR2_out_13,
   I1 => ROTR2_out_25,
   I2 => ROTR2_out_2,
   I3 => b_reg_n_0_30,
   I4 => c_reg_n_0_30,
   I5 => ROTR2_out_15,
   O => T2_31_i_6_n_0
);
T2_31_i_7 : LUT6
  generic map(
   INIT => X"6969699669969696"
  )
 port map (
   I0 => ROTR2_out_14,
   I1 => ROTR2_out_26,
   I2 => ROTR2_out_3,
   I3 => b_reg_n_0_29,
   I4 => c_reg_n_0_29,
   I5 => ROTR2_out_16,
   O => T2_31_i_7_n_0
);
T2_31_i_8 : LUT6
  generic map(
   INIT => X"6969699669969696"
  )
 port map (
   I0 => ROTR2_out_15,
   I1 => ROTR2_out_27,
   I2 => ROTR2_out_4,
   I3 => b_reg_n_0_28,
   I4 => c_reg_n_0_28,
   I5 => ROTR2_out_17,
   O => T2_31_i_8_n_0
);
T2_3_i_2 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => ROTR2_out_29,
   I1 => ROTR2_out_20,
   I2 => ROTR2_out_8,
   O => SIGMA_UCASE_0_3
);
T2_3_i_3 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => ROTR2_out_30,
   I1 => ROTR2_out_21,
   I2 => ROTR2_out_9,
   O => SIGMA_UCASE_0_2
);
T2_3_i_4 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => ROTR2_out_31,
   I1 => ROTR2_out_22,
   I2 => ROTR2_out_10,
   O => SIGMA_UCASE_0_1
);
T2_3_i_5 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => ROTR2_out_32,
   I1 => ROTR2_out_23,
   I2 => ROTR2_out_11,
   O => SIGMA_UCASE_0_0
);
T2_3_i_6 : LUT6
  generic map(
   INIT => X"6969699669969696"
  )
 port map (
   I0 => ROTR2_out_8,
   I1 => ROTR2_out_20,
   I2 => ROTR2_out_29,
   I3 => b_reg_n_0_3,
   I4 => c_reg_n_0_3,
   I5 => ROTR2_out_10,
   O => T2_3_i_6_n_0
);
T2_3_i_7 : LUT6
  generic map(
   INIT => X"6969699669969696"
  )
 port map (
   I0 => ROTR2_out_9,
   I1 => ROTR2_out_21,
   I2 => ROTR2_out_30,
   I3 => b_reg_n_0_2,
   I4 => c_reg_n_0_2,
   I5 => ROTR2_out_11,
   O => T2_3_i_7_n_0
);
T2_3_i_8 : LUT6
  generic map(
   INIT => X"6969699669969696"
  )
 port map (
   I0 => ROTR2_out_10,
   I1 => ROTR2_out_22,
   I2 => ROTR2_out_31,
   I3 => b_reg_n_0_1,
   I4 => c_reg_n_0_1,
   I5 => ROTR2_out_12,
   O => T2_3_i_8_n_0
);
T2_3_i_9 : LUT6
  generic map(
   INIT => X"6969699669969696"
  )
 port map (
   I0 => ROTR2_out_11,
   I1 => ROTR2_out_23,
   I2 => ROTR2_out_32,
   I3 => b_reg_n_0_0,
   I4 => c_reg_n_0_0,
   I5 => ROTR2_out_13,
   O => T2_3_i_9_n_0
);
T2_7_i_2 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => ROTR2_out_25,
   I1 => ROTR2_out_16,
   I2 => ROTR2_out_4,
   O => SIGMA_UCASE_0_7
);
T2_7_i_3 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => ROTR2_out_26,
   I1 => ROTR2_out_17,
   I2 => ROTR2_out_5,
   O => SIGMA_UCASE_0_6
);
T2_7_i_4 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => ROTR2_out_27,
   I1 => ROTR2_out_18,
   I2 => ROTR2_out_6,
   O => SIGMA_UCASE_0_5
);
T2_7_i_5 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => ROTR2_out_28,
   I1 => ROTR2_out_19,
   I2 => ROTR2_out_7,
   O => SIGMA_UCASE_0_4
);
T2_7_i_6 : LUT6
  generic map(
   INIT => X"6969699669969696"
  )
 port map (
   I0 => ROTR2_out_4,
   I1 => ROTR2_out_16,
   I2 => ROTR2_out_25,
   I3 => b_reg_n_0_7,
   I4 => c_reg_n_0_7,
   I5 => ROTR2_out_6,
   O => T2_7_i_6_n_0
);
T2_7_i_7 : LUT6
  generic map(
   INIT => X"6969699669969696"
  )
 port map (
   I0 => ROTR2_out_5,
   I1 => ROTR2_out_17,
   I2 => ROTR2_out_26,
   I3 => b_reg_n_0_6,
   I4 => c_reg_n_0_6,
   I5 => ROTR2_out_7,
   O => T2_7_i_7_n_0
);
T2_7_i_8 : LUT6
  generic map(
   INIT => X"6969699669969696"
  )
 port map (
   I0 => ROTR2_out_6,
   I1 => ROTR2_out_18,
   I2 => ROTR2_out_27,
   I3 => b_reg_n_0_5,
   I4 => c_reg_n_0_5,
   I5 => ROTR2_out_8,
   O => T2_7_i_8_n_0
);
T2_7_i_9 : LUT6
  generic map(
   INIT => X"6969699669969696"
  )
 port map (
   I0 => ROTR2_out_7,
   I1 => ROTR2_out_19,
   I2 => ROTR2_out_28,
   I3 => b_reg_n_0_4,
   I4 => c_reg_n_0_4,
   I5 => ROTR2_out_9,
   O => T2_7_i_9_n_0
);
T2_reg_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T20_0,
   R => '0',
   Q => T2_0
);
T2_reg_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T20_10,
   R => '0',
   Q => T2_10
);
T2_reg_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T20_11,
   R => '0',
   Q => T2_11
);
T2_reg_11_i_1 : CARRY4
 port map (
   CI => T2_reg_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => SIGMA_UCASE_0_8,
   DI(1) => SIGMA_UCASE_0_9,
   DI(2) => SIGMA_UCASE_0_10,
   DI(3) => SIGMA_UCASE_0_11,
   S(0) => T2_11_i_9_n_0,
   S(1) => T2_11_i_8_n_0,
   S(2) => T2_11_i_7_n_0,
   S(3) => T2_11_i_6_n_0,
   CO(0) => T2_reg_11_i_1_n_3,
   CO(1) => T2_reg_11_i_1_n_2,
   CO(2) => T2_reg_11_i_1_n_1,
   CO(3) => T2_reg_11_i_1_n_0,
   O(0) => T20_8,
   O(1) => T20_9,
   O(2) => T20_10,
   O(3) => T20_11
);
T2_reg_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T20_12,
   R => '0',
   Q => T2_12
);
T2_reg_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T20_13,
   R => '0',
   Q => T2_13
);
T2_reg_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T20_14,
   R => '0',
   Q => T2_14
);
T2_reg_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T20_15,
   R => '0',
   Q => T2_15
);
T2_reg_15_i_1 : CARRY4
 port map (
   CI => T2_reg_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => SIGMA_UCASE_0_12,
   DI(1) => SIGMA_UCASE_0_13,
   DI(2) => SIGMA_UCASE_0_14,
   DI(3) => SIGMA_UCASE_0_15,
   S(0) => T2_15_i_9_n_0,
   S(1) => T2_15_i_8_n_0,
   S(2) => T2_15_i_7_n_0,
   S(3) => T2_15_i_6_n_0,
   CO(0) => T2_reg_15_i_1_n_3,
   CO(1) => T2_reg_15_i_1_n_2,
   CO(2) => T2_reg_15_i_1_n_1,
   CO(3) => T2_reg_15_i_1_n_0,
   O(0) => T20_12,
   O(1) => T20_13,
   O(2) => T20_14,
   O(3) => T20_15
);
T2_reg_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T20_16,
   R => '0',
   Q => T2_16
);
T2_reg_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T20_17,
   R => '0',
   Q => T2_17
);
T2_reg_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T20_18,
   R => '0',
   Q => T2_18
);
T2_reg_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T20_19,
   R => '0',
   Q => T2_19
);
T2_reg_19_i_1 : CARRY4
 port map (
   CI => T2_reg_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => SIGMA_UCASE_0_16,
   DI(1) => SIGMA_UCASE_0_17,
   DI(2) => SIGMA_UCASE_0_18,
   DI(3) => SIGMA_UCASE_0_19,
   S(0) => T2_19_i_9_n_0,
   S(1) => T2_19_i_8_n_0,
   S(2) => T2_19_i_7_n_0,
   S(3) => T2_19_i_6_n_0,
   CO(0) => T2_reg_19_i_1_n_3,
   CO(1) => T2_reg_19_i_1_n_2,
   CO(2) => T2_reg_19_i_1_n_1,
   CO(3) => T2_reg_19_i_1_n_0,
   O(0) => T20_16,
   O(1) => T20_17,
   O(2) => T20_18,
   O(3) => T20_19
);
T2_reg_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T20_1,
   R => '0',
   Q => T2_1
);
T2_reg_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T20_20,
   R => '0',
   Q => T2_20
);
T2_reg_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T20_21,
   R => '0',
   Q => T2_21
);
T2_reg_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T20_22,
   R => '0',
   Q => T2_22
);
T2_reg_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T20_23,
   R => '0',
   Q => T2_23
);
T2_reg_23_i_1 : CARRY4
 port map (
   CI => T2_reg_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => SIGMA_UCASE_0_20,
   DI(1) => SIGMA_UCASE_0_21,
   DI(2) => SIGMA_UCASE_0_22,
   DI(3) => SIGMA_UCASE_0_23,
   S(0) => T2_23_i_9_n_0,
   S(1) => T2_23_i_8_n_0,
   S(2) => T2_23_i_7_n_0,
   S(3) => T2_23_i_6_n_0,
   CO(0) => T2_reg_23_i_1_n_3,
   CO(1) => T2_reg_23_i_1_n_2,
   CO(2) => T2_reg_23_i_1_n_1,
   CO(3) => T2_reg_23_i_1_n_0,
   O(0) => T20_20,
   O(1) => T20_21,
   O(2) => T20_22,
   O(3) => T20_23
);
T2_reg_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T20_24,
   R => '0',
   Q => T2_24
);
T2_reg_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T20_25,
   R => '0',
   Q => T2_25
);
T2_reg_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T20_26,
   R => '0',
   Q => T2_26
);
T2_reg_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T20_27,
   R => '0',
   Q => T2_27
);
T2_reg_27_i_1 : CARRY4
 port map (
   CI => T2_reg_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => SIGMA_UCASE_0_24,
   DI(1) => SIGMA_UCASE_0_25,
   DI(2) => SIGMA_UCASE_0_26,
   DI(3) => SIGMA_UCASE_0_27,
   S(0) => T2_27_i_9_n_0,
   S(1) => T2_27_i_8_n_0,
   S(2) => T2_27_i_7_n_0,
   S(3) => T2_27_i_6_n_0,
   CO(0) => T2_reg_27_i_1_n_3,
   CO(1) => T2_reg_27_i_1_n_2,
   CO(2) => T2_reg_27_i_1_n_1,
   CO(3) => T2_reg_27_i_1_n_0,
   O(0) => T20_24,
   O(1) => T20_25,
   O(2) => T20_26,
   O(3) => T20_27
);
T2_reg_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T20_28,
   R => '0',
   Q => T2_28
);
T2_reg_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T20_29,
   R => '0',
   Q => T2_29
);
T2_reg_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T20_2,
   R => '0',
   Q => T2_2
);
T2_reg_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T20_30,
   R => '0',
   Q => T2_30
);
T2_reg_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T20_31,
   R => '0',
   Q => T2_31
);
T2_reg_31_i_1 : CARRY4
 port map (
   CI => T2_reg_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => SIGMA_UCASE_0_28,
   DI(1) => SIGMA_UCASE_0_29,
   DI(2) => SIGMA_UCASE_0_30,
   DI(3) => '0',
   S(0) => T2_31_i_8_n_0,
   S(1) => T2_31_i_7_n_0,
   S(2) => T2_31_i_6_n_0,
   S(3) => T2_31_i_5_n_0,
   CO(0) => T2_reg_31_i_1_n_3,
   CO(1) => T2_reg_31_i_1_n_2,
   CO(2) => T2_reg_31_i_1_n_1,
   CO(3) => NLW_T2_reg_31_i_1_CO_UNCONNECTED_3,
   O(0) => T20_28,
   O(1) => T20_29,
   O(2) => T20_30,
   O(3) => T20_31
);
T2_reg_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T20_3,
   R => '0',
   Q => T2_3
);
T2_reg_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => SIGMA_UCASE_0_0,
   DI(1) => SIGMA_UCASE_0_1,
   DI(2) => SIGMA_UCASE_0_2,
   DI(3) => SIGMA_UCASE_0_3,
   S(0) => T2_3_i_9_n_0,
   S(1) => T2_3_i_8_n_0,
   S(2) => T2_3_i_7_n_0,
   S(3) => T2_3_i_6_n_0,
   CO(0) => T2_reg_3_i_1_n_3,
   CO(1) => T2_reg_3_i_1_n_2,
   CO(2) => T2_reg_3_i_1_n_1,
   CO(3) => T2_reg_3_i_1_n_0,
   O(0) => T20_0,
   O(1) => T20_1,
   O(2) => T20_2,
   O(3) => T20_3
);
T2_reg_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T20_4,
   R => '0',
   Q => T2_4
);
T2_reg_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T20_5,
   R => '0',
   Q => T2_5
);
T2_reg_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T20_6,
   R => '0',
   Q => T2_6
);
T2_reg_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T20_7,
   R => '0',
   Q => T2_7
);
T2_reg_7_i_1 : CARRY4
 port map (
   CI => T2_reg_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => SIGMA_UCASE_0_4,
   DI(1) => SIGMA_UCASE_0_5,
   DI(2) => SIGMA_UCASE_0_6,
   DI(3) => SIGMA_UCASE_0_7,
   S(0) => T2_7_i_9_n_0,
   S(1) => T2_7_i_8_n_0,
   S(2) => T2_7_i_7_n_0,
   S(3) => T2_7_i_6_n_0,
   CO(0) => T2_reg_7_i_1_n_3,
   CO(1) => T2_reg_7_i_1_n_2,
   CO(2) => T2_reg_7_i_1_n_1,
   CO(3) => T2_reg_7_i_1_n_0,
   O(0) => T20_4,
   O(1) => T20_5,
   O(2) => T20_6,
   O(3) => T20_7
);
T2_reg_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T20_8,
   R => '0',
   Q => T2_8
);
T2_reg_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => T1_31_i_1_n_0,
   D => T20_9,
   R => '0',
   Q => T2_9
);
W_0_31_i_1 : LUT2
  generic map(
   INIT => X"2"
  )
 port map (
   I0 => W_0,
   I1 => rst_IBUF,
   O => W_reg_0_0
);
W_16_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_0_10,
   I1 => M_reg_9_10,
   I2 => M_reg_1_28,
   I3 => M_reg_1_17,
   I4 => M_reg_1_13,
   O => W_16_11_i_10_n_0
);
W_16_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_9_9,
   I1 => M_reg_1_12,
   I2 => M_reg_1_16,
   I3 => M_reg_1_27,
   I4 => M_reg_0_9,
   O => W_16_11_i_11_n_0
);
W_16_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_0_9,
   I1 => M_reg_9_9,
   I2 => M_reg_1_27,
   I3 => M_reg_1_16,
   I4 => M_reg_1_12,
   O => W_16_11_i_12_n_0
);
W_16_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_9_8,
   I1 => M_reg_1_11,
   I2 => M_reg_1_15,
   I3 => M_reg_1_26,
   I4 => M_reg_0_8,
   O => W_16_11_i_13_n_0
);
W_16_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_0_8,
   I1 => M_reg_9_8,
   I2 => M_reg_1_26,
   I3 => M_reg_1_15,
   I4 => M_reg_1_11,
   O => W_16_11_i_14_n_0
);
W_16_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_9_7,
   I1 => M_reg_1_10,
   I2 => M_reg_1_14,
   I3 => M_reg_1_25,
   I4 => M_reg_0_7,
   O => W_16_11_i_15_n_0
);
W_16_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_0_7,
   I1 => M_reg_9_7,
   I2 => M_reg_1_25,
   I3 => M_reg_1_14,
   I4 => M_reg_1_10,
   O => W_16_11_i_16_n_0
);
W_16_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_9_6,
   I1 => M_reg_1_9,
   I2 => M_reg_1_13,
   I3 => M_reg_1_24,
   I4 => M_reg_0_6,
   O => W_16_11_i_17_n_0
);
W_16_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => M_reg_14_20,
   I1 => M_reg_14_27,
   I2 => M_reg_14_29,
   I3 => W_16_11_i_10_n_0,
   I4 => W_16_11_i_11_n_0,
   O => W_16_11_i_2_n_0
);
W_16_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => M_reg_14_19,
   I1 => M_reg_14_26,
   I2 => M_reg_14_28,
   I3 => W_16_11_i_12_n_0,
   I4 => W_16_11_i_13_n_0,
   O => W_16_11_i_3_n_0
);
W_16_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => M_reg_14_18,
   I1 => M_reg_14_25,
   I2 => M_reg_14_27,
   I3 => W_16_11_i_14_n_0,
   I4 => W_16_11_i_15_n_0,
   O => W_16_11_i_4_n_0
);
W_16_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => M_reg_14_17,
   I1 => M_reg_14_24,
   I2 => M_reg_14_26,
   I3 => W_16_11_i_16_n_0,
   I4 => W_16_11_i_17_n_0,
   O => W_16_11_i_5_n_0
);
W_16_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_16_11_i_2_n_0,
   I1 => W_16_15_i_16_n_0,
   I2 => M_reg_14_21,
   I3 => M_reg_14_28,
   I4 => M_reg_14_30,
   I5 => W_16_15_i_17_n_0,
   O => W_16_11_i_6_n_0
);
W_16_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_16_11_i_3_n_0,
   I1 => W_16_11_i_10_n_0,
   I2 => M_reg_14_20,
   I3 => M_reg_14_27,
   I4 => M_reg_14_29,
   I5 => W_16_11_i_11_n_0,
   O => W_16_11_i_7_n_0
);
W_16_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_16_11_i_4_n_0,
   I1 => W_16_11_i_12_n_0,
   I2 => M_reg_14_19,
   I3 => M_reg_14_26,
   I4 => M_reg_14_28,
   I5 => W_16_11_i_13_n_0,
   O => W_16_11_i_8_n_0
);
W_16_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_16_11_i_5_n_0,
   I1 => W_16_11_i_14_n_0,
   I2 => M_reg_14_18,
   I3 => M_reg_14_25,
   I4 => M_reg_14_27,
   I5 => W_16_11_i_15_n_0,
   O => W_16_11_i_9_n_0
);
W_16_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_0_14,
   I1 => M_reg_9_14,
   I2 => M_reg_1_0,
   I3 => M_reg_1_21,
   I4 => M_reg_1_17,
   O => W_16_15_i_10_n_0
);
W_16_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_9_13,
   I1 => M_reg_1_16,
   I2 => M_reg_1_20,
   I3 => M_reg_1_31,
   I4 => M_reg_0_13,
   O => W_16_15_i_11_n_0
);
W_16_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_0_13,
   I1 => M_reg_9_13,
   I2 => M_reg_1_31,
   I3 => M_reg_1_20,
   I4 => M_reg_1_16,
   O => W_16_15_i_12_n_0
);
W_16_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_9_12,
   I1 => M_reg_1_15,
   I2 => M_reg_1_19,
   I3 => M_reg_1_30,
   I4 => M_reg_0_12,
   O => W_16_15_i_13_n_0
);
W_16_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_0_12,
   I1 => M_reg_9_12,
   I2 => M_reg_1_30,
   I3 => M_reg_1_19,
   I4 => M_reg_1_15,
   O => W_16_15_i_14_n_0
);
W_16_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_9_11,
   I1 => M_reg_1_14,
   I2 => M_reg_1_18,
   I3 => M_reg_1_29,
   I4 => M_reg_0_11,
   O => W_16_15_i_15_n_0
);
W_16_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_0_11,
   I1 => M_reg_9_11,
   I2 => M_reg_1_29,
   I3 => M_reg_1_18,
   I4 => M_reg_1_14,
   O => W_16_15_i_16_n_0
);
W_16_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_9_10,
   I1 => M_reg_1_13,
   I2 => M_reg_1_17,
   I3 => M_reg_1_28,
   I4 => M_reg_0_10,
   O => W_16_15_i_17_n_0
);
W_16_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => M_reg_14_24,
   I1 => M_reg_14_31,
   I2 => M_reg_14_1,
   I3 => W_16_15_i_10_n_0,
   I4 => W_16_15_i_11_n_0,
   O => W_16_15_i_2_n_0
);
W_16_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => M_reg_14_23,
   I1 => M_reg_14_30,
   I2 => M_reg_14_0,
   I3 => W_16_15_i_12_n_0,
   I4 => W_16_15_i_13_n_0,
   O => W_16_15_i_3_n_0
);
W_16_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => M_reg_14_22,
   I1 => M_reg_14_29,
   I2 => M_reg_14_31,
   I3 => W_16_15_i_14_n_0,
   I4 => W_16_15_i_15_n_0,
   O => W_16_15_i_4_n_0
);
W_16_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => M_reg_14_21,
   I1 => M_reg_14_28,
   I2 => M_reg_14_30,
   I3 => W_16_15_i_16_n_0,
   I4 => W_16_15_i_17_n_0,
   O => W_16_15_i_5_n_0
);
W_16_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_16_15_i_2_n_0,
   I1 => W_16_19_i_16_n_0,
   I2 => M_reg_14_25,
   I3 => M_reg_14_0,
   I4 => M_reg_14_2,
   I5 => W_16_19_i_17_n_0,
   O => W_16_15_i_6_n_0
);
W_16_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_16_15_i_3_n_0,
   I1 => W_16_15_i_10_n_0,
   I2 => M_reg_14_24,
   I3 => M_reg_14_31,
   I4 => M_reg_14_1,
   I5 => W_16_15_i_11_n_0,
   O => W_16_15_i_7_n_0
);
W_16_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_16_15_i_4_n_0,
   I1 => W_16_15_i_12_n_0,
   I2 => M_reg_14_23,
   I3 => M_reg_14_30,
   I4 => M_reg_14_0,
   I5 => W_16_15_i_13_n_0,
   O => W_16_15_i_8_n_0
);
W_16_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_16_15_i_5_n_0,
   I1 => W_16_15_i_14_n_0,
   I2 => M_reg_14_22,
   I3 => M_reg_14_29,
   I4 => M_reg_14_31,
   I5 => W_16_15_i_15_n_0,
   O => W_16_15_i_9_n_0
);
W_16_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_0_18,
   I1 => M_reg_9_18,
   I2 => M_reg_1_4,
   I3 => M_reg_1_25,
   I4 => M_reg_1_21,
   O => W_16_19_i_10_n_0
);
W_16_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_9_17,
   I1 => M_reg_1_20,
   I2 => M_reg_1_24,
   I3 => M_reg_1_3,
   I4 => M_reg_0_17,
   O => W_16_19_i_11_n_0
);
W_16_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_0_17,
   I1 => M_reg_9_17,
   I2 => M_reg_1_3,
   I3 => M_reg_1_24,
   I4 => M_reg_1_20,
   O => W_16_19_i_12_n_0
);
W_16_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_9_16,
   I1 => M_reg_1_19,
   I2 => M_reg_1_23,
   I3 => M_reg_1_2,
   I4 => M_reg_0_16,
   O => W_16_19_i_13_n_0
);
W_16_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_0_16,
   I1 => M_reg_9_16,
   I2 => M_reg_1_2,
   I3 => M_reg_1_23,
   I4 => M_reg_1_19,
   O => W_16_19_i_14_n_0
);
W_16_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_9_15,
   I1 => M_reg_1_18,
   I2 => M_reg_1_22,
   I3 => M_reg_1_1,
   I4 => M_reg_0_15,
   O => W_16_19_i_15_n_0
);
W_16_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_0_15,
   I1 => M_reg_9_15,
   I2 => M_reg_1_1,
   I3 => M_reg_1_22,
   I4 => M_reg_1_18,
   O => W_16_19_i_16_n_0
);
W_16_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_9_14,
   I1 => M_reg_1_17,
   I2 => M_reg_1_21,
   I3 => M_reg_1_0,
   I4 => M_reg_0_14,
   O => W_16_19_i_17_n_0
);
W_16_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => M_reg_14_28,
   I1 => M_reg_14_3,
   I2 => M_reg_14_5,
   I3 => W_16_19_i_10_n_0,
   I4 => W_16_19_i_11_n_0,
   O => W_16_19_i_2_n_0
);
W_16_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => M_reg_14_27,
   I1 => M_reg_14_2,
   I2 => M_reg_14_4,
   I3 => W_16_19_i_12_n_0,
   I4 => W_16_19_i_13_n_0,
   O => W_16_19_i_3_n_0
);
W_16_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => M_reg_14_26,
   I1 => M_reg_14_1,
   I2 => M_reg_14_3,
   I3 => W_16_19_i_14_n_0,
   I4 => W_16_19_i_15_n_0,
   O => W_16_19_i_4_n_0
);
W_16_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => M_reg_14_25,
   I1 => M_reg_14_0,
   I2 => M_reg_14_2,
   I3 => W_16_19_i_16_n_0,
   I4 => W_16_19_i_17_n_0,
   O => W_16_19_i_5_n_0
);
W_16_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_16_19_i_2_n_0,
   I1 => W_16_23_i_16_n_0,
   I2 => M_reg_14_29,
   I3 => M_reg_14_4,
   I4 => M_reg_14_6,
   I5 => W_16_23_i_17_n_0,
   O => W_16_19_i_6_n_0
);
W_16_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_16_19_i_3_n_0,
   I1 => W_16_19_i_10_n_0,
   I2 => M_reg_14_28,
   I3 => M_reg_14_3,
   I4 => M_reg_14_5,
   I5 => W_16_19_i_11_n_0,
   O => W_16_19_i_7_n_0
);
W_16_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_16_19_i_4_n_0,
   I1 => W_16_19_i_12_n_0,
   I2 => M_reg_14_27,
   I3 => M_reg_14_2,
   I4 => M_reg_14_4,
   I5 => W_16_19_i_13_n_0,
   O => W_16_19_i_8_n_0
);
W_16_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_16_19_i_5_n_0,
   I1 => W_16_19_i_14_n_0,
   I2 => M_reg_14_26,
   I3 => M_reg_14_1,
   I4 => M_reg_14_3,
   I5 => W_16_19_i_15_n_0,
   O => W_16_19_i_9_n_0
);
W_16_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_0_22,
   I1 => M_reg_9_22,
   I2 => M_reg_1_8,
   I3 => M_reg_1_29,
   I4 => M_reg_1_25,
   O => W_16_23_i_10_n_0
);
W_16_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_9_21,
   I1 => M_reg_1_24,
   I2 => M_reg_1_28,
   I3 => M_reg_1_7,
   I4 => M_reg_0_21,
   O => W_16_23_i_11_n_0
);
W_16_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_0_21,
   I1 => M_reg_9_21,
   I2 => M_reg_1_7,
   I3 => M_reg_1_28,
   I4 => M_reg_1_24,
   O => W_16_23_i_12_n_0
);
W_16_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_9_20,
   I1 => M_reg_1_23,
   I2 => M_reg_1_27,
   I3 => M_reg_1_6,
   I4 => M_reg_0_20,
   O => W_16_23_i_13_n_0
);
W_16_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_0_20,
   I1 => M_reg_9_20,
   I2 => M_reg_1_6,
   I3 => M_reg_1_27,
   I4 => M_reg_1_23,
   O => W_16_23_i_14_n_0
);
W_16_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_9_19,
   I1 => M_reg_1_22,
   I2 => M_reg_1_26,
   I3 => M_reg_1_5,
   I4 => M_reg_0_19,
   O => W_16_23_i_15_n_0
);
W_16_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_0_19,
   I1 => M_reg_9_19,
   I2 => M_reg_1_5,
   I3 => M_reg_1_26,
   I4 => M_reg_1_22,
   O => W_16_23_i_16_n_0
);
W_16_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_9_18,
   I1 => M_reg_1_21,
   I2 => M_reg_1_25,
   I3 => M_reg_1_4,
   I4 => M_reg_0_18,
   O => W_16_23_i_17_n_0
);
W_16_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => M_reg_14_7,
   I1 => M_reg_14_9,
   I2 => W_16_23_i_10_n_0,
   I3 => W_16_23_i_11_n_0,
   O => W_16_23_i_2_n_0
);
W_16_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => M_reg_14_31,
   I1 => M_reg_14_6,
   I2 => M_reg_14_8,
   I3 => W_16_23_i_12_n_0,
   I4 => W_16_23_i_13_n_0,
   O => W_16_23_i_3_n_0
);
W_16_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => M_reg_14_30,
   I1 => M_reg_14_5,
   I2 => M_reg_14_7,
   I3 => W_16_23_i_14_n_0,
   I4 => W_16_23_i_15_n_0,
   O => W_16_23_i_4_n_0
);
W_16_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => M_reg_14_29,
   I1 => M_reg_14_4,
   I2 => M_reg_14_6,
   I3 => W_16_23_i_16_n_0,
   I4 => W_16_23_i_17_n_0,
   O => W_16_23_i_5_n_0
);
W_16_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_14_8,
   I1 => M_reg_14_10,
   I2 => W_16_27_i_16_n_0,
   I3 => W_16_27_i_17_n_0,
   I4 => W_16_23_i_2_n_0,
   O => W_16_23_i_6_n_0
);
W_16_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_14_7,
   I1 => M_reg_14_9,
   I2 => W_16_23_i_10_n_0,
   I3 => W_16_23_i_11_n_0,
   I4 => W_16_23_i_3_n_0,
   O => W_16_23_i_7_n_0
);
W_16_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_16_23_i_4_n_0,
   I1 => W_16_23_i_12_n_0,
   I2 => M_reg_14_31,
   I3 => M_reg_14_6,
   I4 => M_reg_14_8,
   I5 => W_16_23_i_13_n_0,
   O => W_16_23_i_8_n_0
);
W_16_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_16_23_i_5_n_0,
   I1 => W_16_23_i_14_n_0,
   I2 => M_reg_14_30,
   I3 => M_reg_14_5,
   I4 => M_reg_14_7,
   I5 => W_16_23_i_15_n_0,
   O => W_16_23_i_9_n_0
);
W_16_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_0_26,
   I1 => M_reg_9_26,
   I2 => M_reg_1_12,
   I3 => M_reg_1_1,
   I4 => M_reg_1_29,
   O => W_16_27_i_10_n_0
);
W_16_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_9_25,
   I1 => M_reg_1_28,
   I2 => M_reg_1_0,
   I3 => M_reg_1_11,
   I4 => M_reg_0_25,
   O => W_16_27_i_11_n_0
);
W_16_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_0_25,
   I1 => M_reg_9_25,
   I2 => M_reg_1_11,
   I3 => M_reg_1_0,
   I4 => M_reg_1_28,
   O => W_16_27_i_12_n_0
);
W_16_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_9_24,
   I1 => M_reg_1_27,
   I2 => M_reg_1_31,
   I3 => M_reg_1_10,
   I4 => M_reg_0_24,
   O => W_16_27_i_13_n_0
);
W_16_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_0_24,
   I1 => M_reg_9_24,
   I2 => M_reg_1_10,
   I3 => M_reg_1_31,
   I4 => M_reg_1_27,
   O => W_16_27_i_14_n_0
);
W_16_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_9_23,
   I1 => M_reg_1_26,
   I2 => M_reg_1_30,
   I3 => M_reg_1_9,
   I4 => M_reg_0_23,
   O => W_16_27_i_15_n_0
);
W_16_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_0_23,
   I1 => M_reg_9_23,
   I2 => M_reg_1_9,
   I3 => M_reg_1_30,
   I4 => M_reg_1_26,
   O => W_16_27_i_16_n_0
);
W_16_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_9_22,
   I1 => M_reg_1_25,
   I2 => M_reg_1_29,
   I3 => M_reg_1_8,
   I4 => M_reg_0_22,
   O => W_16_27_i_17_n_0
);
W_16_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => M_reg_14_11,
   I1 => M_reg_14_13,
   I2 => W_16_27_i_10_n_0,
   I3 => W_16_27_i_11_n_0,
   O => W_16_27_i_2_n_0
);
W_16_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => M_reg_14_10,
   I1 => M_reg_14_12,
   I2 => W_16_27_i_12_n_0,
   I3 => W_16_27_i_13_n_0,
   O => W_16_27_i_3_n_0
);
W_16_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => M_reg_14_9,
   I1 => M_reg_14_11,
   I2 => W_16_27_i_14_n_0,
   I3 => W_16_27_i_15_n_0,
   O => W_16_27_i_4_n_0
);
W_16_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => M_reg_14_8,
   I1 => M_reg_14_10,
   I2 => W_16_27_i_16_n_0,
   I3 => W_16_27_i_17_n_0,
   O => W_16_27_i_5_n_0
);
W_16_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_14_12,
   I1 => M_reg_14_14,
   I2 => W_16_31_i_14_n_0,
   I3 => W_16_31_i_15_n_0,
   I4 => W_16_27_i_2_n_0,
   O => W_16_27_i_6_n_0
);
W_16_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_14_11,
   I1 => M_reg_14_13,
   I2 => W_16_27_i_10_n_0,
   I3 => W_16_27_i_11_n_0,
   I4 => W_16_27_i_3_n_0,
   O => W_16_27_i_7_n_0
);
W_16_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_14_10,
   I1 => M_reg_14_12,
   I2 => W_16_27_i_12_n_0,
   I3 => W_16_27_i_13_n_0,
   I4 => W_16_27_i_4_n_0,
   O => W_16_27_i_8_n_0
);
W_16_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_14_9,
   I1 => M_reg_14_11,
   I2 => W_16_27_i_14_n_0,
   I3 => W_16_27_i_15_n_0,
   I4 => W_16_27_i_5_n_0,
   O => W_16_27_i_9_n_0
);
W_16_31_i_1 : LUT2
  generic map(
   INIT => X"2"
  )
 port map (
   I0 => W_16,
   I1 => rst_IBUF,
   O => W_reg_16_0
);
W_16_31_i_10 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => M_reg_0_29,
   I1 => M_reg_9_29,
   I2 => M_reg_1_15,
   I3 => M_reg_1_4,
   O => W_16_31_i_10_n_0
);
W_16_31_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_9_28,
   I1 => M_reg_1_31,
   I2 => M_reg_1_3,
   I3 => M_reg_1_14,
   I4 => M_reg_0_28,
   O => W_16_31_i_11_n_0
);
W_16_31_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_0_28,
   I1 => M_reg_9_28,
   I2 => M_reg_1_14,
   I3 => M_reg_1_3,
   I4 => M_reg_1_31,
   O => W_16_31_i_12_n_0
);
W_16_31_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_9_27,
   I1 => M_reg_1_30,
   I2 => M_reg_1_2,
   I3 => M_reg_1_13,
   I4 => M_reg_0_27,
   O => W_16_31_i_13_n_0
);
W_16_31_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_0_27,
   I1 => M_reg_9_27,
   I2 => M_reg_1_13,
   I3 => M_reg_1_2,
   I4 => M_reg_1_30,
   O => W_16_31_i_14_n_0
);
W_16_31_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_9_26,
   I1 => M_reg_1_29,
   I2 => M_reg_1_1,
   I3 => M_reg_1_12,
   I4 => M_reg_0_26,
   O => W_16_31_i_15_n_0
);
W_16_31_i_16 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => M_reg_9_29,
   I1 => M_reg_1_4,
   I2 => M_reg_1_15,
   I3 => M_reg_0_29,
   O => W_16_31_i_16_n_0
);
W_16_31_i_17 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => M_reg_14_17,
   I1 => M_reg_14_15,
   O => SIGMA_LCASE_1387_out_30
);
W_16_31_i_18 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => M_reg_1_6,
   I1 => M_reg_1_17,
   I2 => M_reg_9_31,
   I3 => M_reg_0_31,
   I4 => M_reg_14_16,
   I5 => M_reg_14_18,
   O => W_16_31_i_18_n_0
);
W_16_31_i_19 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => M_reg_1_16,
   I1 => M_reg_1_5,
   O => SIGMA_LCASE_0383_out_30
);
W_16_31_i_20 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => M_reg_0_30,
   I1 => M_reg_9_30,
   I2 => M_reg_1_16,
   I3 => M_reg_1_5,
   O => W_16_31_i_20_n_0
);
W_16_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => M_reg_14_14,
   I1 => M_reg_14_16,
   I2 => W_16_31_i_10_n_0,
   I3 => W_16_31_i_11_n_0,
   O => W_16_31_i_3_n_0
);
W_16_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => M_reg_14_13,
   I1 => M_reg_14_15,
   I2 => W_16_31_i_12_n_0,
   I3 => W_16_31_i_13_n_0,
   O => W_16_31_i_4_n_0
);
W_16_31_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => M_reg_14_12,
   I1 => M_reg_14_14,
   I2 => W_16_31_i_14_n_0,
   I3 => W_16_31_i_15_n_0,
   O => W_16_31_i_5_n_0
);
W_16_31_i_6 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_16_31_i_16_n_0,
   I1 => SIGMA_LCASE_1387_out_30,
   I2 => W_16_31_i_18_n_0,
   I3 => M_reg_9_30,
   I4 => SIGMA_LCASE_0383_out_30,
   I5 => M_reg_0_30,
   O => W_16_31_i_6_n_0
);
W_16_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_16_31_i_3_n_0,
   I1 => W_16_31_i_20_n_0,
   I2 => M_reg_14_15,
   I3 => M_reg_14_17,
   I4 => W_16_31_i_16_n_0,
   O => W_16_31_i_7_n_0
);
W_16_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_14_14,
   I1 => M_reg_14_16,
   I2 => W_16_31_i_10_n_0,
   I3 => W_16_31_i_11_n_0,
   I4 => W_16_31_i_4_n_0,
   O => W_16_31_i_8_n_0
);
W_16_31_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_14_13,
   I1 => M_reg_14_15,
   I2 => W_16_31_i_12_n_0,
   I3 => W_16_31_i_13_n_0,
   I4 => W_16_31_i_5_n_0,
   O => W_16_31_i_9_n_0
);
W_16_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_0_2,
   I1 => M_reg_9_2,
   I2 => M_reg_1_20,
   I3 => M_reg_1_9,
   I4 => M_reg_1_5,
   O => W_16_3_i_10_n_0
);
W_16_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_9_1,
   I1 => M_reg_1_4,
   I2 => M_reg_1_8,
   I3 => M_reg_1_19,
   I4 => M_reg_0_1,
   O => W_16_3_i_11_n_0
);
W_16_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => M_reg_1_19,
   I1 => M_reg_1_8,
   I2 => M_reg_1_4,
   O => SIGMA_LCASE_0383_out_1
);
W_16_3_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_0_1,
   I1 => M_reg_9_1,
   I2 => M_reg_1_19,
   I3 => M_reg_1_8,
   I4 => M_reg_1_4,
   O => W_16_3_i_13_n_0
);
W_16_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => M_reg_14_12,
   I1 => M_reg_14_19,
   I2 => M_reg_14_21,
   I3 => W_16_3_i_10_n_0,
   I4 => W_16_3_i_11_n_0,
   O => W_16_3_i_2_n_0
);
W_16_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_16_3_i_11_n_0,
   I1 => M_reg_14_21,
   I2 => M_reg_14_19,
   I3 => M_reg_14_12,
   I4 => W_16_3_i_10_n_0,
   O => W_16_3_i_3_n_0
);
W_16_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_0383_out_1,
   I1 => M_reg_9_1,
   I2 => M_reg_0_1,
   I3 => M_reg_14_11,
   I4 => M_reg_14_18,
   I5 => M_reg_14_20,
   O => W_16_3_i_4_n_0
);
W_16_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_0_0,
   I1 => M_reg_9_0,
   I2 => M_reg_1_18,
   I3 => M_reg_1_7,
   I4 => M_reg_1_3,
   O => W_16_3_i_5_n_0
);
W_16_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_16_3_i_2_n_0,
   I1 => W_16_7_i_16_n_0,
   I2 => M_reg_14_13,
   I3 => M_reg_14_20,
   I4 => M_reg_14_22,
   I5 => W_16_7_i_17_n_0,
   O => W_16_3_i_6_n_0
);
W_16_3_i_7 : LUT5
  generic map(
   INIT => X"6aa6a66a"
  )
 port map (
   I0 => W_16_3_i_3_n_0,
   I1 => W_16_3_i_13_n_0,
   I2 => M_reg_14_20,
   I3 => M_reg_14_18,
   I4 => M_reg_14_11,
   O => W_16_3_i_7_n_0
);
W_16_3_i_8 : LUT6
  generic map(
   INIT => X"566565566aa6a66a"
  )
 port map (
   I0 => W_16_3_i_4_n_0,
   I1 => M_reg_0_0,
   I2 => M_reg_1_18,
   I3 => M_reg_1_7,
   I4 => M_reg_1_3,
   I5 => M_reg_9_0,
   O => W_16_3_i_8_n_0
);
W_16_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_16_3_i_5_n_0,
   I1 => M_reg_14_10,
   I2 => M_reg_14_17,
   I3 => M_reg_14_19,
   O => W_16_3_i_9_n_0
);
W_16_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_0_6,
   I1 => M_reg_9_6,
   I2 => M_reg_1_24,
   I3 => M_reg_1_13,
   I4 => M_reg_1_9,
   O => W_16_7_i_10_n_0
);
W_16_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_9_5,
   I1 => M_reg_1_8,
   I2 => M_reg_1_12,
   I3 => M_reg_1_23,
   I4 => M_reg_0_5,
   O => W_16_7_i_11_n_0
);
W_16_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_0_5,
   I1 => M_reg_9_5,
   I2 => M_reg_1_23,
   I3 => M_reg_1_12,
   I4 => M_reg_1_8,
   O => W_16_7_i_12_n_0
);
W_16_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_9_4,
   I1 => M_reg_1_7,
   I2 => M_reg_1_11,
   I3 => M_reg_1_22,
   I4 => M_reg_0_4,
   O => W_16_7_i_13_n_0
);
W_16_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_0_4,
   I1 => M_reg_9_4,
   I2 => M_reg_1_22,
   I3 => M_reg_1_11,
   I4 => M_reg_1_7,
   O => W_16_7_i_14_n_0
);
W_16_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_9_3,
   I1 => M_reg_1_6,
   I2 => M_reg_1_10,
   I3 => M_reg_1_21,
   I4 => M_reg_0_3,
   O => W_16_7_i_15_n_0
);
W_16_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_0_3,
   I1 => M_reg_9_3,
   I2 => M_reg_1_21,
   I3 => M_reg_1_10,
   I4 => M_reg_1_6,
   O => W_16_7_i_16_n_0
);
W_16_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_9_2,
   I1 => M_reg_1_5,
   I2 => M_reg_1_9,
   I3 => M_reg_1_20,
   I4 => M_reg_0_2,
   O => W_16_7_i_17_n_0
);
W_16_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => M_reg_14_16,
   I1 => M_reg_14_23,
   I2 => M_reg_14_25,
   I3 => W_16_7_i_10_n_0,
   I4 => W_16_7_i_11_n_0,
   O => W_16_7_i_2_n_0
);
W_16_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => M_reg_14_15,
   I1 => M_reg_14_22,
   I2 => M_reg_14_24,
   I3 => W_16_7_i_12_n_0,
   I4 => W_16_7_i_13_n_0,
   O => W_16_7_i_3_n_0
);
W_16_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => M_reg_14_14,
   I1 => M_reg_14_21,
   I2 => M_reg_14_23,
   I3 => W_16_7_i_14_n_0,
   I4 => W_16_7_i_15_n_0,
   O => W_16_7_i_4_n_0
);
W_16_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => M_reg_14_13,
   I1 => M_reg_14_20,
   I2 => M_reg_14_22,
   I3 => W_16_7_i_16_n_0,
   I4 => W_16_7_i_17_n_0,
   O => W_16_7_i_5_n_0
);
W_16_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_16_7_i_2_n_0,
   I1 => W_16_11_i_16_n_0,
   I2 => M_reg_14_17,
   I3 => M_reg_14_24,
   I4 => M_reg_14_26,
   I5 => W_16_11_i_17_n_0,
   O => W_16_7_i_6_n_0
);
W_16_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_16_7_i_3_n_0,
   I1 => W_16_7_i_10_n_0,
   I2 => M_reg_14_16,
   I3 => M_reg_14_23,
   I4 => M_reg_14_25,
   I5 => W_16_7_i_11_n_0,
   O => W_16_7_i_7_n_0
);
W_16_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_16_7_i_4_n_0,
   I1 => W_16_7_i_12_n_0,
   I2 => M_reg_14_15,
   I3 => M_reg_14_22,
   I4 => M_reg_14_24,
   I5 => W_16_7_i_13_n_0,
   O => W_16_7_i_8_n_0
);
W_16_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_16_7_i_5_n_0,
   I1 => W_16_7_i_14_n_0,
   I2 => M_reg_14_14,
   I3 => M_reg_14_21,
   I4 => M_reg_14_23,
   I5 => W_16_7_i_15_n_0,
   O => W_16_7_i_9_n_0
);
W_17_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_1_10,
   I1 => M_reg_10_10,
   I2 => M_reg_2_28,
   I3 => M_reg_2_17,
   I4 => M_reg_2_13,
   O => W_17_11_i_10_n_0
);
W_17_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_10_9,
   I1 => M_reg_2_12,
   I2 => M_reg_2_16,
   I3 => M_reg_2_27,
   I4 => M_reg_1_9,
   O => W_17_11_i_11_n_0
);
W_17_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_1_9,
   I1 => M_reg_10_9,
   I2 => M_reg_2_27,
   I3 => M_reg_2_16,
   I4 => M_reg_2_12,
   O => W_17_11_i_12_n_0
);
W_17_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_10_8,
   I1 => M_reg_2_11,
   I2 => M_reg_2_15,
   I3 => M_reg_2_26,
   I4 => M_reg_1_8,
   O => W_17_11_i_13_n_0
);
W_17_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_1_8,
   I1 => M_reg_10_8,
   I2 => M_reg_2_26,
   I3 => M_reg_2_15,
   I4 => M_reg_2_11,
   O => W_17_11_i_14_n_0
);
W_17_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_10_7,
   I1 => M_reg_2_10,
   I2 => M_reg_2_14,
   I3 => M_reg_2_25,
   I4 => M_reg_1_7,
   O => W_17_11_i_15_n_0
);
W_17_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_1_7,
   I1 => M_reg_10_7,
   I2 => M_reg_2_25,
   I3 => M_reg_2_14,
   I4 => M_reg_2_10,
   O => W_17_11_i_16_n_0
);
W_17_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_10_6,
   I1 => M_reg_2_9,
   I2 => M_reg_2_13,
   I3 => M_reg_2_24,
   I4 => M_reg_1_6,
   O => W_17_11_i_17_n_0
);
W_17_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => M_reg_15_20,
   I1 => M_reg_15_27,
   I2 => M_reg_15_29,
   I3 => W_17_11_i_10_n_0,
   I4 => W_17_11_i_11_n_0,
   O => W_17_11_i_2_n_0
);
W_17_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => M_reg_15_19,
   I1 => M_reg_15_26,
   I2 => M_reg_15_28,
   I3 => W_17_11_i_12_n_0,
   I4 => W_17_11_i_13_n_0,
   O => W_17_11_i_3_n_0
);
W_17_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => M_reg_15_18,
   I1 => M_reg_15_25,
   I2 => M_reg_15_27,
   I3 => W_17_11_i_14_n_0,
   I4 => W_17_11_i_15_n_0,
   O => W_17_11_i_4_n_0
);
W_17_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => M_reg_15_17,
   I1 => M_reg_15_24,
   I2 => M_reg_15_26,
   I3 => W_17_11_i_16_n_0,
   I4 => W_17_11_i_17_n_0,
   O => W_17_11_i_5_n_0
);
W_17_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_17_11_i_2_n_0,
   I1 => W_17_15_i_16_n_0,
   I2 => M_reg_15_21,
   I3 => M_reg_15_28,
   I4 => M_reg_15_30,
   I5 => W_17_15_i_17_n_0,
   O => W_17_11_i_6_n_0
);
W_17_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_17_11_i_3_n_0,
   I1 => W_17_11_i_10_n_0,
   I2 => M_reg_15_20,
   I3 => M_reg_15_27,
   I4 => M_reg_15_29,
   I5 => W_17_11_i_11_n_0,
   O => W_17_11_i_7_n_0
);
W_17_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_17_11_i_4_n_0,
   I1 => W_17_11_i_12_n_0,
   I2 => M_reg_15_19,
   I3 => M_reg_15_26,
   I4 => M_reg_15_28,
   I5 => W_17_11_i_13_n_0,
   O => W_17_11_i_8_n_0
);
W_17_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_17_11_i_5_n_0,
   I1 => W_17_11_i_14_n_0,
   I2 => M_reg_15_18,
   I3 => M_reg_15_25,
   I4 => M_reg_15_27,
   I5 => W_17_11_i_15_n_0,
   O => W_17_11_i_9_n_0
);
W_17_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_1_14,
   I1 => M_reg_10_14,
   I2 => M_reg_2_0,
   I3 => M_reg_2_21,
   I4 => M_reg_2_17,
   O => W_17_15_i_10_n_0
);
W_17_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_10_13,
   I1 => M_reg_2_16,
   I2 => M_reg_2_20,
   I3 => M_reg_2_31,
   I4 => M_reg_1_13,
   O => W_17_15_i_11_n_0
);
W_17_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_1_13,
   I1 => M_reg_10_13,
   I2 => M_reg_2_31,
   I3 => M_reg_2_20,
   I4 => M_reg_2_16,
   O => W_17_15_i_12_n_0
);
W_17_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_10_12,
   I1 => M_reg_2_15,
   I2 => M_reg_2_19,
   I3 => M_reg_2_30,
   I4 => M_reg_1_12,
   O => W_17_15_i_13_n_0
);
W_17_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_1_12,
   I1 => M_reg_10_12,
   I2 => M_reg_2_30,
   I3 => M_reg_2_19,
   I4 => M_reg_2_15,
   O => W_17_15_i_14_n_0
);
W_17_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_10_11,
   I1 => M_reg_2_14,
   I2 => M_reg_2_18,
   I3 => M_reg_2_29,
   I4 => M_reg_1_11,
   O => W_17_15_i_15_n_0
);
W_17_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_1_11,
   I1 => M_reg_10_11,
   I2 => M_reg_2_29,
   I3 => M_reg_2_18,
   I4 => M_reg_2_14,
   O => W_17_15_i_16_n_0
);
W_17_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_10_10,
   I1 => M_reg_2_13,
   I2 => M_reg_2_17,
   I3 => M_reg_2_28,
   I4 => M_reg_1_10,
   O => W_17_15_i_17_n_0
);
W_17_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => M_reg_15_24,
   I1 => M_reg_15_31,
   I2 => M_reg_15_1,
   I3 => W_17_15_i_10_n_0,
   I4 => W_17_15_i_11_n_0,
   O => W_17_15_i_2_n_0
);
W_17_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => M_reg_15_23,
   I1 => M_reg_15_30,
   I2 => M_reg_15_0,
   I3 => W_17_15_i_12_n_0,
   I4 => W_17_15_i_13_n_0,
   O => W_17_15_i_3_n_0
);
W_17_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => M_reg_15_22,
   I1 => M_reg_15_29,
   I2 => M_reg_15_31,
   I3 => W_17_15_i_14_n_0,
   I4 => W_17_15_i_15_n_0,
   O => W_17_15_i_4_n_0
);
W_17_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => M_reg_15_21,
   I1 => M_reg_15_28,
   I2 => M_reg_15_30,
   I3 => W_17_15_i_16_n_0,
   I4 => W_17_15_i_17_n_0,
   O => W_17_15_i_5_n_0
);
W_17_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_17_15_i_2_n_0,
   I1 => W_17_19_i_16_n_0,
   I2 => M_reg_15_25,
   I3 => M_reg_15_0,
   I4 => M_reg_15_2,
   I5 => W_17_19_i_17_n_0,
   O => W_17_15_i_6_n_0
);
W_17_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_17_15_i_3_n_0,
   I1 => W_17_15_i_10_n_0,
   I2 => M_reg_15_24,
   I3 => M_reg_15_31,
   I4 => M_reg_15_1,
   I5 => W_17_15_i_11_n_0,
   O => W_17_15_i_7_n_0
);
W_17_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_17_15_i_4_n_0,
   I1 => W_17_15_i_12_n_0,
   I2 => M_reg_15_23,
   I3 => M_reg_15_30,
   I4 => M_reg_15_0,
   I5 => W_17_15_i_13_n_0,
   O => W_17_15_i_8_n_0
);
W_17_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_17_15_i_5_n_0,
   I1 => W_17_15_i_14_n_0,
   I2 => M_reg_15_22,
   I3 => M_reg_15_29,
   I4 => M_reg_15_31,
   I5 => W_17_15_i_15_n_0,
   O => W_17_15_i_9_n_0
);
W_17_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_1_18,
   I1 => M_reg_10_18,
   I2 => M_reg_2_4,
   I3 => M_reg_2_25,
   I4 => M_reg_2_21,
   O => W_17_19_i_10_n_0
);
W_17_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_10_17,
   I1 => M_reg_2_20,
   I2 => M_reg_2_24,
   I3 => M_reg_2_3,
   I4 => M_reg_1_17,
   O => W_17_19_i_11_n_0
);
W_17_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_1_17,
   I1 => M_reg_10_17,
   I2 => M_reg_2_3,
   I3 => M_reg_2_24,
   I4 => M_reg_2_20,
   O => W_17_19_i_12_n_0
);
W_17_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_10_16,
   I1 => M_reg_2_19,
   I2 => M_reg_2_23,
   I3 => M_reg_2_2,
   I4 => M_reg_1_16,
   O => W_17_19_i_13_n_0
);
W_17_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_1_16,
   I1 => M_reg_10_16,
   I2 => M_reg_2_2,
   I3 => M_reg_2_23,
   I4 => M_reg_2_19,
   O => W_17_19_i_14_n_0
);
W_17_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_10_15,
   I1 => M_reg_2_18,
   I2 => M_reg_2_22,
   I3 => M_reg_2_1,
   I4 => M_reg_1_15,
   O => W_17_19_i_15_n_0
);
W_17_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_1_15,
   I1 => M_reg_10_15,
   I2 => M_reg_2_1,
   I3 => M_reg_2_22,
   I4 => M_reg_2_18,
   O => W_17_19_i_16_n_0
);
W_17_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_10_14,
   I1 => M_reg_2_17,
   I2 => M_reg_2_21,
   I3 => M_reg_2_0,
   I4 => M_reg_1_14,
   O => W_17_19_i_17_n_0
);
W_17_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => M_reg_15_28,
   I1 => M_reg_15_3,
   I2 => M_reg_15_5,
   I3 => W_17_19_i_10_n_0,
   I4 => W_17_19_i_11_n_0,
   O => W_17_19_i_2_n_0
);
W_17_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => M_reg_15_27,
   I1 => M_reg_15_2,
   I2 => M_reg_15_4,
   I3 => W_17_19_i_12_n_0,
   I4 => W_17_19_i_13_n_0,
   O => W_17_19_i_3_n_0
);
W_17_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => M_reg_15_26,
   I1 => M_reg_15_1,
   I2 => M_reg_15_3,
   I3 => W_17_19_i_14_n_0,
   I4 => W_17_19_i_15_n_0,
   O => W_17_19_i_4_n_0
);
W_17_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => M_reg_15_25,
   I1 => M_reg_15_0,
   I2 => M_reg_15_2,
   I3 => W_17_19_i_16_n_0,
   I4 => W_17_19_i_17_n_0,
   O => W_17_19_i_5_n_0
);
W_17_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_17_19_i_2_n_0,
   I1 => W_17_23_i_16_n_0,
   I2 => M_reg_15_29,
   I3 => M_reg_15_4,
   I4 => M_reg_15_6,
   I5 => W_17_23_i_17_n_0,
   O => W_17_19_i_6_n_0
);
W_17_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_17_19_i_3_n_0,
   I1 => W_17_19_i_10_n_0,
   I2 => M_reg_15_28,
   I3 => M_reg_15_3,
   I4 => M_reg_15_5,
   I5 => W_17_19_i_11_n_0,
   O => W_17_19_i_7_n_0
);
W_17_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_17_19_i_4_n_0,
   I1 => W_17_19_i_12_n_0,
   I2 => M_reg_15_27,
   I3 => M_reg_15_2,
   I4 => M_reg_15_4,
   I5 => W_17_19_i_13_n_0,
   O => W_17_19_i_8_n_0
);
W_17_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_17_19_i_5_n_0,
   I1 => W_17_19_i_14_n_0,
   I2 => M_reg_15_26,
   I3 => M_reg_15_1,
   I4 => M_reg_15_3,
   I5 => W_17_19_i_15_n_0,
   O => W_17_19_i_9_n_0
);
W_17_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_1_22,
   I1 => M_reg_10_22,
   I2 => M_reg_2_8,
   I3 => M_reg_2_29,
   I4 => M_reg_2_25,
   O => W_17_23_i_10_n_0
);
W_17_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_10_21,
   I1 => M_reg_2_24,
   I2 => M_reg_2_28,
   I3 => M_reg_2_7,
   I4 => M_reg_1_21,
   O => W_17_23_i_11_n_0
);
W_17_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_1_21,
   I1 => M_reg_10_21,
   I2 => M_reg_2_7,
   I3 => M_reg_2_28,
   I4 => M_reg_2_24,
   O => W_17_23_i_12_n_0
);
W_17_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_10_20,
   I1 => M_reg_2_23,
   I2 => M_reg_2_27,
   I3 => M_reg_2_6,
   I4 => M_reg_1_20,
   O => W_17_23_i_13_n_0
);
W_17_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_1_20,
   I1 => M_reg_10_20,
   I2 => M_reg_2_6,
   I3 => M_reg_2_27,
   I4 => M_reg_2_23,
   O => W_17_23_i_14_n_0
);
W_17_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_10_19,
   I1 => M_reg_2_22,
   I2 => M_reg_2_26,
   I3 => M_reg_2_5,
   I4 => M_reg_1_19,
   O => W_17_23_i_15_n_0
);
W_17_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_1_19,
   I1 => M_reg_10_19,
   I2 => M_reg_2_5,
   I3 => M_reg_2_26,
   I4 => M_reg_2_22,
   O => W_17_23_i_16_n_0
);
W_17_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_10_18,
   I1 => M_reg_2_21,
   I2 => M_reg_2_25,
   I3 => M_reg_2_4,
   I4 => M_reg_1_18,
   O => W_17_23_i_17_n_0
);
W_17_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => M_reg_15_7,
   I1 => M_reg_15_9,
   I2 => W_17_23_i_10_n_0,
   I3 => W_17_23_i_11_n_0,
   O => W_17_23_i_2_n_0
);
W_17_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => M_reg_15_31,
   I1 => M_reg_15_6,
   I2 => M_reg_15_8,
   I3 => W_17_23_i_12_n_0,
   I4 => W_17_23_i_13_n_0,
   O => W_17_23_i_3_n_0
);
W_17_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => M_reg_15_30,
   I1 => M_reg_15_5,
   I2 => M_reg_15_7,
   I3 => W_17_23_i_14_n_0,
   I4 => W_17_23_i_15_n_0,
   O => W_17_23_i_4_n_0
);
W_17_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => M_reg_15_29,
   I1 => M_reg_15_4,
   I2 => M_reg_15_6,
   I3 => W_17_23_i_16_n_0,
   I4 => W_17_23_i_17_n_0,
   O => W_17_23_i_5_n_0
);
W_17_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_15_8,
   I1 => M_reg_15_10,
   I2 => W_17_27_i_16_n_0,
   I3 => W_17_27_i_17_n_0,
   I4 => W_17_23_i_2_n_0,
   O => W_17_23_i_6_n_0
);
W_17_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_15_7,
   I1 => M_reg_15_9,
   I2 => W_17_23_i_10_n_0,
   I3 => W_17_23_i_11_n_0,
   I4 => W_17_23_i_3_n_0,
   O => W_17_23_i_7_n_0
);
W_17_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_17_23_i_4_n_0,
   I1 => W_17_23_i_12_n_0,
   I2 => M_reg_15_31,
   I3 => M_reg_15_6,
   I4 => M_reg_15_8,
   I5 => W_17_23_i_13_n_0,
   O => W_17_23_i_8_n_0
);
W_17_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_17_23_i_5_n_0,
   I1 => W_17_23_i_14_n_0,
   I2 => M_reg_15_30,
   I3 => M_reg_15_5,
   I4 => M_reg_15_7,
   I5 => W_17_23_i_15_n_0,
   O => W_17_23_i_9_n_0
);
W_17_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_1_26,
   I1 => M_reg_10_26,
   I2 => M_reg_2_12,
   I3 => M_reg_2_1,
   I4 => M_reg_2_29,
   O => W_17_27_i_10_n_0
);
W_17_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_10_25,
   I1 => M_reg_2_28,
   I2 => M_reg_2_0,
   I3 => M_reg_2_11,
   I4 => M_reg_1_25,
   O => W_17_27_i_11_n_0
);
W_17_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_1_25,
   I1 => M_reg_10_25,
   I2 => M_reg_2_11,
   I3 => M_reg_2_0,
   I4 => M_reg_2_28,
   O => W_17_27_i_12_n_0
);
W_17_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_10_24,
   I1 => M_reg_2_27,
   I2 => M_reg_2_31,
   I3 => M_reg_2_10,
   I4 => M_reg_1_24,
   O => W_17_27_i_13_n_0
);
W_17_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_1_24,
   I1 => M_reg_10_24,
   I2 => M_reg_2_10,
   I3 => M_reg_2_31,
   I4 => M_reg_2_27,
   O => W_17_27_i_14_n_0
);
W_17_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_10_23,
   I1 => M_reg_2_26,
   I2 => M_reg_2_30,
   I3 => M_reg_2_9,
   I4 => M_reg_1_23,
   O => W_17_27_i_15_n_0
);
W_17_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_1_23,
   I1 => M_reg_10_23,
   I2 => M_reg_2_9,
   I3 => M_reg_2_30,
   I4 => M_reg_2_26,
   O => W_17_27_i_16_n_0
);
W_17_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_10_22,
   I1 => M_reg_2_25,
   I2 => M_reg_2_29,
   I3 => M_reg_2_8,
   I4 => M_reg_1_22,
   O => W_17_27_i_17_n_0
);
W_17_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => M_reg_15_11,
   I1 => M_reg_15_13,
   I2 => W_17_27_i_10_n_0,
   I3 => W_17_27_i_11_n_0,
   O => W_17_27_i_2_n_0
);
W_17_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => M_reg_15_10,
   I1 => M_reg_15_12,
   I2 => W_17_27_i_12_n_0,
   I3 => W_17_27_i_13_n_0,
   O => W_17_27_i_3_n_0
);
W_17_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => M_reg_15_9,
   I1 => M_reg_15_11,
   I2 => W_17_27_i_14_n_0,
   I3 => W_17_27_i_15_n_0,
   O => W_17_27_i_4_n_0
);
W_17_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => M_reg_15_8,
   I1 => M_reg_15_10,
   I2 => W_17_27_i_16_n_0,
   I3 => W_17_27_i_17_n_0,
   O => W_17_27_i_5_n_0
);
W_17_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_15_12,
   I1 => M_reg_15_14,
   I2 => W_17_31_i_13_n_0,
   I3 => W_17_31_i_14_n_0,
   I4 => W_17_27_i_2_n_0,
   O => W_17_27_i_6_n_0
);
W_17_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_15_11,
   I1 => M_reg_15_13,
   I2 => W_17_27_i_10_n_0,
   I3 => W_17_27_i_11_n_0,
   I4 => W_17_27_i_3_n_0,
   O => W_17_27_i_7_n_0
);
W_17_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_15_10,
   I1 => M_reg_15_12,
   I2 => W_17_27_i_12_n_0,
   I3 => W_17_27_i_13_n_0,
   I4 => W_17_27_i_4_n_0,
   O => W_17_27_i_8_n_0
);
W_17_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_15_9,
   I1 => M_reg_15_11,
   I2 => W_17_27_i_14_n_0,
   I3 => W_17_27_i_15_n_0,
   I4 => W_17_27_i_5_n_0,
   O => W_17_27_i_9_n_0
);
W_17_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_10_28,
   I1 => M_reg_2_31,
   I2 => M_reg_2_3,
   I3 => M_reg_2_14,
   I4 => M_reg_1_28,
   O => W_17_31_i_10_n_0
);
W_17_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_1_28,
   I1 => M_reg_10_28,
   I2 => M_reg_2_14,
   I3 => M_reg_2_3,
   I4 => M_reg_2_31,
   O => W_17_31_i_11_n_0
);
W_17_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_10_27,
   I1 => M_reg_2_30,
   I2 => M_reg_2_2,
   I3 => M_reg_2_13,
   I4 => M_reg_1_27,
   O => W_17_31_i_12_n_0
);
W_17_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_1_27,
   I1 => M_reg_10_27,
   I2 => M_reg_2_13,
   I3 => M_reg_2_2,
   I4 => M_reg_2_30,
   O => W_17_31_i_13_n_0
);
W_17_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_10_26,
   I1 => M_reg_2_29,
   I2 => M_reg_2_1,
   I3 => M_reg_2_12,
   I4 => M_reg_1_26,
   O => W_17_31_i_14_n_0
);
W_17_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => M_reg_10_29,
   I1 => M_reg_2_4,
   I2 => M_reg_2_15,
   I3 => M_reg_1_29,
   O => W_17_31_i_15_n_0
);
W_17_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => M_reg_15_17,
   I1 => M_reg_15_15,
   O => SIGMA_LCASE_1379_out_30
);
W_17_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => M_reg_2_6,
   I1 => M_reg_2_17,
   I2 => M_reg_10_31,
   I3 => M_reg_1_31,
   I4 => M_reg_15_16,
   I5 => M_reg_15_18,
   O => W_17_31_i_17_n_0
);
W_17_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => M_reg_2_16,
   I1 => M_reg_2_5,
   O => SIGMA_LCASE_0375_out_30
);
W_17_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => M_reg_1_30,
   I1 => M_reg_10_30,
   I2 => M_reg_2_16,
   I3 => M_reg_2_5,
   O => W_17_31_i_19_n_0
);
W_17_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => M_reg_15_14,
   I1 => M_reg_15_16,
   I2 => W_17_31_i_9_n_0,
   I3 => W_17_31_i_10_n_0,
   O => W_17_31_i_2_n_0
);
W_17_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => M_reg_15_13,
   I1 => M_reg_15_15,
   I2 => W_17_31_i_11_n_0,
   I3 => W_17_31_i_12_n_0,
   O => W_17_31_i_3_n_0
);
W_17_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => M_reg_15_12,
   I1 => M_reg_15_14,
   I2 => W_17_31_i_13_n_0,
   I3 => W_17_31_i_14_n_0,
   O => W_17_31_i_4_n_0
);
W_17_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_17_31_i_15_n_0,
   I1 => SIGMA_LCASE_1379_out_30,
   I2 => W_17_31_i_17_n_0,
   I3 => M_reg_10_30,
   I4 => SIGMA_LCASE_0375_out_30,
   I5 => M_reg_1_30,
   O => W_17_31_i_5_n_0
);
W_17_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_17_31_i_2_n_0,
   I1 => W_17_31_i_19_n_0,
   I2 => M_reg_15_15,
   I3 => M_reg_15_17,
   I4 => W_17_31_i_15_n_0,
   O => W_17_31_i_6_n_0
);
W_17_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_15_14,
   I1 => M_reg_15_16,
   I2 => W_17_31_i_9_n_0,
   I3 => W_17_31_i_10_n_0,
   I4 => W_17_31_i_3_n_0,
   O => W_17_31_i_7_n_0
);
W_17_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_15_13,
   I1 => M_reg_15_15,
   I2 => W_17_31_i_11_n_0,
   I3 => W_17_31_i_12_n_0,
   I4 => W_17_31_i_4_n_0,
   O => W_17_31_i_8_n_0
);
W_17_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => M_reg_1_29,
   I1 => M_reg_10_29,
   I2 => M_reg_2_15,
   I3 => M_reg_2_4,
   O => W_17_31_i_9_n_0
);
W_17_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_1_2,
   I1 => M_reg_10_2,
   I2 => M_reg_2_20,
   I3 => M_reg_2_9,
   I4 => M_reg_2_5,
   O => W_17_3_i_10_n_0
);
W_17_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_10_1,
   I1 => M_reg_2_4,
   I2 => M_reg_2_8,
   I3 => M_reg_2_19,
   I4 => M_reg_1_1,
   O => W_17_3_i_11_n_0
);
W_17_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => M_reg_2_19,
   I1 => M_reg_2_8,
   I2 => M_reg_2_4,
   O => SIGMA_LCASE_0375_out_1
);
W_17_3_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_1_1,
   I1 => M_reg_10_1,
   I2 => M_reg_2_19,
   I3 => M_reg_2_8,
   I4 => M_reg_2_4,
   O => W_17_3_i_13_n_0
);
W_17_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => M_reg_15_12,
   I1 => M_reg_15_19,
   I2 => M_reg_15_21,
   I3 => W_17_3_i_10_n_0,
   I4 => W_17_3_i_11_n_0,
   O => W_17_3_i_2_n_0
);
W_17_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_17_3_i_11_n_0,
   I1 => M_reg_15_21,
   I2 => M_reg_15_19,
   I3 => M_reg_15_12,
   I4 => W_17_3_i_10_n_0,
   O => W_17_3_i_3_n_0
);
W_17_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_0375_out_1,
   I1 => M_reg_10_1,
   I2 => M_reg_1_1,
   I3 => M_reg_15_11,
   I4 => M_reg_15_18,
   I5 => M_reg_15_20,
   O => W_17_3_i_4_n_0
);
W_17_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_1_0,
   I1 => M_reg_10_0,
   I2 => M_reg_2_18,
   I3 => M_reg_2_7,
   I4 => M_reg_2_3,
   O => W_17_3_i_5_n_0
);
W_17_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_17_3_i_2_n_0,
   I1 => W_17_7_i_16_n_0,
   I2 => M_reg_15_13,
   I3 => M_reg_15_20,
   I4 => M_reg_15_22,
   I5 => W_17_7_i_17_n_0,
   O => W_17_3_i_6_n_0
);
W_17_3_i_7 : LUT5
  generic map(
   INIT => X"6aa6a66a"
  )
 port map (
   I0 => W_17_3_i_3_n_0,
   I1 => W_17_3_i_13_n_0,
   I2 => M_reg_15_20,
   I3 => M_reg_15_18,
   I4 => M_reg_15_11,
   O => W_17_3_i_7_n_0
);
W_17_3_i_8 : LUT6
  generic map(
   INIT => X"566565566aa6a66a"
  )
 port map (
   I0 => W_17_3_i_4_n_0,
   I1 => M_reg_1_0,
   I2 => M_reg_2_18,
   I3 => M_reg_2_7,
   I4 => M_reg_2_3,
   I5 => M_reg_10_0,
   O => W_17_3_i_8_n_0
);
W_17_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_17_3_i_5_n_0,
   I1 => M_reg_15_10,
   I2 => M_reg_15_17,
   I3 => M_reg_15_19,
   O => W_17_3_i_9_n_0
);
W_17_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_1_6,
   I1 => M_reg_10_6,
   I2 => M_reg_2_24,
   I3 => M_reg_2_13,
   I4 => M_reg_2_9,
   O => W_17_7_i_10_n_0
);
W_17_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_10_5,
   I1 => M_reg_2_8,
   I2 => M_reg_2_12,
   I3 => M_reg_2_23,
   I4 => M_reg_1_5,
   O => W_17_7_i_11_n_0
);
W_17_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_1_5,
   I1 => M_reg_10_5,
   I2 => M_reg_2_23,
   I3 => M_reg_2_12,
   I4 => M_reg_2_8,
   O => W_17_7_i_12_n_0
);
W_17_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_10_4,
   I1 => M_reg_2_7,
   I2 => M_reg_2_11,
   I3 => M_reg_2_22,
   I4 => M_reg_1_4,
   O => W_17_7_i_13_n_0
);
W_17_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_1_4,
   I1 => M_reg_10_4,
   I2 => M_reg_2_22,
   I3 => M_reg_2_11,
   I4 => M_reg_2_7,
   O => W_17_7_i_14_n_0
);
W_17_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_10_3,
   I1 => M_reg_2_6,
   I2 => M_reg_2_10,
   I3 => M_reg_2_21,
   I4 => M_reg_1_3,
   O => W_17_7_i_15_n_0
);
W_17_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_1_3,
   I1 => M_reg_10_3,
   I2 => M_reg_2_21,
   I3 => M_reg_2_10,
   I4 => M_reg_2_6,
   O => W_17_7_i_16_n_0
);
W_17_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_10_2,
   I1 => M_reg_2_5,
   I2 => M_reg_2_9,
   I3 => M_reg_2_20,
   I4 => M_reg_1_2,
   O => W_17_7_i_17_n_0
);
W_17_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => M_reg_15_16,
   I1 => M_reg_15_23,
   I2 => M_reg_15_25,
   I3 => W_17_7_i_10_n_0,
   I4 => W_17_7_i_11_n_0,
   O => W_17_7_i_2_n_0
);
W_17_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => M_reg_15_15,
   I1 => M_reg_15_22,
   I2 => M_reg_15_24,
   I3 => W_17_7_i_12_n_0,
   I4 => W_17_7_i_13_n_0,
   O => W_17_7_i_3_n_0
);
W_17_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => M_reg_15_14,
   I1 => M_reg_15_21,
   I2 => M_reg_15_23,
   I3 => W_17_7_i_14_n_0,
   I4 => W_17_7_i_15_n_0,
   O => W_17_7_i_4_n_0
);
W_17_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => M_reg_15_13,
   I1 => M_reg_15_20,
   I2 => M_reg_15_22,
   I3 => W_17_7_i_16_n_0,
   I4 => W_17_7_i_17_n_0,
   O => W_17_7_i_5_n_0
);
W_17_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_17_7_i_2_n_0,
   I1 => W_17_11_i_16_n_0,
   I2 => M_reg_15_17,
   I3 => M_reg_15_24,
   I4 => M_reg_15_26,
   I5 => W_17_11_i_17_n_0,
   O => W_17_7_i_6_n_0
);
W_17_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_17_7_i_3_n_0,
   I1 => W_17_7_i_10_n_0,
   I2 => M_reg_15_16,
   I3 => M_reg_15_23,
   I4 => M_reg_15_25,
   I5 => W_17_7_i_11_n_0,
   O => W_17_7_i_7_n_0
);
W_17_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_17_7_i_4_n_0,
   I1 => W_17_7_i_12_n_0,
   I2 => M_reg_15_15,
   I3 => M_reg_15_22,
   I4 => M_reg_15_24,
   I5 => W_17_7_i_13_n_0,
   O => W_17_7_i_8_n_0
);
W_17_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_17_7_i_5_n_0,
   I1 => W_17_7_i_14_n_0,
   I2 => M_reg_15_14,
   I3 => M_reg_15_21,
   I4 => M_reg_15_23,
   I5 => W_17_7_i_15_n_0,
   O => W_17_7_i_9_n_0
);
W_18_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_2_10,
   I1 => M_reg_11_10,
   I2 => M_reg_3_28,
   I3 => M_reg_3_17,
   I4 => M_reg_3_13,
   O => W_18_11_i_10_n_0
);
W_18_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_11_9,
   I1 => M_reg_3_12,
   I2 => M_reg_3_16,
   I3 => M_reg_3_27,
   I4 => M_reg_2_9,
   O => W_18_11_i_11_n_0
);
W_18_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_2_9,
   I1 => M_reg_11_9,
   I2 => M_reg_3_27,
   I3 => M_reg_3_16,
   I4 => M_reg_3_12,
   O => W_18_11_i_12_n_0
);
W_18_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_11_8,
   I1 => M_reg_3_11,
   I2 => M_reg_3_15,
   I3 => M_reg_3_26,
   I4 => M_reg_2_8,
   O => W_18_11_i_13_n_0
);
W_18_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_2_8,
   I1 => M_reg_11_8,
   I2 => M_reg_3_26,
   I3 => M_reg_3_15,
   I4 => M_reg_3_11,
   O => W_18_11_i_14_n_0
);
W_18_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_11_7,
   I1 => M_reg_3_10,
   I2 => M_reg_3_14,
   I3 => M_reg_3_25,
   I4 => M_reg_2_7,
   O => W_18_11_i_15_n_0
);
W_18_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_2_7,
   I1 => M_reg_11_7,
   I2 => M_reg_3_25,
   I3 => M_reg_3_14,
   I4 => M_reg_3_10,
   O => W_18_11_i_16_n_0
);
W_18_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_11_6,
   I1 => M_reg_3_9,
   I2 => M_reg_3_13,
   I3 => M_reg_3_24,
   I4 => M_reg_2_6,
   O => W_18_11_i_17_n_0
);
W_18_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x117_out_20,
   I1 => x117_out_27,
   I2 => x117_out_29,
   I3 => W_18_11_i_10_n_0,
   I4 => W_18_11_i_11_n_0,
   O => W_18_11_i_2_n_0
);
W_18_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x117_out_19,
   I1 => x117_out_26,
   I2 => x117_out_28,
   I3 => W_18_11_i_12_n_0,
   I4 => W_18_11_i_13_n_0,
   O => W_18_11_i_3_n_0
);
W_18_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x117_out_18,
   I1 => x117_out_25,
   I2 => x117_out_27,
   I3 => W_18_11_i_14_n_0,
   I4 => W_18_11_i_15_n_0,
   O => W_18_11_i_4_n_0
);
W_18_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x117_out_17,
   I1 => x117_out_24,
   I2 => x117_out_26,
   I3 => W_18_11_i_16_n_0,
   I4 => W_18_11_i_17_n_0,
   O => W_18_11_i_5_n_0
);
W_18_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_18_11_i_2_n_0,
   I1 => W_18_15_i_16_n_0,
   I2 => x117_out_21,
   I3 => x117_out_28,
   I4 => x117_out_30,
   I5 => W_18_15_i_17_n_0,
   O => W_18_11_i_6_n_0
);
W_18_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_18_11_i_3_n_0,
   I1 => W_18_11_i_10_n_0,
   I2 => x117_out_20,
   I3 => x117_out_27,
   I4 => x117_out_29,
   I5 => W_18_11_i_11_n_0,
   O => W_18_11_i_7_n_0
);
W_18_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_18_11_i_4_n_0,
   I1 => W_18_11_i_12_n_0,
   I2 => x117_out_19,
   I3 => x117_out_26,
   I4 => x117_out_28,
   I5 => W_18_11_i_13_n_0,
   O => W_18_11_i_8_n_0
);
W_18_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_18_11_i_5_n_0,
   I1 => W_18_11_i_14_n_0,
   I2 => x117_out_18,
   I3 => x117_out_25,
   I4 => x117_out_27,
   I5 => W_18_11_i_15_n_0,
   O => W_18_11_i_9_n_0
);
W_18_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_2_14,
   I1 => M_reg_11_14,
   I2 => M_reg_3_0,
   I3 => M_reg_3_21,
   I4 => M_reg_3_17,
   O => W_18_15_i_10_n_0
);
W_18_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_11_13,
   I1 => M_reg_3_16,
   I2 => M_reg_3_20,
   I3 => M_reg_3_31,
   I4 => M_reg_2_13,
   O => W_18_15_i_11_n_0
);
W_18_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_2_13,
   I1 => M_reg_11_13,
   I2 => M_reg_3_31,
   I3 => M_reg_3_20,
   I4 => M_reg_3_16,
   O => W_18_15_i_12_n_0
);
W_18_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_11_12,
   I1 => M_reg_3_15,
   I2 => M_reg_3_19,
   I3 => M_reg_3_30,
   I4 => M_reg_2_12,
   O => W_18_15_i_13_n_0
);
W_18_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_2_12,
   I1 => M_reg_11_12,
   I2 => M_reg_3_30,
   I3 => M_reg_3_19,
   I4 => M_reg_3_15,
   O => W_18_15_i_14_n_0
);
W_18_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_11_11,
   I1 => M_reg_3_14,
   I2 => M_reg_3_18,
   I3 => M_reg_3_29,
   I4 => M_reg_2_11,
   O => W_18_15_i_15_n_0
);
W_18_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_2_11,
   I1 => M_reg_11_11,
   I2 => M_reg_3_29,
   I3 => M_reg_3_18,
   I4 => M_reg_3_14,
   O => W_18_15_i_16_n_0
);
W_18_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_11_10,
   I1 => M_reg_3_13,
   I2 => M_reg_3_17,
   I3 => M_reg_3_28,
   I4 => M_reg_2_10,
   O => W_18_15_i_17_n_0
);
W_18_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x117_out_24,
   I1 => x117_out_31,
   I2 => x117_out_1,
   I3 => W_18_15_i_10_n_0,
   I4 => W_18_15_i_11_n_0,
   O => W_18_15_i_2_n_0
);
W_18_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x117_out_23,
   I1 => x117_out_30,
   I2 => x117_out_0,
   I3 => W_18_15_i_12_n_0,
   I4 => W_18_15_i_13_n_0,
   O => W_18_15_i_3_n_0
);
W_18_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x117_out_22,
   I1 => x117_out_29,
   I2 => x117_out_31,
   I3 => W_18_15_i_14_n_0,
   I4 => W_18_15_i_15_n_0,
   O => W_18_15_i_4_n_0
);
W_18_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x117_out_21,
   I1 => x117_out_28,
   I2 => x117_out_30,
   I3 => W_18_15_i_16_n_0,
   I4 => W_18_15_i_17_n_0,
   O => W_18_15_i_5_n_0
);
W_18_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_18_15_i_2_n_0,
   I1 => W_18_19_i_16_n_0,
   I2 => x117_out_25,
   I3 => x117_out_0,
   I4 => x117_out_2,
   I5 => W_18_19_i_17_n_0,
   O => W_18_15_i_6_n_0
);
W_18_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_18_15_i_3_n_0,
   I1 => W_18_15_i_10_n_0,
   I2 => x117_out_24,
   I3 => x117_out_31,
   I4 => x117_out_1,
   I5 => W_18_15_i_11_n_0,
   O => W_18_15_i_7_n_0
);
W_18_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_18_15_i_4_n_0,
   I1 => W_18_15_i_12_n_0,
   I2 => x117_out_23,
   I3 => x117_out_30,
   I4 => x117_out_0,
   I5 => W_18_15_i_13_n_0,
   O => W_18_15_i_8_n_0
);
W_18_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_18_15_i_5_n_0,
   I1 => W_18_15_i_14_n_0,
   I2 => x117_out_22,
   I3 => x117_out_29,
   I4 => x117_out_31,
   I5 => W_18_15_i_15_n_0,
   O => W_18_15_i_9_n_0
);
W_18_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_2_18,
   I1 => M_reg_11_18,
   I2 => M_reg_3_4,
   I3 => M_reg_3_25,
   I4 => M_reg_3_21,
   O => W_18_19_i_10_n_0
);
W_18_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_11_17,
   I1 => M_reg_3_20,
   I2 => M_reg_3_24,
   I3 => M_reg_3_3,
   I4 => M_reg_2_17,
   O => W_18_19_i_11_n_0
);
W_18_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_2_17,
   I1 => M_reg_11_17,
   I2 => M_reg_3_3,
   I3 => M_reg_3_24,
   I4 => M_reg_3_20,
   O => W_18_19_i_12_n_0
);
W_18_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_11_16,
   I1 => M_reg_3_19,
   I2 => M_reg_3_23,
   I3 => M_reg_3_2,
   I4 => M_reg_2_16,
   O => W_18_19_i_13_n_0
);
W_18_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_2_16,
   I1 => M_reg_11_16,
   I2 => M_reg_3_2,
   I3 => M_reg_3_23,
   I4 => M_reg_3_19,
   O => W_18_19_i_14_n_0
);
W_18_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_11_15,
   I1 => M_reg_3_18,
   I2 => M_reg_3_22,
   I3 => M_reg_3_1,
   I4 => M_reg_2_15,
   O => W_18_19_i_15_n_0
);
W_18_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_2_15,
   I1 => M_reg_11_15,
   I2 => M_reg_3_1,
   I3 => M_reg_3_22,
   I4 => M_reg_3_18,
   O => W_18_19_i_16_n_0
);
W_18_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_11_14,
   I1 => M_reg_3_17,
   I2 => M_reg_3_21,
   I3 => M_reg_3_0,
   I4 => M_reg_2_14,
   O => W_18_19_i_17_n_0
);
W_18_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x117_out_28,
   I1 => x117_out_3,
   I2 => x117_out_5,
   I3 => W_18_19_i_10_n_0,
   I4 => W_18_19_i_11_n_0,
   O => W_18_19_i_2_n_0
);
W_18_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x117_out_27,
   I1 => x117_out_2,
   I2 => x117_out_4,
   I3 => W_18_19_i_12_n_0,
   I4 => W_18_19_i_13_n_0,
   O => W_18_19_i_3_n_0
);
W_18_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x117_out_26,
   I1 => x117_out_1,
   I2 => x117_out_3,
   I3 => W_18_19_i_14_n_0,
   I4 => W_18_19_i_15_n_0,
   O => W_18_19_i_4_n_0
);
W_18_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x117_out_25,
   I1 => x117_out_0,
   I2 => x117_out_2,
   I3 => W_18_19_i_16_n_0,
   I4 => W_18_19_i_17_n_0,
   O => W_18_19_i_5_n_0
);
W_18_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_18_19_i_2_n_0,
   I1 => W_18_23_i_16_n_0,
   I2 => x117_out_29,
   I3 => x117_out_4,
   I4 => x117_out_6,
   I5 => W_18_23_i_17_n_0,
   O => W_18_19_i_6_n_0
);
W_18_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_18_19_i_3_n_0,
   I1 => W_18_19_i_10_n_0,
   I2 => x117_out_28,
   I3 => x117_out_3,
   I4 => x117_out_5,
   I5 => W_18_19_i_11_n_0,
   O => W_18_19_i_7_n_0
);
W_18_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_18_19_i_4_n_0,
   I1 => W_18_19_i_12_n_0,
   I2 => x117_out_27,
   I3 => x117_out_2,
   I4 => x117_out_4,
   I5 => W_18_19_i_13_n_0,
   O => W_18_19_i_8_n_0
);
W_18_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_18_19_i_5_n_0,
   I1 => W_18_19_i_14_n_0,
   I2 => x117_out_26,
   I3 => x117_out_1,
   I4 => x117_out_3,
   I5 => W_18_19_i_15_n_0,
   O => W_18_19_i_9_n_0
);
W_18_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_2_22,
   I1 => M_reg_11_22,
   I2 => M_reg_3_8,
   I3 => M_reg_3_29,
   I4 => M_reg_3_25,
   O => W_18_23_i_10_n_0
);
W_18_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_11_21,
   I1 => M_reg_3_24,
   I2 => M_reg_3_28,
   I3 => M_reg_3_7,
   I4 => M_reg_2_21,
   O => W_18_23_i_11_n_0
);
W_18_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_2_21,
   I1 => M_reg_11_21,
   I2 => M_reg_3_7,
   I3 => M_reg_3_28,
   I4 => M_reg_3_24,
   O => W_18_23_i_12_n_0
);
W_18_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_11_20,
   I1 => M_reg_3_23,
   I2 => M_reg_3_27,
   I3 => M_reg_3_6,
   I4 => M_reg_2_20,
   O => W_18_23_i_13_n_0
);
W_18_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_2_20,
   I1 => M_reg_11_20,
   I2 => M_reg_3_6,
   I3 => M_reg_3_27,
   I4 => M_reg_3_23,
   O => W_18_23_i_14_n_0
);
W_18_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_11_19,
   I1 => M_reg_3_22,
   I2 => M_reg_3_26,
   I3 => M_reg_3_5,
   I4 => M_reg_2_19,
   O => W_18_23_i_15_n_0
);
W_18_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_2_19,
   I1 => M_reg_11_19,
   I2 => M_reg_3_5,
   I3 => M_reg_3_26,
   I4 => M_reg_3_22,
   O => W_18_23_i_16_n_0
);
W_18_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_11_18,
   I1 => M_reg_3_21,
   I2 => M_reg_3_25,
   I3 => M_reg_3_4,
   I4 => M_reg_2_18,
   O => W_18_23_i_17_n_0
);
W_18_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x117_out_7,
   I1 => x117_out_9,
   I2 => W_18_23_i_10_n_0,
   I3 => W_18_23_i_11_n_0,
   O => W_18_23_i_2_n_0
);
W_18_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x117_out_31,
   I1 => x117_out_6,
   I2 => x117_out_8,
   I3 => W_18_23_i_12_n_0,
   I4 => W_18_23_i_13_n_0,
   O => W_18_23_i_3_n_0
);
W_18_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x117_out_30,
   I1 => x117_out_5,
   I2 => x117_out_7,
   I3 => W_18_23_i_14_n_0,
   I4 => W_18_23_i_15_n_0,
   O => W_18_23_i_4_n_0
);
W_18_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x117_out_29,
   I1 => x117_out_4,
   I2 => x117_out_6,
   I3 => W_18_23_i_16_n_0,
   I4 => W_18_23_i_17_n_0,
   O => W_18_23_i_5_n_0
);
W_18_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x117_out_8,
   I1 => x117_out_10,
   I2 => W_18_27_i_16_n_0,
   I3 => W_18_27_i_17_n_0,
   I4 => W_18_23_i_2_n_0,
   O => W_18_23_i_6_n_0
);
W_18_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x117_out_7,
   I1 => x117_out_9,
   I2 => W_18_23_i_10_n_0,
   I3 => W_18_23_i_11_n_0,
   I4 => W_18_23_i_3_n_0,
   O => W_18_23_i_7_n_0
);
W_18_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_18_23_i_4_n_0,
   I1 => W_18_23_i_12_n_0,
   I2 => x117_out_31,
   I3 => x117_out_6,
   I4 => x117_out_8,
   I5 => W_18_23_i_13_n_0,
   O => W_18_23_i_8_n_0
);
W_18_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_18_23_i_5_n_0,
   I1 => W_18_23_i_14_n_0,
   I2 => x117_out_30,
   I3 => x117_out_5,
   I4 => x117_out_7,
   I5 => W_18_23_i_15_n_0,
   O => W_18_23_i_9_n_0
);
W_18_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_2_26,
   I1 => M_reg_11_26,
   I2 => M_reg_3_12,
   I3 => M_reg_3_1,
   I4 => M_reg_3_29,
   O => W_18_27_i_10_n_0
);
W_18_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_11_25,
   I1 => M_reg_3_28,
   I2 => M_reg_3_0,
   I3 => M_reg_3_11,
   I4 => M_reg_2_25,
   O => W_18_27_i_11_n_0
);
W_18_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_2_25,
   I1 => M_reg_11_25,
   I2 => M_reg_3_11,
   I3 => M_reg_3_0,
   I4 => M_reg_3_28,
   O => W_18_27_i_12_n_0
);
W_18_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_11_24,
   I1 => M_reg_3_27,
   I2 => M_reg_3_31,
   I3 => M_reg_3_10,
   I4 => M_reg_2_24,
   O => W_18_27_i_13_n_0
);
W_18_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_2_24,
   I1 => M_reg_11_24,
   I2 => M_reg_3_10,
   I3 => M_reg_3_31,
   I4 => M_reg_3_27,
   O => W_18_27_i_14_n_0
);
W_18_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_11_23,
   I1 => M_reg_3_26,
   I2 => M_reg_3_30,
   I3 => M_reg_3_9,
   I4 => M_reg_2_23,
   O => W_18_27_i_15_n_0
);
W_18_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_2_23,
   I1 => M_reg_11_23,
   I2 => M_reg_3_9,
   I3 => M_reg_3_30,
   I4 => M_reg_3_26,
   O => W_18_27_i_16_n_0
);
W_18_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_11_22,
   I1 => M_reg_3_25,
   I2 => M_reg_3_29,
   I3 => M_reg_3_8,
   I4 => M_reg_2_22,
   O => W_18_27_i_17_n_0
);
W_18_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x117_out_11,
   I1 => x117_out_13,
   I2 => W_18_27_i_10_n_0,
   I3 => W_18_27_i_11_n_0,
   O => W_18_27_i_2_n_0
);
W_18_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x117_out_10,
   I1 => x117_out_12,
   I2 => W_18_27_i_12_n_0,
   I3 => W_18_27_i_13_n_0,
   O => W_18_27_i_3_n_0
);
W_18_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x117_out_9,
   I1 => x117_out_11,
   I2 => W_18_27_i_14_n_0,
   I3 => W_18_27_i_15_n_0,
   O => W_18_27_i_4_n_0
);
W_18_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x117_out_8,
   I1 => x117_out_10,
   I2 => W_18_27_i_16_n_0,
   I3 => W_18_27_i_17_n_0,
   O => W_18_27_i_5_n_0
);
W_18_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x117_out_12,
   I1 => x117_out_14,
   I2 => W_18_31_i_13_n_0,
   I3 => W_18_31_i_14_n_0,
   I4 => W_18_27_i_2_n_0,
   O => W_18_27_i_6_n_0
);
W_18_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x117_out_11,
   I1 => x117_out_13,
   I2 => W_18_27_i_10_n_0,
   I3 => W_18_27_i_11_n_0,
   I4 => W_18_27_i_3_n_0,
   O => W_18_27_i_7_n_0
);
W_18_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x117_out_10,
   I1 => x117_out_12,
   I2 => W_18_27_i_12_n_0,
   I3 => W_18_27_i_13_n_0,
   I4 => W_18_27_i_4_n_0,
   O => W_18_27_i_8_n_0
);
W_18_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x117_out_9,
   I1 => x117_out_11,
   I2 => W_18_27_i_14_n_0,
   I3 => W_18_27_i_15_n_0,
   I4 => W_18_27_i_5_n_0,
   O => W_18_27_i_9_n_0
);
W_18_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_11_28,
   I1 => M_reg_3_31,
   I2 => M_reg_3_3,
   I3 => M_reg_3_14,
   I4 => M_reg_2_28,
   O => W_18_31_i_10_n_0
);
W_18_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_2_28,
   I1 => M_reg_11_28,
   I2 => M_reg_3_14,
   I3 => M_reg_3_3,
   I4 => M_reg_3_31,
   O => W_18_31_i_11_n_0
);
W_18_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_11_27,
   I1 => M_reg_3_30,
   I2 => M_reg_3_2,
   I3 => M_reg_3_13,
   I4 => M_reg_2_27,
   O => W_18_31_i_12_n_0
);
W_18_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_2_27,
   I1 => M_reg_11_27,
   I2 => M_reg_3_13,
   I3 => M_reg_3_2,
   I4 => M_reg_3_30,
   O => W_18_31_i_13_n_0
);
W_18_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_11_26,
   I1 => M_reg_3_29,
   I2 => M_reg_3_1,
   I3 => M_reg_3_12,
   I4 => M_reg_2_26,
   O => W_18_31_i_14_n_0
);
W_18_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => M_reg_11_29,
   I1 => M_reg_3_4,
   I2 => M_reg_3_15,
   I3 => M_reg_2_29,
   O => W_18_31_i_15_n_0
);
W_18_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x117_out_17,
   I1 => x117_out_15,
   O => SIGMA_LCASE_1371_out_30
);
W_18_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => M_reg_3_6,
   I1 => M_reg_3_17,
   I2 => M_reg_11_31,
   I3 => M_reg_2_31,
   I4 => x117_out_16,
   I5 => x117_out_18,
   O => W_18_31_i_17_n_0
);
W_18_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => M_reg_3_16,
   I1 => M_reg_3_5,
   O => SIGMA_LCASE_0367_out_30
);
W_18_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => M_reg_2_30,
   I1 => M_reg_11_30,
   I2 => M_reg_3_16,
   I3 => M_reg_3_5,
   O => W_18_31_i_19_n_0
);
W_18_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x117_out_14,
   I1 => x117_out_16,
   I2 => W_18_31_i_9_n_0,
   I3 => W_18_31_i_10_n_0,
   O => W_18_31_i_2_n_0
);
W_18_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x117_out_13,
   I1 => x117_out_15,
   I2 => W_18_31_i_11_n_0,
   I3 => W_18_31_i_12_n_0,
   O => W_18_31_i_3_n_0
);
W_18_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x117_out_12,
   I1 => x117_out_14,
   I2 => W_18_31_i_13_n_0,
   I3 => W_18_31_i_14_n_0,
   O => W_18_31_i_4_n_0
);
W_18_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_18_31_i_15_n_0,
   I1 => SIGMA_LCASE_1371_out_30,
   I2 => W_18_31_i_17_n_0,
   I3 => M_reg_11_30,
   I4 => SIGMA_LCASE_0367_out_30,
   I5 => M_reg_2_30,
   O => W_18_31_i_5_n_0
);
W_18_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_18_31_i_2_n_0,
   I1 => W_18_31_i_19_n_0,
   I2 => x117_out_15,
   I3 => x117_out_17,
   I4 => W_18_31_i_15_n_0,
   O => W_18_31_i_6_n_0
);
W_18_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x117_out_14,
   I1 => x117_out_16,
   I2 => W_18_31_i_9_n_0,
   I3 => W_18_31_i_10_n_0,
   I4 => W_18_31_i_3_n_0,
   O => W_18_31_i_7_n_0
);
W_18_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x117_out_13,
   I1 => x117_out_15,
   I2 => W_18_31_i_11_n_0,
   I3 => W_18_31_i_12_n_0,
   I4 => W_18_31_i_4_n_0,
   O => W_18_31_i_8_n_0
);
W_18_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => M_reg_2_29,
   I1 => M_reg_11_29,
   I2 => M_reg_3_15,
   I3 => M_reg_3_4,
   O => W_18_31_i_9_n_0
);
W_18_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_2_2,
   I1 => M_reg_11_2,
   I2 => M_reg_3_20,
   I3 => M_reg_3_9,
   I4 => M_reg_3_5,
   O => W_18_3_i_10_n_0
);
W_18_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_11_1,
   I1 => M_reg_3_4,
   I2 => M_reg_3_8,
   I3 => M_reg_3_19,
   I4 => M_reg_2_1,
   O => W_18_3_i_11_n_0
);
W_18_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => M_reg_3_19,
   I1 => M_reg_3_8,
   I2 => M_reg_3_4,
   O => SIGMA_LCASE_0367_out_1
);
W_18_3_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_2_1,
   I1 => M_reg_11_1,
   I2 => M_reg_3_19,
   I3 => M_reg_3_8,
   I4 => M_reg_3_4,
   O => W_18_3_i_13_n_0
);
W_18_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x117_out_12,
   I1 => x117_out_19,
   I2 => x117_out_21,
   I3 => W_18_3_i_10_n_0,
   I4 => W_18_3_i_11_n_0,
   O => W_18_3_i_2_n_0
);
W_18_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_18_3_i_11_n_0,
   I1 => x117_out_21,
   I2 => x117_out_19,
   I3 => x117_out_12,
   I4 => W_18_3_i_10_n_0,
   O => W_18_3_i_3_n_0
);
W_18_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_0367_out_1,
   I1 => M_reg_11_1,
   I2 => M_reg_2_1,
   I3 => x117_out_11,
   I4 => x117_out_18,
   I5 => x117_out_20,
   O => W_18_3_i_4_n_0
);
W_18_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_2_0,
   I1 => M_reg_11_0,
   I2 => M_reg_3_18,
   I3 => M_reg_3_7,
   I4 => M_reg_3_3,
   O => W_18_3_i_5_n_0
);
W_18_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_18_3_i_2_n_0,
   I1 => W_18_7_i_16_n_0,
   I2 => x117_out_13,
   I3 => x117_out_20,
   I4 => x117_out_22,
   I5 => W_18_7_i_17_n_0,
   O => W_18_3_i_6_n_0
);
W_18_3_i_7 : LUT5
  generic map(
   INIT => X"6aa6a66a"
  )
 port map (
   I0 => W_18_3_i_3_n_0,
   I1 => W_18_3_i_13_n_0,
   I2 => x117_out_20,
   I3 => x117_out_18,
   I4 => x117_out_11,
   O => W_18_3_i_7_n_0
);
W_18_3_i_8 : LUT6
  generic map(
   INIT => X"566565566aa6a66a"
  )
 port map (
   I0 => W_18_3_i_4_n_0,
   I1 => M_reg_2_0,
   I2 => M_reg_3_18,
   I3 => M_reg_3_7,
   I4 => M_reg_3_3,
   I5 => M_reg_11_0,
   O => W_18_3_i_8_n_0
);
W_18_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_18_3_i_5_n_0,
   I1 => x117_out_10,
   I2 => x117_out_17,
   I3 => x117_out_19,
   O => W_18_3_i_9_n_0
);
W_18_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_2_6,
   I1 => M_reg_11_6,
   I2 => M_reg_3_24,
   I3 => M_reg_3_13,
   I4 => M_reg_3_9,
   O => W_18_7_i_10_n_0
);
W_18_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_11_5,
   I1 => M_reg_3_8,
   I2 => M_reg_3_12,
   I3 => M_reg_3_23,
   I4 => M_reg_2_5,
   O => W_18_7_i_11_n_0
);
W_18_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_2_5,
   I1 => M_reg_11_5,
   I2 => M_reg_3_23,
   I3 => M_reg_3_12,
   I4 => M_reg_3_8,
   O => W_18_7_i_12_n_0
);
W_18_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_11_4,
   I1 => M_reg_3_7,
   I2 => M_reg_3_11,
   I3 => M_reg_3_22,
   I4 => M_reg_2_4,
   O => W_18_7_i_13_n_0
);
W_18_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_2_4,
   I1 => M_reg_11_4,
   I2 => M_reg_3_22,
   I3 => M_reg_3_11,
   I4 => M_reg_3_7,
   O => W_18_7_i_14_n_0
);
W_18_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_11_3,
   I1 => M_reg_3_6,
   I2 => M_reg_3_10,
   I3 => M_reg_3_21,
   I4 => M_reg_2_3,
   O => W_18_7_i_15_n_0
);
W_18_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_2_3,
   I1 => M_reg_11_3,
   I2 => M_reg_3_21,
   I3 => M_reg_3_10,
   I4 => M_reg_3_6,
   O => W_18_7_i_16_n_0
);
W_18_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_11_2,
   I1 => M_reg_3_5,
   I2 => M_reg_3_9,
   I3 => M_reg_3_20,
   I4 => M_reg_2_2,
   O => W_18_7_i_17_n_0
);
W_18_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x117_out_16,
   I1 => x117_out_23,
   I2 => x117_out_25,
   I3 => W_18_7_i_10_n_0,
   I4 => W_18_7_i_11_n_0,
   O => W_18_7_i_2_n_0
);
W_18_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x117_out_15,
   I1 => x117_out_22,
   I2 => x117_out_24,
   I3 => W_18_7_i_12_n_0,
   I4 => W_18_7_i_13_n_0,
   O => W_18_7_i_3_n_0
);
W_18_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x117_out_14,
   I1 => x117_out_21,
   I2 => x117_out_23,
   I3 => W_18_7_i_14_n_0,
   I4 => W_18_7_i_15_n_0,
   O => W_18_7_i_4_n_0
);
W_18_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x117_out_13,
   I1 => x117_out_20,
   I2 => x117_out_22,
   I3 => W_18_7_i_16_n_0,
   I4 => W_18_7_i_17_n_0,
   O => W_18_7_i_5_n_0
);
W_18_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_18_7_i_2_n_0,
   I1 => W_18_11_i_16_n_0,
   I2 => x117_out_17,
   I3 => x117_out_24,
   I4 => x117_out_26,
   I5 => W_18_11_i_17_n_0,
   O => W_18_7_i_6_n_0
);
W_18_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_18_7_i_3_n_0,
   I1 => W_18_7_i_10_n_0,
   I2 => x117_out_16,
   I3 => x117_out_23,
   I4 => x117_out_25,
   I5 => W_18_7_i_11_n_0,
   O => W_18_7_i_7_n_0
);
W_18_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_18_7_i_4_n_0,
   I1 => W_18_7_i_12_n_0,
   I2 => x117_out_15,
   I3 => x117_out_22,
   I4 => x117_out_24,
   I5 => W_18_7_i_13_n_0,
   O => W_18_7_i_8_n_0
);
W_18_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_18_7_i_5_n_0,
   I1 => W_18_7_i_14_n_0,
   I2 => x117_out_14,
   I3 => x117_out_21,
   I4 => x117_out_23,
   I5 => W_18_7_i_15_n_0,
   O => W_18_7_i_9_n_0
);
W_19_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_3_10,
   I1 => M_reg_12_10,
   I2 => M_reg_4_28,
   I3 => M_reg_4_17,
   I4 => M_reg_4_13,
   O => W_19_11_i_10_n_0
);
W_19_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_12_9,
   I1 => M_reg_4_12,
   I2 => M_reg_4_16,
   I3 => M_reg_4_27,
   I4 => M_reg_3_9,
   O => W_19_11_i_11_n_0
);
W_19_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_3_9,
   I1 => M_reg_12_9,
   I2 => M_reg_4_27,
   I3 => M_reg_4_16,
   I4 => M_reg_4_12,
   O => W_19_11_i_12_n_0
);
W_19_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_12_8,
   I1 => M_reg_4_11,
   I2 => M_reg_4_15,
   I3 => M_reg_4_26,
   I4 => M_reg_3_8,
   O => W_19_11_i_13_n_0
);
W_19_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_3_8,
   I1 => M_reg_12_8,
   I2 => M_reg_4_26,
   I3 => M_reg_4_15,
   I4 => M_reg_4_11,
   O => W_19_11_i_14_n_0
);
W_19_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_12_7,
   I1 => M_reg_4_10,
   I2 => M_reg_4_14,
   I3 => M_reg_4_25,
   I4 => M_reg_3_7,
   O => W_19_11_i_15_n_0
);
W_19_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_3_7,
   I1 => M_reg_12_7,
   I2 => M_reg_4_25,
   I3 => M_reg_4_14,
   I4 => M_reg_4_10,
   O => W_19_11_i_16_n_0
);
W_19_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_12_6,
   I1 => M_reg_4_9,
   I2 => M_reg_4_13,
   I3 => M_reg_4_24,
   I4 => M_reg_3_6,
   O => W_19_11_i_17_n_0
);
W_19_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x116_out_20,
   I1 => x116_out_27,
   I2 => x116_out_29,
   I3 => W_19_11_i_10_n_0,
   I4 => W_19_11_i_11_n_0,
   O => W_19_11_i_2_n_0
);
W_19_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x116_out_19,
   I1 => x116_out_26,
   I2 => x116_out_28,
   I3 => W_19_11_i_12_n_0,
   I4 => W_19_11_i_13_n_0,
   O => W_19_11_i_3_n_0
);
W_19_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x116_out_18,
   I1 => x116_out_25,
   I2 => x116_out_27,
   I3 => W_19_11_i_14_n_0,
   I4 => W_19_11_i_15_n_0,
   O => W_19_11_i_4_n_0
);
W_19_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x116_out_17,
   I1 => x116_out_24,
   I2 => x116_out_26,
   I3 => W_19_11_i_16_n_0,
   I4 => W_19_11_i_17_n_0,
   O => W_19_11_i_5_n_0
);
W_19_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_19_11_i_2_n_0,
   I1 => W_19_15_i_16_n_0,
   I2 => x116_out_21,
   I3 => x116_out_28,
   I4 => x116_out_30,
   I5 => W_19_15_i_17_n_0,
   O => W_19_11_i_6_n_0
);
W_19_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_19_11_i_3_n_0,
   I1 => W_19_11_i_10_n_0,
   I2 => x116_out_20,
   I3 => x116_out_27,
   I4 => x116_out_29,
   I5 => W_19_11_i_11_n_0,
   O => W_19_11_i_7_n_0
);
W_19_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_19_11_i_4_n_0,
   I1 => W_19_11_i_12_n_0,
   I2 => x116_out_19,
   I3 => x116_out_26,
   I4 => x116_out_28,
   I5 => W_19_11_i_13_n_0,
   O => W_19_11_i_8_n_0
);
W_19_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_19_11_i_5_n_0,
   I1 => W_19_11_i_14_n_0,
   I2 => x116_out_18,
   I3 => x116_out_25,
   I4 => x116_out_27,
   I5 => W_19_11_i_15_n_0,
   O => W_19_11_i_9_n_0
);
W_19_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_3_14,
   I1 => M_reg_12_14,
   I2 => M_reg_4_0,
   I3 => M_reg_4_21,
   I4 => M_reg_4_17,
   O => W_19_15_i_10_n_0
);
W_19_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_12_13,
   I1 => M_reg_4_16,
   I2 => M_reg_4_20,
   I3 => M_reg_4_31,
   I4 => M_reg_3_13,
   O => W_19_15_i_11_n_0
);
W_19_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_3_13,
   I1 => M_reg_12_13,
   I2 => M_reg_4_31,
   I3 => M_reg_4_20,
   I4 => M_reg_4_16,
   O => W_19_15_i_12_n_0
);
W_19_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_12_12,
   I1 => M_reg_4_15,
   I2 => M_reg_4_19,
   I3 => M_reg_4_30,
   I4 => M_reg_3_12,
   O => W_19_15_i_13_n_0
);
W_19_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_3_12,
   I1 => M_reg_12_12,
   I2 => M_reg_4_30,
   I3 => M_reg_4_19,
   I4 => M_reg_4_15,
   O => W_19_15_i_14_n_0
);
W_19_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_12_11,
   I1 => M_reg_4_14,
   I2 => M_reg_4_18,
   I3 => M_reg_4_29,
   I4 => M_reg_3_11,
   O => W_19_15_i_15_n_0
);
W_19_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_3_11,
   I1 => M_reg_12_11,
   I2 => M_reg_4_29,
   I3 => M_reg_4_18,
   I4 => M_reg_4_14,
   O => W_19_15_i_16_n_0
);
W_19_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_12_10,
   I1 => M_reg_4_13,
   I2 => M_reg_4_17,
   I3 => M_reg_4_28,
   I4 => M_reg_3_10,
   O => W_19_15_i_17_n_0
);
W_19_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x116_out_24,
   I1 => x116_out_31,
   I2 => x116_out_1,
   I3 => W_19_15_i_10_n_0,
   I4 => W_19_15_i_11_n_0,
   O => W_19_15_i_2_n_0
);
W_19_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x116_out_23,
   I1 => x116_out_30,
   I2 => x116_out_0,
   I3 => W_19_15_i_12_n_0,
   I4 => W_19_15_i_13_n_0,
   O => W_19_15_i_3_n_0
);
W_19_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x116_out_22,
   I1 => x116_out_29,
   I2 => x116_out_31,
   I3 => W_19_15_i_14_n_0,
   I4 => W_19_15_i_15_n_0,
   O => W_19_15_i_4_n_0
);
W_19_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x116_out_21,
   I1 => x116_out_28,
   I2 => x116_out_30,
   I3 => W_19_15_i_16_n_0,
   I4 => W_19_15_i_17_n_0,
   O => W_19_15_i_5_n_0
);
W_19_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_19_15_i_2_n_0,
   I1 => W_19_19_i_16_n_0,
   I2 => x116_out_25,
   I3 => x116_out_0,
   I4 => x116_out_2,
   I5 => W_19_19_i_17_n_0,
   O => W_19_15_i_6_n_0
);
W_19_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_19_15_i_3_n_0,
   I1 => W_19_15_i_10_n_0,
   I2 => x116_out_24,
   I3 => x116_out_31,
   I4 => x116_out_1,
   I5 => W_19_15_i_11_n_0,
   O => W_19_15_i_7_n_0
);
W_19_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_19_15_i_4_n_0,
   I1 => W_19_15_i_12_n_0,
   I2 => x116_out_23,
   I3 => x116_out_30,
   I4 => x116_out_0,
   I5 => W_19_15_i_13_n_0,
   O => W_19_15_i_8_n_0
);
W_19_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_19_15_i_5_n_0,
   I1 => W_19_15_i_14_n_0,
   I2 => x116_out_22,
   I3 => x116_out_29,
   I4 => x116_out_31,
   I5 => W_19_15_i_15_n_0,
   O => W_19_15_i_9_n_0
);
W_19_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_3_18,
   I1 => M_reg_12_18,
   I2 => M_reg_4_4,
   I3 => M_reg_4_25,
   I4 => M_reg_4_21,
   O => W_19_19_i_10_n_0
);
W_19_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_12_17,
   I1 => M_reg_4_20,
   I2 => M_reg_4_24,
   I3 => M_reg_4_3,
   I4 => M_reg_3_17,
   O => W_19_19_i_11_n_0
);
W_19_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_3_17,
   I1 => M_reg_12_17,
   I2 => M_reg_4_3,
   I3 => M_reg_4_24,
   I4 => M_reg_4_20,
   O => W_19_19_i_12_n_0
);
W_19_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_12_16,
   I1 => M_reg_4_19,
   I2 => M_reg_4_23,
   I3 => M_reg_4_2,
   I4 => M_reg_3_16,
   O => W_19_19_i_13_n_0
);
W_19_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_3_16,
   I1 => M_reg_12_16,
   I2 => M_reg_4_2,
   I3 => M_reg_4_23,
   I4 => M_reg_4_19,
   O => W_19_19_i_14_n_0
);
W_19_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_12_15,
   I1 => M_reg_4_18,
   I2 => M_reg_4_22,
   I3 => M_reg_4_1,
   I4 => M_reg_3_15,
   O => W_19_19_i_15_n_0
);
W_19_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_3_15,
   I1 => M_reg_12_15,
   I2 => M_reg_4_1,
   I3 => M_reg_4_22,
   I4 => M_reg_4_18,
   O => W_19_19_i_16_n_0
);
W_19_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_12_14,
   I1 => M_reg_4_17,
   I2 => M_reg_4_21,
   I3 => M_reg_4_0,
   I4 => M_reg_3_14,
   O => W_19_19_i_17_n_0
);
W_19_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x116_out_28,
   I1 => x116_out_3,
   I2 => x116_out_5,
   I3 => W_19_19_i_10_n_0,
   I4 => W_19_19_i_11_n_0,
   O => W_19_19_i_2_n_0
);
W_19_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x116_out_27,
   I1 => x116_out_2,
   I2 => x116_out_4,
   I3 => W_19_19_i_12_n_0,
   I4 => W_19_19_i_13_n_0,
   O => W_19_19_i_3_n_0
);
W_19_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x116_out_26,
   I1 => x116_out_1,
   I2 => x116_out_3,
   I3 => W_19_19_i_14_n_0,
   I4 => W_19_19_i_15_n_0,
   O => W_19_19_i_4_n_0
);
W_19_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x116_out_25,
   I1 => x116_out_0,
   I2 => x116_out_2,
   I3 => W_19_19_i_16_n_0,
   I4 => W_19_19_i_17_n_0,
   O => W_19_19_i_5_n_0
);
W_19_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_19_19_i_2_n_0,
   I1 => W_19_23_i_16_n_0,
   I2 => x116_out_29,
   I3 => x116_out_4,
   I4 => x116_out_6,
   I5 => W_19_23_i_17_n_0,
   O => W_19_19_i_6_n_0
);
W_19_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_19_19_i_3_n_0,
   I1 => W_19_19_i_10_n_0,
   I2 => x116_out_28,
   I3 => x116_out_3,
   I4 => x116_out_5,
   I5 => W_19_19_i_11_n_0,
   O => W_19_19_i_7_n_0
);
W_19_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_19_19_i_4_n_0,
   I1 => W_19_19_i_12_n_0,
   I2 => x116_out_27,
   I3 => x116_out_2,
   I4 => x116_out_4,
   I5 => W_19_19_i_13_n_0,
   O => W_19_19_i_8_n_0
);
W_19_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_19_19_i_5_n_0,
   I1 => W_19_19_i_14_n_0,
   I2 => x116_out_26,
   I3 => x116_out_1,
   I4 => x116_out_3,
   I5 => W_19_19_i_15_n_0,
   O => W_19_19_i_9_n_0
);
W_19_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_3_22,
   I1 => M_reg_12_22,
   I2 => M_reg_4_8,
   I3 => M_reg_4_29,
   I4 => M_reg_4_25,
   O => W_19_23_i_10_n_0
);
W_19_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_12_21,
   I1 => M_reg_4_24,
   I2 => M_reg_4_28,
   I3 => M_reg_4_7,
   I4 => M_reg_3_21,
   O => W_19_23_i_11_n_0
);
W_19_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_3_21,
   I1 => M_reg_12_21,
   I2 => M_reg_4_7,
   I3 => M_reg_4_28,
   I4 => M_reg_4_24,
   O => W_19_23_i_12_n_0
);
W_19_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_12_20,
   I1 => M_reg_4_23,
   I2 => M_reg_4_27,
   I3 => M_reg_4_6,
   I4 => M_reg_3_20,
   O => W_19_23_i_13_n_0
);
W_19_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_3_20,
   I1 => M_reg_12_20,
   I2 => M_reg_4_6,
   I3 => M_reg_4_27,
   I4 => M_reg_4_23,
   O => W_19_23_i_14_n_0
);
W_19_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_12_19,
   I1 => M_reg_4_22,
   I2 => M_reg_4_26,
   I3 => M_reg_4_5,
   I4 => M_reg_3_19,
   O => W_19_23_i_15_n_0
);
W_19_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_3_19,
   I1 => M_reg_12_19,
   I2 => M_reg_4_5,
   I3 => M_reg_4_26,
   I4 => M_reg_4_22,
   O => W_19_23_i_16_n_0
);
W_19_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_12_18,
   I1 => M_reg_4_21,
   I2 => M_reg_4_25,
   I3 => M_reg_4_4,
   I4 => M_reg_3_18,
   O => W_19_23_i_17_n_0
);
W_19_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x116_out_7,
   I1 => x116_out_9,
   I2 => W_19_23_i_10_n_0,
   I3 => W_19_23_i_11_n_0,
   O => W_19_23_i_2_n_0
);
W_19_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x116_out_31,
   I1 => x116_out_6,
   I2 => x116_out_8,
   I3 => W_19_23_i_12_n_0,
   I4 => W_19_23_i_13_n_0,
   O => W_19_23_i_3_n_0
);
W_19_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x116_out_30,
   I1 => x116_out_5,
   I2 => x116_out_7,
   I3 => W_19_23_i_14_n_0,
   I4 => W_19_23_i_15_n_0,
   O => W_19_23_i_4_n_0
);
W_19_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x116_out_29,
   I1 => x116_out_4,
   I2 => x116_out_6,
   I3 => W_19_23_i_16_n_0,
   I4 => W_19_23_i_17_n_0,
   O => W_19_23_i_5_n_0
);
W_19_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x116_out_8,
   I1 => x116_out_10,
   I2 => W_19_27_i_16_n_0,
   I3 => W_19_27_i_17_n_0,
   I4 => W_19_23_i_2_n_0,
   O => W_19_23_i_6_n_0
);
W_19_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x116_out_7,
   I1 => x116_out_9,
   I2 => W_19_23_i_10_n_0,
   I3 => W_19_23_i_11_n_0,
   I4 => W_19_23_i_3_n_0,
   O => W_19_23_i_7_n_0
);
W_19_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_19_23_i_4_n_0,
   I1 => W_19_23_i_12_n_0,
   I2 => x116_out_31,
   I3 => x116_out_6,
   I4 => x116_out_8,
   I5 => W_19_23_i_13_n_0,
   O => W_19_23_i_8_n_0
);
W_19_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_19_23_i_5_n_0,
   I1 => W_19_23_i_14_n_0,
   I2 => x116_out_30,
   I3 => x116_out_5,
   I4 => x116_out_7,
   I5 => W_19_23_i_15_n_0,
   O => W_19_23_i_9_n_0
);
W_19_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_3_26,
   I1 => M_reg_12_26,
   I2 => M_reg_4_12,
   I3 => M_reg_4_1,
   I4 => M_reg_4_29,
   O => W_19_27_i_10_n_0
);
W_19_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_12_25,
   I1 => M_reg_4_28,
   I2 => M_reg_4_0,
   I3 => M_reg_4_11,
   I4 => M_reg_3_25,
   O => W_19_27_i_11_n_0
);
W_19_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_3_25,
   I1 => M_reg_12_25,
   I2 => M_reg_4_11,
   I3 => M_reg_4_0,
   I4 => M_reg_4_28,
   O => W_19_27_i_12_n_0
);
W_19_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_12_24,
   I1 => M_reg_4_27,
   I2 => M_reg_4_31,
   I3 => M_reg_4_10,
   I4 => M_reg_3_24,
   O => W_19_27_i_13_n_0
);
W_19_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_3_24,
   I1 => M_reg_12_24,
   I2 => M_reg_4_10,
   I3 => M_reg_4_31,
   I4 => M_reg_4_27,
   O => W_19_27_i_14_n_0
);
W_19_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_12_23,
   I1 => M_reg_4_26,
   I2 => M_reg_4_30,
   I3 => M_reg_4_9,
   I4 => M_reg_3_23,
   O => W_19_27_i_15_n_0
);
W_19_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_3_23,
   I1 => M_reg_12_23,
   I2 => M_reg_4_9,
   I3 => M_reg_4_30,
   I4 => M_reg_4_26,
   O => W_19_27_i_16_n_0
);
W_19_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_12_22,
   I1 => M_reg_4_25,
   I2 => M_reg_4_29,
   I3 => M_reg_4_8,
   I4 => M_reg_3_22,
   O => W_19_27_i_17_n_0
);
W_19_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x116_out_11,
   I1 => x116_out_13,
   I2 => W_19_27_i_10_n_0,
   I3 => W_19_27_i_11_n_0,
   O => W_19_27_i_2_n_0
);
W_19_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x116_out_10,
   I1 => x116_out_12,
   I2 => W_19_27_i_12_n_0,
   I3 => W_19_27_i_13_n_0,
   O => W_19_27_i_3_n_0
);
W_19_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x116_out_9,
   I1 => x116_out_11,
   I2 => W_19_27_i_14_n_0,
   I3 => W_19_27_i_15_n_0,
   O => W_19_27_i_4_n_0
);
W_19_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x116_out_8,
   I1 => x116_out_10,
   I2 => W_19_27_i_16_n_0,
   I3 => W_19_27_i_17_n_0,
   O => W_19_27_i_5_n_0
);
W_19_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x116_out_12,
   I1 => x116_out_14,
   I2 => W_19_31_i_13_n_0,
   I3 => W_19_31_i_14_n_0,
   I4 => W_19_27_i_2_n_0,
   O => W_19_27_i_6_n_0
);
W_19_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x116_out_11,
   I1 => x116_out_13,
   I2 => W_19_27_i_10_n_0,
   I3 => W_19_27_i_11_n_0,
   I4 => W_19_27_i_3_n_0,
   O => W_19_27_i_7_n_0
);
W_19_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x116_out_10,
   I1 => x116_out_12,
   I2 => W_19_27_i_12_n_0,
   I3 => W_19_27_i_13_n_0,
   I4 => W_19_27_i_4_n_0,
   O => W_19_27_i_8_n_0
);
W_19_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x116_out_9,
   I1 => x116_out_11,
   I2 => W_19_27_i_14_n_0,
   I3 => W_19_27_i_15_n_0,
   I4 => W_19_27_i_5_n_0,
   O => W_19_27_i_9_n_0
);
W_19_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_12_28,
   I1 => M_reg_4_31,
   I2 => M_reg_4_3,
   I3 => M_reg_4_14,
   I4 => M_reg_3_28,
   O => W_19_31_i_10_n_0
);
W_19_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_3_28,
   I1 => M_reg_12_28,
   I2 => M_reg_4_14,
   I3 => M_reg_4_3,
   I4 => M_reg_4_31,
   O => W_19_31_i_11_n_0
);
W_19_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_12_27,
   I1 => M_reg_4_30,
   I2 => M_reg_4_2,
   I3 => M_reg_4_13,
   I4 => M_reg_3_27,
   O => W_19_31_i_12_n_0
);
W_19_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_3_27,
   I1 => M_reg_12_27,
   I2 => M_reg_4_13,
   I3 => M_reg_4_2,
   I4 => M_reg_4_30,
   O => W_19_31_i_13_n_0
);
W_19_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_12_26,
   I1 => M_reg_4_29,
   I2 => M_reg_4_1,
   I3 => M_reg_4_12,
   I4 => M_reg_3_26,
   O => W_19_31_i_14_n_0
);
W_19_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => M_reg_12_29,
   I1 => M_reg_4_4,
   I2 => M_reg_4_15,
   I3 => M_reg_3_29,
   O => W_19_31_i_15_n_0
);
W_19_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x116_out_17,
   I1 => x116_out_15,
   O => SIGMA_LCASE_1363_out_30
);
W_19_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => M_reg_4_6,
   I1 => M_reg_4_17,
   I2 => M_reg_12_31,
   I3 => M_reg_3_31,
   I4 => x116_out_16,
   I5 => x116_out_18,
   O => W_19_31_i_17_n_0
);
W_19_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => M_reg_4_16,
   I1 => M_reg_4_5,
   O => SIGMA_LCASE_0359_out_30
);
W_19_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => M_reg_3_30,
   I1 => M_reg_12_30,
   I2 => M_reg_4_16,
   I3 => M_reg_4_5,
   O => W_19_31_i_19_n_0
);
W_19_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x116_out_14,
   I1 => x116_out_16,
   I2 => W_19_31_i_9_n_0,
   I3 => W_19_31_i_10_n_0,
   O => W_19_31_i_2_n_0
);
W_19_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x116_out_13,
   I1 => x116_out_15,
   I2 => W_19_31_i_11_n_0,
   I3 => W_19_31_i_12_n_0,
   O => W_19_31_i_3_n_0
);
W_19_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x116_out_12,
   I1 => x116_out_14,
   I2 => W_19_31_i_13_n_0,
   I3 => W_19_31_i_14_n_0,
   O => W_19_31_i_4_n_0
);
W_19_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_19_31_i_15_n_0,
   I1 => SIGMA_LCASE_1363_out_30,
   I2 => W_19_31_i_17_n_0,
   I3 => M_reg_12_30,
   I4 => SIGMA_LCASE_0359_out_30,
   I5 => M_reg_3_30,
   O => W_19_31_i_5_n_0
);
W_19_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_19_31_i_2_n_0,
   I1 => W_19_31_i_19_n_0,
   I2 => x116_out_15,
   I3 => x116_out_17,
   I4 => W_19_31_i_15_n_0,
   O => W_19_31_i_6_n_0
);
W_19_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x116_out_14,
   I1 => x116_out_16,
   I2 => W_19_31_i_9_n_0,
   I3 => W_19_31_i_10_n_0,
   I4 => W_19_31_i_3_n_0,
   O => W_19_31_i_7_n_0
);
W_19_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x116_out_13,
   I1 => x116_out_15,
   I2 => W_19_31_i_11_n_0,
   I3 => W_19_31_i_12_n_0,
   I4 => W_19_31_i_4_n_0,
   O => W_19_31_i_8_n_0
);
W_19_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => M_reg_3_29,
   I1 => M_reg_12_29,
   I2 => M_reg_4_15,
   I3 => M_reg_4_4,
   O => W_19_31_i_9_n_0
);
W_19_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_3_2,
   I1 => M_reg_12_2,
   I2 => M_reg_4_20,
   I3 => M_reg_4_9,
   I4 => M_reg_4_5,
   O => W_19_3_i_10_n_0
);
W_19_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_12_1,
   I1 => M_reg_4_4,
   I2 => M_reg_4_8,
   I3 => M_reg_4_19,
   I4 => M_reg_3_1,
   O => W_19_3_i_11_n_0
);
W_19_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => M_reg_4_19,
   I1 => M_reg_4_8,
   I2 => M_reg_4_4,
   O => SIGMA_LCASE_0359_out_1
);
W_19_3_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_3_1,
   I1 => M_reg_12_1,
   I2 => M_reg_4_19,
   I3 => M_reg_4_8,
   I4 => M_reg_4_4,
   O => W_19_3_i_13_n_0
);
W_19_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x116_out_12,
   I1 => x116_out_19,
   I2 => x116_out_21,
   I3 => W_19_3_i_10_n_0,
   I4 => W_19_3_i_11_n_0,
   O => W_19_3_i_2_n_0
);
W_19_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_19_3_i_11_n_0,
   I1 => x116_out_21,
   I2 => x116_out_19,
   I3 => x116_out_12,
   I4 => W_19_3_i_10_n_0,
   O => W_19_3_i_3_n_0
);
W_19_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_0359_out_1,
   I1 => M_reg_12_1,
   I2 => M_reg_3_1,
   I3 => x116_out_11,
   I4 => x116_out_18,
   I5 => x116_out_20,
   O => W_19_3_i_4_n_0
);
W_19_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_3_0,
   I1 => M_reg_12_0,
   I2 => M_reg_4_18,
   I3 => M_reg_4_7,
   I4 => M_reg_4_3,
   O => W_19_3_i_5_n_0
);
W_19_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_19_3_i_2_n_0,
   I1 => W_19_7_i_16_n_0,
   I2 => x116_out_13,
   I3 => x116_out_20,
   I4 => x116_out_22,
   I5 => W_19_7_i_17_n_0,
   O => W_19_3_i_6_n_0
);
W_19_3_i_7 : LUT5
  generic map(
   INIT => X"6aa6a66a"
  )
 port map (
   I0 => W_19_3_i_3_n_0,
   I1 => W_19_3_i_13_n_0,
   I2 => x116_out_20,
   I3 => x116_out_18,
   I4 => x116_out_11,
   O => W_19_3_i_7_n_0
);
W_19_3_i_8 : LUT6
  generic map(
   INIT => X"566565566aa6a66a"
  )
 port map (
   I0 => W_19_3_i_4_n_0,
   I1 => M_reg_3_0,
   I2 => M_reg_4_18,
   I3 => M_reg_4_7,
   I4 => M_reg_4_3,
   I5 => M_reg_12_0,
   O => W_19_3_i_8_n_0
);
W_19_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_19_3_i_5_n_0,
   I1 => x116_out_10,
   I2 => x116_out_17,
   I3 => x116_out_19,
   O => W_19_3_i_9_n_0
);
W_19_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_3_6,
   I1 => M_reg_12_6,
   I2 => M_reg_4_24,
   I3 => M_reg_4_13,
   I4 => M_reg_4_9,
   O => W_19_7_i_10_n_0
);
W_19_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_12_5,
   I1 => M_reg_4_8,
   I2 => M_reg_4_12,
   I3 => M_reg_4_23,
   I4 => M_reg_3_5,
   O => W_19_7_i_11_n_0
);
W_19_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_3_5,
   I1 => M_reg_12_5,
   I2 => M_reg_4_23,
   I3 => M_reg_4_12,
   I4 => M_reg_4_8,
   O => W_19_7_i_12_n_0
);
W_19_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_12_4,
   I1 => M_reg_4_7,
   I2 => M_reg_4_11,
   I3 => M_reg_4_22,
   I4 => M_reg_3_4,
   O => W_19_7_i_13_n_0
);
W_19_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_3_4,
   I1 => M_reg_12_4,
   I2 => M_reg_4_22,
   I3 => M_reg_4_11,
   I4 => M_reg_4_7,
   O => W_19_7_i_14_n_0
);
W_19_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_12_3,
   I1 => M_reg_4_6,
   I2 => M_reg_4_10,
   I3 => M_reg_4_21,
   I4 => M_reg_3_3,
   O => W_19_7_i_15_n_0
);
W_19_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_3_3,
   I1 => M_reg_12_3,
   I2 => M_reg_4_21,
   I3 => M_reg_4_10,
   I4 => M_reg_4_6,
   O => W_19_7_i_16_n_0
);
W_19_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_12_2,
   I1 => M_reg_4_5,
   I2 => M_reg_4_9,
   I3 => M_reg_4_20,
   I4 => M_reg_3_2,
   O => W_19_7_i_17_n_0
);
W_19_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x116_out_16,
   I1 => x116_out_23,
   I2 => x116_out_25,
   I3 => W_19_7_i_10_n_0,
   I4 => W_19_7_i_11_n_0,
   O => W_19_7_i_2_n_0
);
W_19_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x116_out_15,
   I1 => x116_out_22,
   I2 => x116_out_24,
   I3 => W_19_7_i_12_n_0,
   I4 => W_19_7_i_13_n_0,
   O => W_19_7_i_3_n_0
);
W_19_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x116_out_14,
   I1 => x116_out_21,
   I2 => x116_out_23,
   I3 => W_19_7_i_14_n_0,
   I4 => W_19_7_i_15_n_0,
   O => W_19_7_i_4_n_0
);
W_19_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x116_out_13,
   I1 => x116_out_20,
   I2 => x116_out_22,
   I3 => W_19_7_i_16_n_0,
   I4 => W_19_7_i_17_n_0,
   O => W_19_7_i_5_n_0
);
W_19_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_19_7_i_2_n_0,
   I1 => W_19_11_i_16_n_0,
   I2 => x116_out_17,
   I3 => x116_out_24,
   I4 => x116_out_26,
   I5 => W_19_11_i_17_n_0,
   O => W_19_7_i_6_n_0
);
W_19_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_19_7_i_3_n_0,
   I1 => W_19_7_i_10_n_0,
   I2 => x116_out_16,
   I3 => x116_out_23,
   I4 => x116_out_25,
   I5 => W_19_7_i_11_n_0,
   O => W_19_7_i_7_n_0
);
W_19_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_19_7_i_4_n_0,
   I1 => W_19_7_i_12_n_0,
   I2 => x116_out_15,
   I3 => x116_out_22,
   I4 => x116_out_24,
   I5 => W_19_7_i_13_n_0,
   O => W_19_7_i_8_n_0
);
W_19_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_19_7_i_5_n_0,
   I1 => W_19_7_i_14_n_0,
   I2 => x116_out_14,
   I3 => x116_out_21,
   I4 => x116_out_23,
   I5 => W_19_7_i_15_n_0,
   O => W_19_7_i_9_n_0
);
W_20_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_4_10,
   I1 => M_reg_13_10,
   I2 => M_reg_5_28,
   I3 => M_reg_5_17,
   I4 => M_reg_5_13,
   O => W_20_11_i_10_n_0
);
W_20_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_13_9,
   I1 => M_reg_5_12,
   I2 => M_reg_5_16,
   I3 => M_reg_5_27,
   I4 => M_reg_4_9,
   O => W_20_11_i_11_n_0
);
W_20_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_4_9,
   I1 => M_reg_13_9,
   I2 => M_reg_5_27,
   I3 => M_reg_5_16,
   I4 => M_reg_5_12,
   O => W_20_11_i_12_n_0
);
W_20_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_13_8,
   I1 => M_reg_5_11,
   I2 => M_reg_5_15,
   I3 => M_reg_5_26,
   I4 => M_reg_4_8,
   O => W_20_11_i_13_n_0
);
W_20_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_4_8,
   I1 => M_reg_13_8,
   I2 => M_reg_5_26,
   I3 => M_reg_5_15,
   I4 => M_reg_5_11,
   O => W_20_11_i_14_n_0
);
W_20_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_13_7,
   I1 => M_reg_5_10,
   I2 => M_reg_5_14,
   I3 => M_reg_5_25,
   I4 => M_reg_4_7,
   O => W_20_11_i_15_n_0
);
W_20_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_4_7,
   I1 => M_reg_13_7,
   I2 => M_reg_5_25,
   I3 => M_reg_5_14,
   I4 => M_reg_5_10,
   O => W_20_11_i_16_n_0
);
W_20_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_13_6,
   I1 => M_reg_5_9,
   I2 => M_reg_5_13,
   I3 => M_reg_5_24,
   I4 => M_reg_4_6,
   O => W_20_11_i_17_n_0
);
W_20_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x115_out_20,
   I1 => x115_out_27,
   I2 => x115_out_29,
   I3 => W_20_11_i_10_n_0,
   I4 => W_20_11_i_11_n_0,
   O => W_20_11_i_2_n_0
);
W_20_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x115_out_19,
   I1 => x115_out_26,
   I2 => x115_out_28,
   I3 => W_20_11_i_12_n_0,
   I4 => W_20_11_i_13_n_0,
   O => W_20_11_i_3_n_0
);
W_20_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x115_out_18,
   I1 => x115_out_25,
   I2 => x115_out_27,
   I3 => W_20_11_i_14_n_0,
   I4 => W_20_11_i_15_n_0,
   O => W_20_11_i_4_n_0
);
W_20_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x115_out_17,
   I1 => x115_out_24,
   I2 => x115_out_26,
   I3 => W_20_11_i_16_n_0,
   I4 => W_20_11_i_17_n_0,
   O => W_20_11_i_5_n_0
);
W_20_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_20_11_i_2_n_0,
   I1 => W_20_15_i_16_n_0,
   I2 => x115_out_21,
   I3 => x115_out_28,
   I4 => x115_out_30,
   I5 => W_20_15_i_17_n_0,
   O => W_20_11_i_6_n_0
);
W_20_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_20_11_i_3_n_0,
   I1 => W_20_11_i_10_n_0,
   I2 => x115_out_20,
   I3 => x115_out_27,
   I4 => x115_out_29,
   I5 => W_20_11_i_11_n_0,
   O => W_20_11_i_7_n_0
);
W_20_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_20_11_i_4_n_0,
   I1 => W_20_11_i_12_n_0,
   I2 => x115_out_19,
   I3 => x115_out_26,
   I4 => x115_out_28,
   I5 => W_20_11_i_13_n_0,
   O => W_20_11_i_8_n_0
);
W_20_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_20_11_i_5_n_0,
   I1 => W_20_11_i_14_n_0,
   I2 => x115_out_18,
   I3 => x115_out_25,
   I4 => x115_out_27,
   I5 => W_20_11_i_15_n_0,
   O => W_20_11_i_9_n_0
);
W_20_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_4_14,
   I1 => M_reg_13_14,
   I2 => M_reg_5_0,
   I3 => M_reg_5_21,
   I4 => M_reg_5_17,
   O => W_20_15_i_10_n_0
);
W_20_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_13_13,
   I1 => M_reg_5_16,
   I2 => M_reg_5_20,
   I3 => M_reg_5_31,
   I4 => M_reg_4_13,
   O => W_20_15_i_11_n_0
);
W_20_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_4_13,
   I1 => M_reg_13_13,
   I2 => M_reg_5_31,
   I3 => M_reg_5_20,
   I4 => M_reg_5_16,
   O => W_20_15_i_12_n_0
);
W_20_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_13_12,
   I1 => M_reg_5_15,
   I2 => M_reg_5_19,
   I3 => M_reg_5_30,
   I4 => M_reg_4_12,
   O => W_20_15_i_13_n_0
);
W_20_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_4_12,
   I1 => M_reg_13_12,
   I2 => M_reg_5_30,
   I3 => M_reg_5_19,
   I4 => M_reg_5_15,
   O => W_20_15_i_14_n_0
);
W_20_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_13_11,
   I1 => M_reg_5_14,
   I2 => M_reg_5_18,
   I3 => M_reg_5_29,
   I4 => M_reg_4_11,
   O => W_20_15_i_15_n_0
);
W_20_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_4_11,
   I1 => M_reg_13_11,
   I2 => M_reg_5_29,
   I3 => M_reg_5_18,
   I4 => M_reg_5_14,
   O => W_20_15_i_16_n_0
);
W_20_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_13_10,
   I1 => M_reg_5_13,
   I2 => M_reg_5_17,
   I3 => M_reg_5_28,
   I4 => M_reg_4_10,
   O => W_20_15_i_17_n_0
);
W_20_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x115_out_24,
   I1 => x115_out_31,
   I2 => x115_out_1,
   I3 => W_20_15_i_10_n_0,
   I4 => W_20_15_i_11_n_0,
   O => W_20_15_i_2_n_0
);
W_20_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x115_out_23,
   I1 => x115_out_30,
   I2 => x115_out_0,
   I3 => W_20_15_i_12_n_0,
   I4 => W_20_15_i_13_n_0,
   O => W_20_15_i_3_n_0
);
W_20_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x115_out_22,
   I1 => x115_out_29,
   I2 => x115_out_31,
   I3 => W_20_15_i_14_n_0,
   I4 => W_20_15_i_15_n_0,
   O => W_20_15_i_4_n_0
);
W_20_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x115_out_21,
   I1 => x115_out_28,
   I2 => x115_out_30,
   I3 => W_20_15_i_16_n_0,
   I4 => W_20_15_i_17_n_0,
   O => W_20_15_i_5_n_0
);
W_20_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_20_15_i_2_n_0,
   I1 => W_20_19_i_16_n_0,
   I2 => x115_out_25,
   I3 => x115_out_0,
   I4 => x115_out_2,
   I5 => W_20_19_i_17_n_0,
   O => W_20_15_i_6_n_0
);
W_20_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_20_15_i_3_n_0,
   I1 => W_20_15_i_10_n_0,
   I2 => x115_out_24,
   I3 => x115_out_31,
   I4 => x115_out_1,
   I5 => W_20_15_i_11_n_0,
   O => W_20_15_i_7_n_0
);
W_20_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_20_15_i_4_n_0,
   I1 => W_20_15_i_12_n_0,
   I2 => x115_out_23,
   I3 => x115_out_30,
   I4 => x115_out_0,
   I5 => W_20_15_i_13_n_0,
   O => W_20_15_i_8_n_0
);
W_20_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_20_15_i_5_n_0,
   I1 => W_20_15_i_14_n_0,
   I2 => x115_out_22,
   I3 => x115_out_29,
   I4 => x115_out_31,
   I5 => W_20_15_i_15_n_0,
   O => W_20_15_i_9_n_0
);
W_20_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_4_18,
   I1 => M_reg_13_18,
   I2 => M_reg_5_4,
   I3 => M_reg_5_25,
   I4 => M_reg_5_21,
   O => W_20_19_i_10_n_0
);
W_20_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_13_17,
   I1 => M_reg_5_20,
   I2 => M_reg_5_24,
   I3 => M_reg_5_3,
   I4 => M_reg_4_17,
   O => W_20_19_i_11_n_0
);
W_20_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_4_17,
   I1 => M_reg_13_17,
   I2 => M_reg_5_3,
   I3 => M_reg_5_24,
   I4 => M_reg_5_20,
   O => W_20_19_i_12_n_0
);
W_20_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_13_16,
   I1 => M_reg_5_19,
   I2 => M_reg_5_23,
   I3 => M_reg_5_2,
   I4 => M_reg_4_16,
   O => W_20_19_i_13_n_0
);
W_20_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_4_16,
   I1 => M_reg_13_16,
   I2 => M_reg_5_2,
   I3 => M_reg_5_23,
   I4 => M_reg_5_19,
   O => W_20_19_i_14_n_0
);
W_20_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_13_15,
   I1 => M_reg_5_18,
   I2 => M_reg_5_22,
   I3 => M_reg_5_1,
   I4 => M_reg_4_15,
   O => W_20_19_i_15_n_0
);
W_20_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_4_15,
   I1 => M_reg_13_15,
   I2 => M_reg_5_1,
   I3 => M_reg_5_22,
   I4 => M_reg_5_18,
   O => W_20_19_i_16_n_0
);
W_20_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_13_14,
   I1 => M_reg_5_17,
   I2 => M_reg_5_21,
   I3 => M_reg_5_0,
   I4 => M_reg_4_14,
   O => W_20_19_i_17_n_0
);
W_20_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x115_out_28,
   I1 => x115_out_3,
   I2 => x115_out_5,
   I3 => W_20_19_i_10_n_0,
   I4 => W_20_19_i_11_n_0,
   O => W_20_19_i_2_n_0
);
W_20_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x115_out_27,
   I1 => x115_out_2,
   I2 => x115_out_4,
   I3 => W_20_19_i_12_n_0,
   I4 => W_20_19_i_13_n_0,
   O => W_20_19_i_3_n_0
);
W_20_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x115_out_26,
   I1 => x115_out_1,
   I2 => x115_out_3,
   I3 => W_20_19_i_14_n_0,
   I4 => W_20_19_i_15_n_0,
   O => W_20_19_i_4_n_0
);
W_20_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x115_out_25,
   I1 => x115_out_0,
   I2 => x115_out_2,
   I3 => W_20_19_i_16_n_0,
   I4 => W_20_19_i_17_n_0,
   O => W_20_19_i_5_n_0
);
W_20_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_20_19_i_2_n_0,
   I1 => W_20_23_i_16_n_0,
   I2 => x115_out_29,
   I3 => x115_out_4,
   I4 => x115_out_6,
   I5 => W_20_23_i_17_n_0,
   O => W_20_19_i_6_n_0
);
W_20_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_20_19_i_3_n_0,
   I1 => W_20_19_i_10_n_0,
   I2 => x115_out_28,
   I3 => x115_out_3,
   I4 => x115_out_5,
   I5 => W_20_19_i_11_n_0,
   O => W_20_19_i_7_n_0
);
W_20_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_20_19_i_4_n_0,
   I1 => W_20_19_i_12_n_0,
   I2 => x115_out_27,
   I3 => x115_out_2,
   I4 => x115_out_4,
   I5 => W_20_19_i_13_n_0,
   O => W_20_19_i_8_n_0
);
W_20_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_20_19_i_5_n_0,
   I1 => W_20_19_i_14_n_0,
   I2 => x115_out_26,
   I3 => x115_out_1,
   I4 => x115_out_3,
   I5 => W_20_19_i_15_n_0,
   O => W_20_19_i_9_n_0
);
W_20_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_4_22,
   I1 => M_reg_13_22,
   I2 => M_reg_5_8,
   I3 => M_reg_5_29,
   I4 => M_reg_5_25,
   O => W_20_23_i_10_n_0
);
W_20_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_13_21,
   I1 => M_reg_5_24,
   I2 => M_reg_5_28,
   I3 => M_reg_5_7,
   I4 => M_reg_4_21,
   O => W_20_23_i_11_n_0
);
W_20_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_4_21,
   I1 => M_reg_13_21,
   I2 => M_reg_5_7,
   I3 => M_reg_5_28,
   I4 => M_reg_5_24,
   O => W_20_23_i_12_n_0
);
W_20_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_13_20,
   I1 => M_reg_5_23,
   I2 => M_reg_5_27,
   I3 => M_reg_5_6,
   I4 => M_reg_4_20,
   O => W_20_23_i_13_n_0
);
W_20_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_4_20,
   I1 => M_reg_13_20,
   I2 => M_reg_5_6,
   I3 => M_reg_5_27,
   I4 => M_reg_5_23,
   O => W_20_23_i_14_n_0
);
W_20_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_13_19,
   I1 => M_reg_5_22,
   I2 => M_reg_5_26,
   I3 => M_reg_5_5,
   I4 => M_reg_4_19,
   O => W_20_23_i_15_n_0
);
W_20_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_4_19,
   I1 => M_reg_13_19,
   I2 => M_reg_5_5,
   I3 => M_reg_5_26,
   I4 => M_reg_5_22,
   O => W_20_23_i_16_n_0
);
W_20_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_13_18,
   I1 => M_reg_5_21,
   I2 => M_reg_5_25,
   I3 => M_reg_5_4,
   I4 => M_reg_4_18,
   O => W_20_23_i_17_n_0
);
W_20_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x115_out_7,
   I1 => x115_out_9,
   I2 => W_20_23_i_10_n_0,
   I3 => W_20_23_i_11_n_0,
   O => W_20_23_i_2_n_0
);
W_20_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x115_out_31,
   I1 => x115_out_6,
   I2 => x115_out_8,
   I3 => W_20_23_i_12_n_0,
   I4 => W_20_23_i_13_n_0,
   O => W_20_23_i_3_n_0
);
W_20_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x115_out_30,
   I1 => x115_out_5,
   I2 => x115_out_7,
   I3 => W_20_23_i_14_n_0,
   I4 => W_20_23_i_15_n_0,
   O => W_20_23_i_4_n_0
);
W_20_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x115_out_29,
   I1 => x115_out_4,
   I2 => x115_out_6,
   I3 => W_20_23_i_16_n_0,
   I4 => W_20_23_i_17_n_0,
   O => W_20_23_i_5_n_0
);
W_20_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x115_out_8,
   I1 => x115_out_10,
   I2 => W_20_27_i_16_n_0,
   I3 => W_20_27_i_17_n_0,
   I4 => W_20_23_i_2_n_0,
   O => W_20_23_i_6_n_0
);
W_20_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x115_out_7,
   I1 => x115_out_9,
   I2 => W_20_23_i_10_n_0,
   I3 => W_20_23_i_11_n_0,
   I4 => W_20_23_i_3_n_0,
   O => W_20_23_i_7_n_0
);
W_20_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_20_23_i_4_n_0,
   I1 => W_20_23_i_12_n_0,
   I2 => x115_out_31,
   I3 => x115_out_6,
   I4 => x115_out_8,
   I5 => W_20_23_i_13_n_0,
   O => W_20_23_i_8_n_0
);
W_20_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_20_23_i_5_n_0,
   I1 => W_20_23_i_14_n_0,
   I2 => x115_out_30,
   I3 => x115_out_5,
   I4 => x115_out_7,
   I5 => W_20_23_i_15_n_0,
   O => W_20_23_i_9_n_0
);
W_20_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_4_26,
   I1 => M_reg_13_26,
   I2 => M_reg_5_12,
   I3 => M_reg_5_1,
   I4 => M_reg_5_29,
   O => W_20_27_i_10_n_0
);
W_20_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_13_25,
   I1 => M_reg_5_28,
   I2 => M_reg_5_0,
   I3 => M_reg_5_11,
   I4 => M_reg_4_25,
   O => W_20_27_i_11_n_0
);
W_20_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_4_25,
   I1 => M_reg_13_25,
   I2 => M_reg_5_11,
   I3 => M_reg_5_0,
   I4 => M_reg_5_28,
   O => W_20_27_i_12_n_0
);
W_20_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_13_24,
   I1 => M_reg_5_27,
   I2 => M_reg_5_31,
   I3 => M_reg_5_10,
   I4 => M_reg_4_24,
   O => W_20_27_i_13_n_0
);
W_20_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_4_24,
   I1 => M_reg_13_24,
   I2 => M_reg_5_10,
   I3 => M_reg_5_31,
   I4 => M_reg_5_27,
   O => W_20_27_i_14_n_0
);
W_20_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_13_23,
   I1 => M_reg_5_26,
   I2 => M_reg_5_30,
   I3 => M_reg_5_9,
   I4 => M_reg_4_23,
   O => W_20_27_i_15_n_0
);
W_20_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_4_23,
   I1 => M_reg_13_23,
   I2 => M_reg_5_9,
   I3 => M_reg_5_30,
   I4 => M_reg_5_26,
   O => W_20_27_i_16_n_0
);
W_20_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_13_22,
   I1 => M_reg_5_25,
   I2 => M_reg_5_29,
   I3 => M_reg_5_8,
   I4 => M_reg_4_22,
   O => W_20_27_i_17_n_0
);
W_20_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x115_out_11,
   I1 => x115_out_13,
   I2 => W_20_27_i_10_n_0,
   I3 => W_20_27_i_11_n_0,
   O => W_20_27_i_2_n_0
);
W_20_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x115_out_10,
   I1 => x115_out_12,
   I2 => W_20_27_i_12_n_0,
   I3 => W_20_27_i_13_n_0,
   O => W_20_27_i_3_n_0
);
W_20_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x115_out_9,
   I1 => x115_out_11,
   I2 => W_20_27_i_14_n_0,
   I3 => W_20_27_i_15_n_0,
   O => W_20_27_i_4_n_0
);
W_20_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x115_out_8,
   I1 => x115_out_10,
   I2 => W_20_27_i_16_n_0,
   I3 => W_20_27_i_17_n_0,
   O => W_20_27_i_5_n_0
);
W_20_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x115_out_12,
   I1 => x115_out_14,
   I2 => W_20_31_i_13_n_0,
   I3 => W_20_31_i_14_n_0,
   I4 => W_20_27_i_2_n_0,
   O => W_20_27_i_6_n_0
);
W_20_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x115_out_11,
   I1 => x115_out_13,
   I2 => W_20_27_i_10_n_0,
   I3 => W_20_27_i_11_n_0,
   I4 => W_20_27_i_3_n_0,
   O => W_20_27_i_7_n_0
);
W_20_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x115_out_10,
   I1 => x115_out_12,
   I2 => W_20_27_i_12_n_0,
   I3 => W_20_27_i_13_n_0,
   I4 => W_20_27_i_4_n_0,
   O => W_20_27_i_8_n_0
);
W_20_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x115_out_9,
   I1 => x115_out_11,
   I2 => W_20_27_i_14_n_0,
   I3 => W_20_27_i_15_n_0,
   I4 => W_20_27_i_5_n_0,
   O => W_20_27_i_9_n_0
);
W_20_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_13_28,
   I1 => M_reg_5_31,
   I2 => M_reg_5_3,
   I3 => M_reg_5_14,
   I4 => M_reg_4_28,
   O => W_20_31_i_10_n_0
);
W_20_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_4_28,
   I1 => M_reg_13_28,
   I2 => M_reg_5_14,
   I3 => M_reg_5_3,
   I4 => M_reg_5_31,
   O => W_20_31_i_11_n_0
);
W_20_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_13_27,
   I1 => M_reg_5_30,
   I2 => M_reg_5_2,
   I3 => M_reg_5_13,
   I4 => M_reg_4_27,
   O => W_20_31_i_12_n_0
);
W_20_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_4_27,
   I1 => M_reg_13_27,
   I2 => M_reg_5_13,
   I3 => M_reg_5_2,
   I4 => M_reg_5_30,
   O => W_20_31_i_13_n_0
);
W_20_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_13_26,
   I1 => M_reg_5_29,
   I2 => M_reg_5_1,
   I3 => M_reg_5_12,
   I4 => M_reg_4_26,
   O => W_20_31_i_14_n_0
);
W_20_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => M_reg_13_29,
   I1 => M_reg_5_4,
   I2 => M_reg_5_15,
   I3 => M_reg_4_29,
   O => W_20_31_i_15_n_0
);
W_20_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x115_out_17,
   I1 => x115_out_15,
   O => SIGMA_LCASE_1355_out_30
);
W_20_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => M_reg_5_6,
   I1 => M_reg_5_17,
   I2 => M_reg_13_31,
   I3 => M_reg_4_31,
   I4 => x115_out_16,
   I5 => x115_out_18,
   O => W_20_31_i_17_n_0
);
W_20_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => M_reg_5_16,
   I1 => M_reg_5_5,
   O => SIGMA_LCASE_0351_out_30
);
W_20_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => M_reg_4_30,
   I1 => M_reg_13_30,
   I2 => M_reg_5_16,
   I3 => M_reg_5_5,
   O => W_20_31_i_19_n_0
);
W_20_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x115_out_14,
   I1 => x115_out_16,
   I2 => W_20_31_i_9_n_0,
   I3 => W_20_31_i_10_n_0,
   O => W_20_31_i_2_n_0
);
W_20_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x115_out_13,
   I1 => x115_out_15,
   I2 => W_20_31_i_11_n_0,
   I3 => W_20_31_i_12_n_0,
   O => W_20_31_i_3_n_0
);
W_20_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x115_out_12,
   I1 => x115_out_14,
   I2 => W_20_31_i_13_n_0,
   I3 => W_20_31_i_14_n_0,
   O => W_20_31_i_4_n_0
);
W_20_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_20_31_i_15_n_0,
   I1 => SIGMA_LCASE_1355_out_30,
   I2 => W_20_31_i_17_n_0,
   I3 => M_reg_13_30,
   I4 => SIGMA_LCASE_0351_out_30,
   I5 => M_reg_4_30,
   O => W_20_31_i_5_n_0
);
W_20_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_20_31_i_2_n_0,
   I1 => W_20_31_i_19_n_0,
   I2 => x115_out_15,
   I3 => x115_out_17,
   I4 => W_20_31_i_15_n_0,
   O => W_20_31_i_6_n_0
);
W_20_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x115_out_14,
   I1 => x115_out_16,
   I2 => W_20_31_i_9_n_0,
   I3 => W_20_31_i_10_n_0,
   I4 => W_20_31_i_3_n_0,
   O => W_20_31_i_7_n_0
);
W_20_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x115_out_13,
   I1 => x115_out_15,
   I2 => W_20_31_i_11_n_0,
   I3 => W_20_31_i_12_n_0,
   I4 => W_20_31_i_4_n_0,
   O => W_20_31_i_8_n_0
);
W_20_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => M_reg_4_29,
   I1 => M_reg_13_29,
   I2 => M_reg_5_15,
   I3 => M_reg_5_4,
   O => W_20_31_i_9_n_0
);
W_20_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_4_2,
   I1 => M_reg_13_2,
   I2 => M_reg_5_20,
   I3 => M_reg_5_9,
   I4 => M_reg_5_5,
   O => W_20_3_i_10_n_0
);
W_20_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_13_1,
   I1 => M_reg_5_4,
   I2 => M_reg_5_8,
   I3 => M_reg_5_19,
   I4 => M_reg_4_1,
   O => W_20_3_i_11_n_0
);
W_20_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => M_reg_5_19,
   I1 => M_reg_5_8,
   I2 => M_reg_5_4,
   O => SIGMA_LCASE_0351_out_1
);
W_20_3_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_4_1,
   I1 => M_reg_13_1,
   I2 => M_reg_5_19,
   I3 => M_reg_5_8,
   I4 => M_reg_5_4,
   O => W_20_3_i_13_n_0
);
W_20_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x115_out_12,
   I1 => x115_out_19,
   I2 => x115_out_21,
   I3 => W_20_3_i_10_n_0,
   I4 => W_20_3_i_11_n_0,
   O => W_20_3_i_2_n_0
);
W_20_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_20_3_i_11_n_0,
   I1 => x115_out_21,
   I2 => x115_out_19,
   I3 => x115_out_12,
   I4 => W_20_3_i_10_n_0,
   O => W_20_3_i_3_n_0
);
W_20_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_0351_out_1,
   I1 => M_reg_13_1,
   I2 => M_reg_4_1,
   I3 => x115_out_11,
   I4 => x115_out_18,
   I5 => x115_out_20,
   O => W_20_3_i_4_n_0
);
W_20_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_4_0,
   I1 => M_reg_13_0,
   I2 => M_reg_5_18,
   I3 => M_reg_5_7,
   I4 => M_reg_5_3,
   O => W_20_3_i_5_n_0
);
W_20_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_20_3_i_2_n_0,
   I1 => W_20_7_i_16_n_0,
   I2 => x115_out_13,
   I3 => x115_out_20,
   I4 => x115_out_22,
   I5 => W_20_7_i_17_n_0,
   O => W_20_3_i_6_n_0
);
W_20_3_i_7 : LUT5
  generic map(
   INIT => X"6aa6a66a"
  )
 port map (
   I0 => W_20_3_i_3_n_0,
   I1 => W_20_3_i_13_n_0,
   I2 => x115_out_20,
   I3 => x115_out_18,
   I4 => x115_out_11,
   O => W_20_3_i_7_n_0
);
W_20_3_i_8 : LUT6
  generic map(
   INIT => X"566565566aa6a66a"
  )
 port map (
   I0 => W_20_3_i_4_n_0,
   I1 => M_reg_4_0,
   I2 => M_reg_5_18,
   I3 => M_reg_5_7,
   I4 => M_reg_5_3,
   I5 => M_reg_13_0,
   O => W_20_3_i_8_n_0
);
W_20_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_20_3_i_5_n_0,
   I1 => x115_out_10,
   I2 => x115_out_17,
   I3 => x115_out_19,
   O => W_20_3_i_9_n_0
);
W_20_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_4_6,
   I1 => M_reg_13_6,
   I2 => M_reg_5_24,
   I3 => M_reg_5_13,
   I4 => M_reg_5_9,
   O => W_20_7_i_10_n_0
);
W_20_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_13_5,
   I1 => M_reg_5_8,
   I2 => M_reg_5_12,
   I3 => M_reg_5_23,
   I4 => M_reg_4_5,
   O => W_20_7_i_11_n_0
);
W_20_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_4_5,
   I1 => M_reg_13_5,
   I2 => M_reg_5_23,
   I3 => M_reg_5_12,
   I4 => M_reg_5_8,
   O => W_20_7_i_12_n_0
);
W_20_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_13_4,
   I1 => M_reg_5_7,
   I2 => M_reg_5_11,
   I3 => M_reg_5_22,
   I4 => M_reg_4_4,
   O => W_20_7_i_13_n_0
);
W_20_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_4_4,
   I1 => M_reg_13_4,
   I2 => M_reg_5_22,
   I3 => M_reg_5_11,
   I4 => M_reg_5_7,
   O => W_20_7_i_14_n_0
);
W_20_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_13_3,
   I1 => M_reg_5_6,
   I2 => M_reg_5_10,
   I3 => M_reg_5_21,
   I4 => M_reg_4_3,
   O => W_20_7_i_15_n_0
);
W_20_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_4_3,
   I1 => M_reg_13_3,
   I2 => M_reg_5_21,
   I3 => M_reg_5_10,
   I4 => M_reg_5_6,
   O => W_20_7_i_16_n_0
);
W_20_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_13_2,
   I1 => M_reg_5_5,
   I2 => M_reg_5_9,
   I3 => M_reg_5_20,
   I4 => M_reg_4_2,
   O => W_20_7_i_17_n_0
);
W_20_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x115_out_16,
   I1 => x115_out_23,
   I2 => x115_out_25,
   I3 => W_20_7_i_10_n_0,
   I4 => W_20_7_i_11_n_0,
   O => W_20_7_i_2_n_0
);
W_20_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x115_out_15,
   I1 => x115_out_22,
   I2 => x115_out_24,
   I3 => W_20_7_i_12_n_0,
   I4 => W_20_7_i_13_n_0,
   O => W_20_7_i_3_n_0
);
W_20_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x115_out_14,
   I1 => x115_out_21,
   I2 => x115_out_23,
   I3 => W_20_7_i_14_n_0,
   I4 => W_20_7_i_15_n_0,
   O => W_20_7_i_4_n_0
);
W_20_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x115_out_13,
   I1 => x115_out_20,
   I2 => x115_out_22,
   I3 => W_20_7_i_16_n_0,
   I4 => W_20_7_i_17_n_0,
   O => W_20_7_i_5_n_0
);
W_20_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_20_7_i_2_n_0,
   I1 => W_20_11_i_16_n_0,
   I2 => x115_out_17,
   I3 => x115_out_24,
   I4 => x115_out_26,
   I5 => W_20_11_i_17_n_0,
   O => W_20_7_i_6_n_0
);
W_20_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_20_7_i_3_n_0,
   I1 => W_20_7_i_10_n_0,
   I2 => x115_out_16,
   I3 => x115_out_23,
   I4 => x115_out_25,
   I5 => W_20_7_i_11_n_0,
   O => W_20_7_i_7_n_0
);
W_20_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_20_7_i_4_n_0,
   I1 => W_20_7_i_12_n_0,
   I2 => x115_out_15,
   I3 => x115_out_22,
   I4 => x115_out_24,
   I5 => W_20_7_i_13_n_0,
   O => W_20_7_i_8_n_0
);
W_20_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_20_7_i_5_n_0,
   I1 => W_20_7_i_14_n_0,
   I2 => x115_out_14,
   I3 => x115_out_21,
   I4 => x115_out_23,
   I5 => W_20_7_i_15_n_0,
   O => W_20_7_i_9_n_0
);
W_21_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_5_10,
   I1 => M_reg_14_10,
   I2 => M_reg_6_28,
   I3 => M_reg_6_17,
   I4 => M_reg_6_13,
   O => W_21_11_i_10_n_0
);
W_21_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_14_9,
   I1 => M_reg_6_12,
   I2 => M_reg_6_16,
   I3 => M_reg_6_27,
   I4 => M_reg_5_9,
   O => W_21_11_i_11_n_0
);
W_21_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_5_9,
   I1 => M_reg_14_9,
   I2 => M_reg_6_27,
   I3 => M_reg_6_16,
   I4 => M_reg_6_12,
   O => W_21_11_i_12_n_0
);
W_21_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_14_8,
   I1 => M_reg_6_11,
   I2 => M_reg_6_15,
   I3 => M_reg_6_26,
   I4 => M_reg_5_8,
   O => W_21_11_i_13_n_0
);
W_21_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_5_8,
   I1 => M_reg_14_8,
   I2 => M_reg_6_26,
   I3 => M_reg_6_15,
   I4 => M_reg_6_11,
   O => W_21_11_i_14_n_0
);
W_21_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_14_7,
   I1 => M_reg_6_10,
   I2 => M_reg_6_14,
   I3 => M_reg_6_25,
   I4 => M_reg_5_7,
   O => W_21_11_i_15_n_0
);
W_21_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_5_7,
   I1 => M_reg_14_7,
   I2 => M_reg_6_25,
   I3 => M_reg_6_14,
   I4 => M_reg_6_10,
   O => W_21_11_i_16_n_0
);
W_21_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_14_6,
   I1 => M_reg_6_9,
   I2 => M_reg_6_13,
   I3 => M_reg_6_24,
   I4 => M_reg_5_6,
   O => W_21_11_i_17_n_0
);
W_21_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x114_out_20,
   I1 => x114_out_27,
   I2 => x114_out_29,
   I3 => W_21_11_i_10_n_0,
   I4 => W_21_11_i_11_n_0,
   O => W_21_11_i_2_n_0
);
W_21_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x114_out_19,
   I1 => x114_out_26,
   I2 => x114_out_28,
   I3 => W_21_11_i_12_n_0,
   I4 => W_21_11_i_13_n_0,
   O => W_21_11_i_3_n_0
);
W_21_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x114_out_18,
   I1 => x114_out_25,
   I2 => x114_out_27,
   I3 => W_21_11_i_14_n_0,
   I4 => W_21_11_i_15_n_0,
   O => W_21_11_i_4_n_0
);
W_21_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x114_out_17,
   I1 => x114_out_24,
   I2 => x114_out_26,
   I3 => W_21_11_i_16_n_0,
   I4 => W_21_11_i_17_n_0,
   O => W_21_11_i_5_n_0
);
W_21_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_21_11_i_2_n_0,
   I1 => W_21_15_i_16_n_0,
   I2 => x114_out_21,
   I3 => x114_out_28,
   I4 => x114_out_30,
   I5 => W_21_15_i_17_n_0,
   O => W_21_11_i_6_n_0
);
W_21_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_21_11_i_3_n_0,
   I1 => W_21_11_i_10_n_0,
   I2 => x114_out_20,
   I3 => x114_out_27,
   I4 => x114_out_29,
   I5 => W_21_11_i_11_n_0,
   O => W_21_11_i_7_n_0
);
W_21_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_21_11_i_4_n_0,
   I1 => W_21_11_i_12_n_0,
   I2 => x114_out_19,
   I3 => x114_out_26,
   I4 => x114_out_28,
   I5 => W_21_11_i_13_n_0,
   O => W_21_11_i_8_n_0
);
W_21_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_21_11_i_5_n_0,
   I1 => W_21_11_i_14_n_0,
   I2 => x114_out_18,
   I3 => x114_out_25,
   I4 => x114_out_27,
   I5 => W_21_11_i_15_n_0,
   O => W_21_11_i_9_n_0
);
W_21_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_5_14,
   I1 => M_reg_14_14,
   I2 => M_reg_6_0,
   I3 => M_reg_6_21,
   I4 => M_reg_6_17,
   O => W_21_15_i_10_n_0
);
W_21_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_14_13,
   I1 => M_reg_6_16,
   I2 => M_reg_6_20,
   I3 => M_reg_6_31,
   I4 => M_reg_5_13,
   O => W_21_15_i_11_n_0
);
W_21_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_5_13,
   I1 => M_reg_14_13,
   I2 => M_reg_6_31,
   I3 => M_reg_6_20,
   I4 => M_reg_6_16,
   O => W_21_15_i_12_n_0
);
W_21_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_14_12,
   I1 => M_reg_6_15,
   I2 => M_reg_6_19,
   I3 => M_reg_6_30,
   I4 => M_reg_5_12,
   O => W_21_15_i_13_n_0
);
W_21_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_5_12,
   I1 => M_reg_14_12,
   I2 => M_reg_6_30,
   I3 => M_reg_6_19,
   I4 => M_reg_6_15,
   O => W_21_15_i_14_n_0
);
W_21_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_14_11,
   I1 => M_reg_6_14,
   I2 => M_reg_6_18,
   I3 => M_reg_6_29,
   I4 => M_reg_5_11,
   O => W_21_15_i_15_n_0
);
W_21_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_5_11,
   I1 => M_reg_14_11,
   I2 => M_reg_6_29,
   I3 => M_reg_6_18,
   I4 => M_reg_6_14,
   O => W_21_15_i_16_n_0
);
W_21_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_14_10,
   I1 => M_reg_6_13,
   I2 => M_reg_6_17,
   I3 => M_reg_6_28,
   I4 => M_reg_5_10,
   O => W_21_15_i_17_n_0
);
W_21_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x114_out_24,
   I1 => x114_out_31,
   I2 => x114_out_1,
   I3 => W_21_15_i_10_n_0,
   I4 => W_21_15_i_11_n_0,
   O => W_21_15_i_2_n_0
);
W_21_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x114_out_23,
   I1 => x114_out_30,
   I2 => x114_out_0,
   I3 => W_21_15_i_12_n_0,
   I4 => W_21_15_i_13_n_0,
   O => W_21_15_i_3_n_0
);
W_21_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x114_out_22,
   I1 => x114_out_29,
   I2 => x114_out_31,
   I3 => W_21_15_i_14_n_0,
   I4 => W_21_15_i_15_n_0,
   O => W_21_15_i_4_n_0
);
W_21_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x114_out_21,
   I1 => x114_out_28,
   I2 => x114_out_30,
   I3 => W_21_15_i_16_n_0,
   I4 => W_21_15_i_17_n_0,
   O => W_21_15_i_5_n_0
);
W_21_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_21_15_i_2_n_0,
   I1 => W_21_19_i_16_n_0,
   I2 => x114_out_25,
   I3 => x114_out_0,
   I4 => x114_out_2,
   I5 => W_21_19_i_17_n_0,
   O => W_21_15_i_6_n_0
);
W_21_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_21_15_i_3_n_0,
   I1 => W_21_15_i_10_n_0,
   I2 => x114_out_24,
   I3 => x114_out_31,
   I4 => x114_out_1,
   I5 => W_21_15_i_11_n_0,
   O => W_21_15_i_7_n_0
);
W_21_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_21_15_i_4_n_0,
   I1 => W_21_15_i_12_n_0,
   I2 => x114_out_23,
   I3 => x114_out_30,
   I4 => x114_out_0,
   I5 => W_21_15_i_13_n_0,
   O => W_21_15_i_8_n_0
);
W_21_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_21_15_i_5_n_0,
   I1 => W_21_15_i_14_n_0,
   I2 => x114_out_22,
   I3 => x114_out_29,
   I4 => x114_out_31,
   I5 => W_21_15_i_15_n_0,
   O => W_21_15_i_9_n_0
);
W_21_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_5_18,
   I1 => M_reg_14_18,
   I2 => M_reg_6_4,
   I3 => M_reg_6_25,
   I4 => M_reg_6_21,
   O => W_21_19_i_10_n_0
);
W_21_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_14_17,
   I1 => M_reg_6_20,
   I2 => M_reg_6_24,
   I3 => M_reg_6_3,
   I4 => M_reg_5_17,
   O => W_21_19_i_11_n_0
);
W_21_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_5_17,
   I1 => M_reg_14_17,
   I2 => M_reg_6_3,
   I3 => M_reg_6_24,
   I4 => M_reg_6_20,
   O => W_21_19_i_12_n_0
);
W_21_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_14_16,
   I1 => M_reg_6_19,
   I2 => M_reg_6_23,
   I3 => M_reg_6_2,
   I4 => M_reg_5_16,
   O => W_21_19_i_13_n_0
);
W_21_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_5_16,
   I1 => M_reg_14_16,
   I2 => M_reg_6_2,
   I3 => M_reg_6_23,
   I4 => M_reg_6_19,
   O => W_21_19_i_14_n_0
);
W_21_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_14_15,
   I1 => M_reg_6_18,
   I2 => M_reg_6_22,
   I3 => M_reg_6_1,
   I4 => M_reg_5_15,
   O => W_21_19_i_15_n_0
);
W_21_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_5_15,
   I1 => M_reg_14_15,
   I2 => M_reg_6_1,
   I3 => M_reg_6_22,
   I4 => M_reg_6_18,
   O => W_21_19_i_16_n_0
);
W_21_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_14_14,
   I1 => M_reg_6_17,
   I2 => M_reg_6_21,
   I3 => M_reg_6_0,
   I4 => M_reg_5_14,
   O => W_21_19_i_17_n_0
);
W_21_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x114_out_28,
   I1 => x114_out_3,
   I2 => x114_out_5,
   I3 => W_21_19_i_10_n_0,
   I4 => W_21_19_i_11_n_0,
   O => W_21_19_i_2_n_0
);
W_21_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x114_out_27,
   I1 => x114_out_2,
   I2 => x114_out_4,
   I3 => W_21_19_i_12_n_0,
   I4 => W_21_19_i_13_n_0,
   O => W_21_19_i_3_n_0
);
W_21_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x114_out_26,
   I1 => x114_out_1,
   I2 => x114_out_3,
   I3 => W_21_19_i_14_n_0,
   I4 => W_21_19_i_15_n_0,
   O => W_21_19_i_4_n_0
);
W_21_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x114_out_25,
   I1 => x114_out_0,
   I2 => x114_out_2,
   I3 => W_21_19_i_16_n_0,
   I4 => W_21_19_i_17_n_0,
   O => W_21_19_i_5_n_0
);
W_21_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_21_19_i_2_n_0,
   I1 => W_21_23_i_16_n_0,
   I2 => x114_out_29,
   I3 => x114_out_4,
   I4 => x114_out_6,
   I5 => W_21_23_i_17_n_0,
   O => W_21_19_i_6_n_0
);
W_21_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_21_19_i_3_n_0,
   I1 => W_21_19_i_10_n_0,
   I2 => x114_out_28,
   I3 => x114_out_3,
   I4 => x114_out_5,
   I5 => W_21_19_i_11_n_0,
   O => W_21_19_i_7_n_0
);
W_21_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_21_19_i_4_n_0,
   I1 => W_21_19_i_12_n_0,
   I2 => x114_out_27,
   I3 => x114_out_2,
   I4 => x114_out_4,
   I5 => W_21_19_i_13_n_0,
   O => W_21_19_i_8_n_0
);
W_21_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_21_19_i_5_n_0,
   I1 => W_21_19_i_14_n_0,
   I2 => x114_out_26,
   I3 => x114_out_1,
   I4 => x114_out_3,
   I5 => W_21_19_i_15_n_0,
   O => W_21_19_i_9_n_0
);
W_21_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_5_22,
   I1 => M_reg_14_22,
   I2 => M_reg_6_8,
   I3 => M_reg_6_29,
   I4 => M_reg_6_25,
   O => W_21_23_i_10_n_0
);
W_21_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_14_21,
   I1 => M_reg_6_24,
   I2 => M_reg_6_28,
   I3 => M_reg_6_7,
   I4 => M_reg_5_21,
   O => W_21_23_i_11_n_0
);
W_21_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_5_21,
   I1 => M_reg_14_21,
   I2 => M_reg_6_7,
   I3 => M_reg_6_28,
   I4 => M_reg_6_24,
   O => W_21_23_i_12_n_0
);
W_21_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_14_20,
   I1 => M_reg_6_23,
   I2 => M_reg_6_27,
   I3 => M_reg_6_6,
   I4 => M_reg_5_20,
   O => W_21_23_i_13_n_0
);
W_21_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_5_20,
   I1 => M_reg_14_20,
   I2 => M_reg_6_6,
   I3 => M_reg_6_27,
   I4 => M_reg_6_23,
   O => W_21_23_i_14_n_0
);
W_21_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_14_19,
   I1 => M_reg_6_22,
   I2 => M_reg_6_26,
   I3 => M_reg_6_5,
   I4 => M_reg_5_19,
   O => W_21_23_i_15_n_0
);
W_21_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_5_19,
   I1 => M_reg_14_19,
   I2 => M_reg_6_5,
   I3 => M_reg_6_26,
   I4 => M_reg_6_22,
   O => W_21_23_i_16_n_0
);
W_21_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_14_18,
   I1 => M_reg_6_21,
   I2 => M_reg_6_25,
   I3 => M_reg_6_4,
   I4 => M_reg_5_18,
   O => W_21_23_i_17_n_0
);
W_21_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x114_out_7,
   I1 => x114_out_9,
   I2 => W_21_23_i_10_n_0,
   I3 => W_21_23_i_11_n_0,
   O => W_21_23_i_2_n_0
);
W_21_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x114_out_31,
   I1 => x114_out_6,
   I2 => x114_out_8,
   I3 => W_21_23_i_12_n_0,
   I4 => W_21_23_i_13_n_0,
   O => W_21_23_i_3_n_0
);
W_21_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x114_out_30,
   I1 => x114_out_5,
   I2 => x114_out_7,
   I3 => W_21_23_i_14_n_0,
   I4 => W_21_23_i_15_n_0,
   O => W_21_23_i_4_n_0
);
W_21_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x114_out_29,
   I1 => x114_out_4,
   I2 => x114_out_6,
   I3 => W_21_23_i_16_n_0,
   I4 => W_21_23_i_17_n_0,
   O => W_21_23_i_5_n_0
);
W_21_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x114_out_8,
   I1 => x114_out_10,
   I2 => W_21_27_i_16_n_0,
   I3 => W_21_27_i_17_n_0,
   I4 => W_21_23_i_2_n_0,
   O => W_21_23_i_6_n_0
);
W_21_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x114_out_7,
   I1 => x114_out_9,
   I2 => W_21_23_i_10_n_0,
   I3 => W_21_23_i_11_n_0,
   I4 => W_21_23_i_3_n_0,
   O => W_21_23_i_7_n_0
);
W_21_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_21_23_i_4_n_0,
   I1 => W_21_23_i_12_n_0,
   I2 => x114_out_31,
   I3 => x114_out_6,
   I4 => x114_out_8,
   I5 => W_21_23_i_13_n_0,
   O => W_21_23_i_8_n_0
);
W_21_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_21_23_i_5_n_0,
   I1 => W_21_23_i_14_n_0,
   I2 => x114_out_30,
   I3 => x114_out_5,
   I4 => x114_out_7,
   I5 => W_21_23_i_15_n_0,
   O => W_21_23_i_9_n_0
);
W_21_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_5_26,
   I1 => M_reg_14_26,
   I2 => M_reg_6_12,
   I3 => M_reg_6_1,
   I4 => M_reg_6_29,
   O => W_21_27_i_10_n_0
);
W_21_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_14_25,
   I1 => M_reg_6_28,
   I2 => M_reg_6_0,
   I3 => M_reg_6_11,
   I4 => M_reg_5_25,
   O => W_21_27_i_11_n_0
);
W_21_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_5_25,
   I1 => M_reg_14_25,
   I2 => M_reg_6_11,
   I3 => M_reg_6_0,
   I4 => M_reg_6_28,
   O => W_21_27_i_12_n_0
);
W_21_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_14_24,
   I1 => M_reg_6_27,
   I2 => M_reg_6_31,
   I3 => M_reg_6_10,
   I4 => M_reg_5_24,
   O => W_21_27_i_13_n_0
);
W_21_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_5_24,
   I1 => M_reg_14_24,
   I2 => M_reg_6_10,
   I3 => M_reg_6_31,
   I4 => M_reg_6_27,
   O => W_21_27_i_14_n_0
);
W_21_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_14_23,
   I1 => M_reg_6_26,
   I2 => M_reg_6_30,
   I3 => M_reg_6_9,
   I4 => M_reg_5_23,
   O => W_21_27_i_15_n_0
);
W_21_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_5_23,
   I1 => M_reg_14_23,
   I2 => M_reg_6_9,
   I3 => M_reg_6_30,
   I4 => M_reg_6_26,
   O => W_21_27_i_16_n_0
);
W_21_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_14_22,
   I1 => M_reg_6_25,
   I2 => M_reg_6_29,
   I3 => M_reg_6_8,
   I4 => M_reg_5_22,
   O => W_21_27_i_17_n_0
);
W_21_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x114_out_11,
   I1 => x114_out_13,
   I2 => W_21_27_i_10_n_0,
   I3 => W_21_27_i_11_n_0,
   O => W_21_27_i_2_n_0
);
W_21_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x114_out_10,
   I1 => x114_out_12,
   I2 => W_21_27_i_12_n_0,
   I3 => W_21_27_i_13_n_0,
   O => W_21_27_i_3_n_0
);
W_21_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x114_out_9,
   I1 => x114_out_11,
   I2 => W_21_27_i_14_n_0,
   I3 => W_21_27_i_15_n_0,
   O => W_21_27_i_4_n_0
);
W_21_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x114_out_8,
   I1 => x114_out_10,
   I2 => W_21_27_i_16_n_0,
   I3 => W_21_27_i_17_n_0,
   O => W_21_27_i_5_n_0
);
W_21_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x114_out_12,
   I1 => x114_out_14,
   I2 => W_21_31_i_13_n_0,
   I3 => W_21_31_i_14_n_0,
   I4 => W_21_27_i_2_n_0,
   O => W_21_27_i_6_n_0
);
W_21_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x114_out_11,
   I1 => x114_out_13,
   I2 => W_21_27_i_10_n_0,
   I3 => W_21_27_i_11_n_0,
   I4 => W_21_27_i_3_n_0,
   O => W_21_27_i_7_n_0
);
W_21_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x114_out_10,
   I1 => x114_out_12,
   I2 => W_21_27_i_12_n_0,
   I3 => W_21_27_i_13_n_0,
   I4 => W_21_27_i_4_n_0,
   O => W_21_27_i_8_n_0
);
W_21_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x114_out_9,
   I1 => x114_out_11,
   I2 => W_21_27_i_14_n_0,
   I3 => W_21_27_i_15_n_0,
   I4 => W_21_27_i_5_n_0,
   O => W_21_27_i_9_n_0
);
W_21_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_14_28,
   I1 => M_reg_6_31,
   I2 => M_reg_6_3,
   I3 => M_reg_6_14,
   I4 => M_reg_5_28,
   O => W_21_31_i_10_n_0
);
W_21_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_5_28,
   I1 => M_reg_14_28,
   I2 => M_reg_6_14,
   I3 => M_reg_6_3,
   I4 => M_reg_6_31,
   O => W_21_31_i_11_n_0
);
W_21_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_14_27,
   I1 => M_reg_6_30,
   I2 => M_reg_6_2,
   I3 => M_reg_6_13,
   I4 => M_reg_5_27,
   O => W_21_31_i_12_n_0
);
W_21_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_5_27,
   I1 => M_reg_14_27,
   I2 => M_reg_6_13,
   I3 => M_reg_6_2,
   I4 => M_reg_6_30,
   O => W_21_31_i_13_n_0
);
W_21_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_14_26,
   I1 => M_reg_6_29,
   I2 => M_reg_6_1,
   I3 => M_reg_6_12,
   I4 => M_reg_5_26,
   O => W_21_31_i_14_n_0
);
W_21_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => M_reg_14_29,
   I1 => M_reg_6_4,
   I2 => M_reg_6_15,
   I3 => M_reg_5_29,
   O => W_21_31_i_15_n_0
);
W_21_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x114_out_17,
   I1 => x114_out_15,
   O => SIGMA_LCASE_1347_out_30
);
W_21_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => M_reg_6_6,
   I1 => M_reg_6_17,
   I2 => M_reg_14_31,
   I3 => M_reg_5_31,
   I4 => x114_out_16,
   I5 => x114_out_18,
   O => W_21_31_i_17_n_0
);
W_21_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => M_reg_6_16,
   I1 => M_reg_6_5,
   O => SIGMA_LCASE_0343_out_30
);
W_21_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => M_reg_5_30,
   I1 => M_reg_14_30,
   I2 => M_reg_6_16,
   I3 => M_reg_6_5,
   O => W_21_31_i_19_n_0
);
W_21_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x114_out_14,
   I1 => x114_out_16,
   I2 => W_21_31_i_9_n_0,
   I3 => W_21_31_i_10_n_0,
   O => W_21_31_i_2_n_0
);
W_21_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x114_out_13,
   I1 => x114_out_15,
   I2 => W_21_31_i_11_n_0,
   I3 => W_21_31_i_12_n_0,
   O => W_21_31_i_3_n_0
);
W_21_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x114_out_12,
   I1 => x114_out_14,
   I2 => W_21_31_i_13_n_0,
   I3 => W_21_31_i_14_n_0,
   O => W_21_31_i_4_n_0
);
W_21_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_21_31_i_15_n_0,
   I1 => SIGMA_LCASE_1347_out_30,
   I2 => W_21_31_i_17_n_0,
   I3 => M_reg_14_30,
   I4 => SIGMA_LCASE_0343_out_30,
   I5 => M_reg_5_30,
   O => W_21_31_i_5_n_0
);
W_21_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_21_31_i_2_n_0,
   I1 => W_21_31_i_19_n_0,
   I2 => x114_out_15,
   I3 => x114_out_17,
   I4 => W_21_31_i_15_n_0,
   O => W_21_31_i_6_n_0
);
W_21_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x114_out_14,
   I1 => x114_out_16,
   I2 => W_21_31_i_9_n_0,
   I3 => W_21_31_i_10_n_0,
   I4 => W_21_31_i_3_n_0,
   O => W_21_31_i_7_n_0
);
W_21_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x114_out_13,
   I1 => x114_out_15,
   I2 => W_21_31_i_11_n_0,
   I3 => W_21_31_i_12_n_0,
   I4 => W_21_31_i_4_n_0,
   O => W_21_31_i_8_n_0
);
W_21_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => M_reg_5_29,
   I1 => M_reg_14_29,
   I2 => M_reg_6_15,
   I3 => M_reg_6_4,
   O => W_21_31_i_9_n_0
);
W_21_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_5_2,
   I1 => M_reg_14_2,
   I2 => M_reg_6_20,
   I3 => M_reg_6_9,
   I4 => M_reg_6_5,
   O => W_21_3_i_10_n_0
);
W_21_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_14_1,
   I1 => M_reg_6_4,
   I2 => M_reg_6_8,
   I3 => M_reg_6_19,
   I4 => M_reg_5_1,
   O => W_21_3_i_11_n_0
);
W_21_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => M_reg_6_19,
   I1 => M_reg_6_8,
   I2 => M_reg_6_4,
   O => SIGMA_LCASE_0343_out_1
);
W_21_3_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_5_1,
   I1 => M_reg_14_1,
   I2 => M_reg_6_19,
   I3 => M_reg_6_8,
   I4 => M_reg_6_4,
   O => W_21_3_i_13_n_0
);
W_21_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x114_out_12,
   I1 => x114_out_19,
   I2 => x114_out_21,
   I3 => W_21_3_i_10_n_0,
   I4 => W_21_3_i_11_n_0,
   O => W_21_3_i_2_n_0
);
W_21_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_21_3_i_11_n_0,
   I1 => x114_out_21,
   I2 => x114_out_19,
   I3 => x114_out_12,
   I4 => W_21_3_i_10_n_0,
   O => W_21_3_i_3_n_0
);
W_21_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_0343_out_1,
   I1 => M_reg_14_1,
   I2 => M_reg_5_1,
   I3 => x114_out_11,
   I4 => x114_out_18,
   I5 => x114_out_20,
   O => W_21_3_i_4_n_0
);
W_21_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_5_0,
   I1 => M_reg_14_0,
   I2 => M_reg_6_18,
   I3 => M_reg_6_7,
   I4 => M_reg_6_3,
   O => W_21_3_i_5_n_0
);
W_21_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_21_3_i_2_n_0,
   I1 => W_21_7_i_16_n_0,
   I2 => x114_out_13,
   I3 => x114_out_20,
   I4 => x114_out_22,
   I5 => W_21_7_i_17_n_0,
   O => W_21_3_i_6_n_0
);
W_21_3_i_7 : LUT5
  generic map(
   INIT => X"6aa6a66a"
  )
 port map (
   I0 => W_21_3_i_3_n_0,
   I1 => W_21_3_i_13_n_0,
   I2 => x114_out_20,
   I3 => x114_out_18,
   I4 => x114_out_11,
   O => W_21_3_i_7_n_0
);
W_21_3_i_8 : LUT6
  generic map(
   INIT => X"566565566aa6a66a"
  )
 port map (
   I0 => W_21_3_i_4_n_0,
   I1 => M_reg_5_0,
   I2 => M_reg_6_18,
   I3 => M_reg_6_7,
   I4 => M_reg_6_3,
   I5 => M_reg_14_0,
   O => W_21_3_i_8_n_0
);
W_21_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_21_3_i_5_n_0,
   I1 => x114_out_10,
   I2 => x114_out_17,
   I3 => x114_out_19,
   O => W_21_3_i_9_n_0
);
W_21_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_5_6,
   I1 => M_reg_14_6,
   I2 => M_reg_6_24,
   I3 => M_reg_6_13,
   I4 => M_reg_6_9,
   O => W_21_7_i_10_n_0
);
W_21_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_14_5,
   I1 => M_reg_6_8,
   I2 => M_reg_6_12,
   I3 => M_reg_6_23,
   I4 => M_reg_5_5,
   O => W_21_7_i_11_n_0
);
W_21_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_5_5,
   I1 => M_reg_14_5,
   I2 => M_reg_6_23,
   I3 => M_reg_6_12,
   I4 => M_reg_6_8,
   O => W_21_7_i_12_n_0
);
W_21_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_14_4,
   I1 => M_reg_6_7,
   I2 => M_reg_6_11,
   I3 => M_reg_6_22,
   I4 => M_reg_5_4,
   O => W_21_7_i_13_n_0
);
W_21_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_5_4,
   I1 => M_reg_14_4,
   I2 => M_reg_6_22,
   I3 => M_reg_6_11,
   I4 => M_reg_6_7,
   O => W_21_7_i_14_n_0
);
W_21_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_14_3,
   I1 => M_reg_6_6,
   I2 => M_reg_6_10,
   I3 => M_reg_6_21,
   I4 => M_reg_5_3,
   O => W_21_7_i_15_n_0
);
W_21_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_5_3,
   I1 => M_reg_14_3,
   I2 => M_reg_6_21,
   I3 => M_reg_6_10,
   I4 => M_reg_6_6,
   O => W_21_7_i_16_n_0
);
W_21_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_14_2,
   I1 => M_reg_6_5,
   I2 => M_reg_6_9,
   I3 => M_reg_6_20,
   I4 => M_reg_5_2,
   O => W_21_7_i_17_n_0
);
W_21_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x114_out_16,
   I1 => x114_out_23,
   I2 => x114_out_25,
   I3 => W_21_7_i_10_n_0,
   I4 => W_21_7_i_11_n_0,
   O => W_21_7_i_2_n_0
);
W_21_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x114_out_15,
   I1 => x114_out_22,
   I2 => x114_out_24,
   I3 => W_21_7_i_12_n_0,
   I4 => W_21_7_i_13_n_0,
   O => W_21_7_i_3_n_0
);
W_21_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x114_out_14,
   I1 => x114_out_21,
   I2 => x114_out_23,
   I3 => W_21_7_i_14_n_0,
   I4 => W_21_7_i_15_n_0,
   O => W_21_7_i_4_n_0
);
W_21_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x114_out_13,
   I1 => x114_out_20,
   I2 => x114_out_22,
   I3 => W_21_7_i_16_n_0,
   I4 => W_21_7_i_17_n_0,
   O => W_21_7_i_5_n_0
);
W_21_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_21_7_i_2_n_0,
   I1 => W_21_11_i_16_n_0,
   I2 => x114_out_17,
   I3 => x114_out_24,
   I4 => x114_out_26,
   I5 => W_21_11_i_17_n_0,
   O => W_21_7_i_6_n_0
);
W_21_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_21_7_i_3_n_0,
   I1 => W_21_7_i_10_n_0,
   I2 => x114_out_16,
   I3 => x114_out_23,
   I4 => x114_out_25,
   I5 => W_21_7_i_11_n_0,
   O => W_21_7_i_7_n_0
);
W_21_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_21_7_i_4_n_0,
   I1 => W_21_7_i_12_n_0,
   I2 => x114_out_15,
   I3 => x114_out_22,
   I4 => x114_out_24,
   I5 => W_21_7_i_13_n_0,
   O => W_21_7_i_8_n_0
);
W_21_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_21_7_i_5_n_0,
   I1 => W_21_7_i_14_n_0,
   I2 => x114_out_14,
   I3 => x114_out_21,
   I4 => x114_out_23,
   I5 => W_21_7_i_15_n_0,
   O => W_21_7_i_9_n_0
);
W_22_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_6_10,
   I1 => M_reg_15_10,
   I2 => M_reg_7_28,
   I3 => M_reg_7_17,
   I4 => M_reg_7_13,
   O => W_22_11_i_10_n_0
);
W_22_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_15_9,
   I1 => M_reg_7_12,
   I2 => M_reg_7_16,
   I3 => M_reg_7_27,
   I4 => M_reg_6_9,
   O => W_22_11_i_11_n_0
);
W_22_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_6_9,
   I1 => M_reg_15_9,
   I2 => M_reg_7_27,
   I3 => M_reg_7_16,
   I4 => M_reg_7_12,
   O => W_22_11_i_12_n_0
);
W_22_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_15_8,
   I1 => M_reg_7_11,
   I2 => M_reg_7_15,
   I3 => M_reg_7_26,
   I4 => M_reg_6_8,
   O => W_22_11_i_13_n_0
);
W_22_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_6_8,
   I1 => M_reg_15_8,
   I2 => M_reg_7_26,
   I3 => M_reg_7_15,
   I4 => M_reg_7_11,
   O => W_22_11_i_14_n_0
);
W_22_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_15_7,
   I1 => M_reg_7_10,
   I2 => M_reg_7_14,
   I3 => M_reg_7_25,
   I4 => M_reg_6_7,
   O => W_22_11_i_15_n_0
);
W_22_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_6_7,
   I1 => M_reg_15_7,
   I2 => M_reg_7_25,
   I3 => M_reg_7_14,
   I4 => M_reg_7_10,
   O => W_22_11_i_16_n_0
);
W_22_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_15_6,
   I1 => M_reg_7_9,
   I2 => M_reg_7_13,
   I3 => M_reg_7_24,
   I4 => M_reg_6_6,
   O => W_22_11_i_17_n_0
);
W_22_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x113_out_20,
   I1 => x113_out_27,
   I2 => x113_out_29,
   I3 => W_22_11_i_10_n_0,
   I4 => W_22_11_i_11_n_0,
   O => W_22_11_i_2_n_0
);
W_22_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x113_out_19,
   I1 => x113_out_26,
   I2 => x113_out_28,
   I3 => W_22_11_i_12_n_0,
   I4 => W_22_11_i_13_n_0,
   O => W_22_11_i_3_n_0
);
W_22_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x113_out_18,
   I1 => x113_out_25,
   I2 => x113_out_27,
   I3 => W_22_11_i_14_n_0,
   I4 => W_22_11_i_15_n_0,
   O => W_22_11_i_4_n_0
);
W_22_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x113_out_17,
   I1 => x113_out_24,
   I2 => x113_out_26,
   I3 => W_22_11_i_16_n_0,
   I4 => W_22_11_i_17_n_0,
   O => W_22_11_i_5_n_0
);
W_22_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_22_11_i_2_n_0,
   I1 => W_22_15_i_16_n_0,
   I2 => x113_out_21,
   I3 => x113_out_28,
   I4 => x113_out_30,
   I5 => W_22_15_i_17_n_0,
   O => W_22_11_i_6_n_0
);
W_22_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_22_11_i_3_n_0,
   I1 => W_22_11_i_10_n_0,
   I2 => x113_out_20,
   I3 => x113_out_27,
   I4 => x113_out_29,
   I5 => W_22_11_i_11_n_0,
   O => W_22_11_i_7_n_0
);
W_22_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_22_11_i_4_n_0,
   I1 => W_22_11_i_12_n_0,
   I2 => x113_out_19,
   I3 => x113_out_26,
   I4 => x113_out_28,
   I5 => W_22_11_i_13_n_0,
   O => W_22_11_i_8_n_0
);
W_22_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_22_11_i_5_n_0,
   I1 => W_22_11_i_14_n_0,
   I2 => x113_out_18,
   I3 => x113_out_25,
   I4 => x113_out_27,
   I5 => W_22_11_i_15_n_0,
   O => W_22_11_i_9_n_0
);
W_22_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_6_14,
   I1 => M_reg_15_14,
   I2 => M_reg_7_0,
   I3 => M_reg_7_21,
   I4 => M_reg_7_17,
   O => W_22_15_i_10_n_0
);
W_22_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_15_13,
   I1 => M_reg_7_16,
   I2 => M_reg_7_20,
   I3 => M_reg_7_31,
   I4 => M_reg_6_13,
   O => W_22_15_i_11_n_0
);
W_22_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_6_13,
   I1 => M_reg_15_13,
   I2 => M_reg_7_31,
   I3 => M_reg_7_20,
   I4 => M_reg_7_16,
   O => W_22_15_i_12_n_0
);
W_22_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_15_12,
   I1 => M_reg_7_15,
   I2 => M_reg_7_19,
   I3 => M_reg_7_30,
   I4 => M_reg_6_12,
   O => W_22_15_i_13_n_0
);
W_22_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_6_12,
   I1 => M_reg_15_12,
   I2 => M_reg_7_30,
   I3 => M_reg_7_19,
   I4 => M_reg_7_15,
   O => W_22_15_i_14_n_0
);
W_22_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_15_11,
   I1 => M_reg_7_14,
   I2 => M_reg_7_18,
   I3 => M_reg_7_29,
   I4 => M_reg_6_11,
   O => W_22_15_i_15_n_0
);
W_22_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_6_11,
   I1 => M_reg_15_11,
   I2 => M_reg_7_29,
   I3 => M_reg_7_18,
   I4 => M_reg_7_14,
   O => W_22_15_i_16_n_0
);
W_22_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_15_10,
   I1 => M_reg_7_13,
   I2 => M_reg_7_17,
   I3 => M_reg_7_28,
   I4 => M_reg_6_10,
   O => W_22_15_i_17_n_0
);
W_22_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x113_out_24,
   I1 => x113_out_31,
   I2 => x113_out_1,
   I3 => W_22_15_i_10_n_0,
   I4 => W_22_15_i_11_n_0,
   O => W_22_15_i_2_n_0
);
W_22_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x113_out_23,
   I1 => x113_out_30,
   I2 => x113_out_0,
   I3 => W_22_15_i_12_n_0,
   I4 => W_22_15_i_13_n_0,
   O => W_22_15_i_3_n_0
);
W_22_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x113_out_22,
   I1 => x113_out_29,
   I2 => x113_out_31,
   I3 => W_22_15_i_14_n_0,
   I4 => W_22_15_i_15_n_0,
   O => W_22_15_i_4_n_0
);
W_22_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x113_out_21,
   I1 => x113_out_28,
   I2 => x113_out_30,
   I3 => W_22_15_i_16_n_0,
   I4 => W_22_15_i_17_n_0,
   O => W_22_15_i_5_n_0
);
W_22_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_22_15_i_2_n_0,
   I1 => W_22_19_i_16_n_0,
   I2 => x113_out_25,
   I3 => x113_out_0,
   I4 => x113_out_2,
   I5 => W_22_19_i_17_n_0,
   O => W_22_15_i_6_n_0
);
W_22_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_22_15_i_3_n_0,
   I1 => W_22_15_i_10_n_0,
   I2 => x113_out_24,
   I3 => x113_out_31,
   I4 => x113_out_1,
   I5 => W_22_15_i_11_n_0,
   O => W_22_15_i_7_n_0
);
W_22_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_22_15_i_4_n_0,
   I1 => W_22_15_i_12_n_0,
   I2 => x113_out_23,
   I3 => x113_out_30,
   I4 => x113_out_0,
   I5 => W_22_15_i_13_n_0,
   O => W_22_15_i_8_n_0
);
W_22_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_22_15_i_5_n_0,
   I1 => W_22_15_i_14_n_0,
   I2 => x113_out_22,
   I3 => x113_out_29,
   I4 => x113_out_31,
   I5 => W_22_15_i_15_n_0,
   O => W_22_15_i_9_n_0
);
W_22_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_6_18,
   I1 => M_reg_15_18,
   I2 => M_reg_7_4,
   I3 => M_reg_7_25,
   I4 => M_reg_7_21,
   O => W_22_19_i_10_n_0
);
W_22_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_15_17,
   I1 => M_reg_7_20,
   I2 => M_reg_7_24,
   I3 => M_reg_7_3,
   I4 => M_reg_6_17,
   O => W_22_19_i_11_n_0
);
W_22_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_6_17,
   I1 => M_reg_15_17,
   I2 => M_reg_7_3,
   I3 => M_reg_7_24,
   I4 => M_reg_7_20,
   O => W_22_19_i_12_n_0
);
W_22_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_15_16,
   I1 => M_reg_7_19,
   I2 => M_reg_7_23,
   I3 => M_reg_7_2,
   I4 => M_reg_6_16,
   O => W_22_19_i_13_n_0
);
W_22_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_6_16,
   I1 => M_reg_15_16,
   I2 => M_reg_7_2,
   I3 => M_reg_7_23,
   I4 => M_reg_7_19,
   O => W_22_19_i_14_n_0
);
W_22_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_15_15,
   I1 => M_reg_7_18,
   I2 => M_reg_7_22,
   I3 => M_reg_7_1,
   I4 => M_reg_6_15,
   O => W_22_19_i_15_n_0
);
W_22_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_6_15,
   I1 => M_reg_15_15,
   I2 => M_reg_7_1,
   I3 => M_reg_7_22,
   I4 => M_reg_7_18,
   O => W_22_19_i_16_n_0
);
W_22_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_15_14,
   I1 => M_reg_7_17,
   I2 => M_reg_7_21,
   I3 => M_reg_7_0,
   I4 => M_reg_6_14,
   O => W_22_19_i_17_n_0
);
W_22_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x113_out_28,
   I1 => x113_out_3,
   I2 => x113_out_5,
   I3 => W_22_19_i_10_n_0,
   I4 => W_22_19_i_11_n_0,
   O => W_22_19_i_2_n_0
);
W_22_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x113_out_27,
   I1 => x113_out_2,
   I2 => x113_out_4,
   I3 => W_22_19_i_12_n_0,
   I4 => W_22_19_i_13_n_0,
   O => W_22_19_i_3_n_0
);
W_22_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x113_out_26,
   I1 => x113_out_1,
   I2 => x113_out_3,
   I3 => W_22_19_i_14_n_0,
   I4 => W_22_19_i_15_n_0,
   O => W_22_19_i_4_n_0
);
W_22_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x113_out_25,
   I1 => x113_out_0,
   I2 => x113_out_2,
   I3 => W_22_19_i_16_n_0,
   I4 => W_22_19_i_17_n_0,
   O => W_22_19_i_5_n_0
);
W_22_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_22_19_i_2_n_0,
   I1 => W_22_23_i_16_n_0,
   I2 => x113_out_29,
   I3 => x113_out_4,
   I4 => x113_out_6,
   I5 => W_22_23_i_17_n_0,
   O => W_22_19_i_6_n_0
);
W_22_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_22_19_i_3_n_0,
   I1 => W_22_19_i_10_n_0,
   I2 => x113_out_28,
   I3 => x113_out_3,
   I4 => x113_out_5,
   I5 => W_22_19_i_11_n_0,
   O => W_22_19_i_7_n_0
);
W_22_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_22_19_i_4_n_0,
   I1 => W_22_19_i_12_n_0,
   I2 => x113_out_27,
   I3 => x113_out_2,
   I4 => x113_out_4,
   I5 => W_22_19_i_13_n_0,
   O => W_22_19_i_8_n_0
);
W_22_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_22_19_i_5_n_0,
   I1 => W_22_19_i_14_n_0,
   I2 => x113_out_26,
   I3 => x113_out_1,
   I4 => x113_out_3,
   I5 => W_22_19_i_15_n_0,
   O => W_22_19_i_9_n_0
);
W_22_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_6_22,
   I1 => M_reg_15_22,
   I2 => M_reg_7_8,
   I3 => M_reg_7_29,
   I4 => M_reg_7_25,
   O => W_22_23_i_10_n_0
);
W_22_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_15_21,
   I1 => M_reg_7_24,
   I2 => M_reg_7_28,
   I3 => M_reg_7_7,
   I4 => M_reg_6_21,
   O => W_22_23_i_11_n_0
);
W_22_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_6_21,
   I1 => M_reg_15_21,
   I2 => M_reg_7_7,
   I3 => M_reg_7_28,
   I4 => M_reg_7_24,
   O => W_22_23_i_12_n_0
);
W_22_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_15_20,
   I1 => M_reg_7_23,
   I2 => M_reg_7_27,
   I3 => M_reg_7_6,
   I4 => M_reg_6_20,
   O => W_22_23_i_13_n_0
);
W_22_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_6_20,
   I1 => M_reg_15_20,
   I2 => M_reg_7_6,
   I3 => M_reg_7_27,
   I4 => M_reg_7_23,
   O => W_22_23_i_14_n_0
);
W_22_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_15_19,
   I1 => M_reg_7_22,
   I2 => M_reg_7_26,
   I3 => M_reg_7_5,
   I4 => M_reg_6_19,
   O => W_22_23_i_15_n_0
);
W_22_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_6_19,
   I1 => M_reg_15_19,
   I2 => M_reg_7_5,
   I3 => M_reg_7_26,
   I4 => M_reg_7_22,
   O => W_22_23_i_16_n_0
);
W_22_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_15_18,
   I1 => M_reg_7_21,
   I2 => M_reg_7_25,
   I3 => M_reg_7_4,
   I4 => M_reg_6_18,
   O => W_22_23_i_17_n_0
);
W_22_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x113_out_7,
   I1 => x113_out_9,
   I2 => W_22_23_i_10_n_0,
   I3 => W_22_23_i_11_n_0,
   O => W_22_23_i_2_n_0
);
W_22_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x113_out_31,
   I1 => x113_out_6,
   I2 => x113_out_8,
   I3 => W_22_23_i_12_n_0,
   I4 => W_22_23_i_13_n_0,
   O => W_22_23_i_3_n_0
);
W_22_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x113_out_30,
   I1 => x113_out_5,
   I2 => x113_out_7,
   I3 => W_22_23_i_14_n_0,
   I4 => W_22_23_i_15_n_0,
   O => W_22_23_i_4_n_0
);
W_22_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x113_out_29,
   I1 => x113_out_4,
   I2 => x113_out_6,
   I3 => W_22_23_i_16_n_0,
   I4 => W_22_23_i_17_n_0,
   O => W_22_23_i_5_n_0
);
W_22_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x113_out_8,
   I1 => x113_out_10,
   I2 => W_22_27_i_16_n_0,
   I3 => W_22_27_i_17_n_0,
   I4 => W_22_23_i_2_n_0,
   O => W_22_23_i_6_n_0
);
W_22_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x113_out_7,
   I1 => x113_out_9,
   I2 => W_22_23_i_10_n_0,
   I3 => W_22_23_i_11_n_0,
   I4 => W_22_23_i_3_n_0,
   O => W_22_23_i_7_n_0
);
W_22_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_22_23_i_4_n_0,
   I1 => W_22_23_i_12_n_0,
   I2 => x113_out_31,
   I3 => x113_out_6,
   I4 => x113_out_8,
   I5 => W_22_23_i_13_n_0,
   O => W_22_23_i_8_n_0
);
W_22_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_22_23_i_5_n_0,
   I1 => W_22_23_i_14_n_0,
   I2 => x113_out_30,
   I3 => x113_out_5,
   I4 => x113_out_7,
   I5 => W_22_23_i_15_n_0,
   O => W_22_23_i_9_n_0
);
W_22_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_6_26,
   I1 => M_reg_15_26,
   I2 => M_reg_7_12,
   I3 => M_reg_7_1,
   I4 => M_reg_7_29,
   O => W_22_27_i_10_n_0
);
W_22_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_15_25,
   I1 => M_reg_7_28,
   I2 => M_reg_7_0,
   I3 => M_reg_7_11,
   I4 => M_reg_6_25,
   O => W_22_27_i_11_n_0
);
W_22_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_6_25,
   I1 => M_reg_15_25,
   I2 => M_reg_7_11,
   I3 => M_reg_7_0,
   I4 => M_reg_7_28,
   O => W_22_27_i_12_n_0
);
W_22_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_15_24,
   I1 => M_reg_7_27,
   I2 => M_reg_7_31,
   I3 => M_reg_7_10,
   I4 => M_reg_6_24,
   O => W_22_27_i_13_n_0
);
W_22_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_6_24,
   I1 => M_reg_15_24,
   I2 => M_reg_7_10,
   I3 => M_reg_7_31,
   I4 => M_reg_7_27,
   O => W_22_27_i_14_n_0
);
W_22_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_15_23,
   I1 => M_reg_7_26,
   I2 => M_reg_7_30,
   I3 => M_reg_7_9,
   I4 => M_reg_6_23,
   O => W_22_27_i_15_n_0
);
W_22_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_6_23,
   I1 => M_reg_15_23,
   I2 => M_reg_7_9,
   I3 => M_reg_7_30,
   I4 => M_reg_7_26,
   O => W_22_27_i_16_n_0
);
W_22_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_15_22,
   I1 => M_reg_7_25,
   I2 => M_reg_7_29,
   I3 => M_reg_7_8,
   I4 => M_reg_6_22,
   O => W_22_27_i_17_n_0
);
W_22_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x113_out_11,
   I1 => x113_out_13,
   I2 => W_22_27_i_10_n_0,
   I3 => W_22_27_i_11_n_0,
   O => W_22_27_i_2_n_0
);
W_22_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x113_out_10,
   I1 => x113_out_12,
   I2 => W_22_27_i_12_n_0,
   I3 => W_22_27_i_13_n_0,
   O => W_22_27_i_3_n_0
);
W_22_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x113_out_9,
   I1 => x113_out_11,
   I2 => W_22_27_i_14_n_0,
   I3 => W_22_27_i_15_n_0,
   O => W_22_27_i_4_n_0
);
W_22_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x113_out_8,
   I1 => x113_out_10,
   I2 => W_22_27_i_16_n_0,
   I3 => W_22_27_i_17_n_0,
   O => W_22_27_i_5_n_0
);
W_22_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x113_out_12,
   I1 => x113_out_14,
   I2 => W_22_31_i_13_n_0,
   I3 => W_22_31_i_14_n_0,
   I4 => W_22_27_i_2_n_0,
   O => W_22_27_i_6_n_0
);
W_22_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x113_out_11,
   I1 => x113_out_13,
   I2 => W_22_27_i_10_n_0,
   I3 => W_22_27_i_11_n_0,
   I4 => W_22_27_i_3_n_0,
   O => W_22_27_i_7_n_0
);
W_22_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x113_out_10,
   I1 => x113_out_12,
   I2 => W_22_27_i_12_n_0,
   I3 => W_22_27_i_13_n_0,
   I4 => W_22_27_i_4_n_0,
   O => W_22_27_i_8_n_0
);
W_22_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x113_out_9,
   I1 => x113_out_11,
   I2 => W_22_27_i_14_n_0,
   I3 => W_22_27_i_15_n_0,
   I4 => W_22_27_i_5_n_0,
   O => W_22_27_i_9_n_0
);
W_22_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_15_28,
   I1 => M_reg_7_31,
   I2 => M_reg_7_3,
   I3 => M_reg_7_14,
   I4 => M_reg_6_28,
   O => W_22_31_i_10_n_0
);
W_22_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_6_28,
   I1 => M_reg_15_28,
   I2 => M_reg_7_14,
   I3 => M_reg_7_3,
   I4 => M_reg_7_31,
   O => W_22_31_i_11_n_0
);
W_22_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_15_27,
   I1 => M_reg_7_30,
   I2 => M_reg_7_2,
   I3 => M_reg_7_13,
   I4 => M_reg_6_27,
   O => W_22_31_i_12_n_0
);
W_22_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_6_27,
   I1 => M_reg_15_27,
   I2 => M_reg_7_13,
   I3 => M_reg_7_2,
   I4 => M_reg_7_30,
   O => W_22_31_i_13_n_0
);
W_22_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_15_26,
   I1 => M_reg_7_29,
   I2 => M_reg_7_1,
   I3 => M_reg_7_12,
   I4 => M_reg_6_26,
   O => W_22_31_i_14_n_0
);
W_22_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => M_reg_15_29,
   I1 => M_reg_7_4,
   I2 => M_reg_7_15,
   I3 => M_reg_6_29,
   O => W_22_31_i_15_n_0
);
W_22_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x113_out_17,
   I1 => x113_out_15,
   O => SIGMA_LCASE_1339_out_30
);
W_22_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => M_reg_7_6,
   I1 => M_reg_7_17,
   I2 => M_reg_15_31,
   I3 => M_reg_6_31,
   I4 => x113_out_16,
   I5 => x113_out_18,
   O => W_22_31_i_17_n_0
);
W_22_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => M_reg_7_16,
   I1 => M_reg_7_5,
   O => SIGMA_LCASE_0335_out_30
);
W_22_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => M_reg_6_30,
   I1 => M_reg_15_30,
   I2 => M_reg_7_16,
   I3 => M_reg_7_5,
   O => W_22_31_i_19_n_0
);
W_22_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x113_out_14,
   I1 => x113_out_16,
   I2 => W_22_31_i_9_n_0,
   I3 => W_22_31_i_10_n_0,
   O => W_22_31_i_2_n_0
);
W_22_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x113_out_13,
   I1 => x113_out_15,
   I2 => W_22_31_i_11_n_0,
   I3 => W_22_31_i_12_n_0,
   O => W_22_31_i_3_n_0
);
W_22_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x113_out_12,
   I1 => x113_out_14,
   I2 => W_22_31_i_13_n_0,
   I3 => W_22_31_i_14_n_0,
   O => W_22_31_i_4_n_0
);
W_22_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_22_31_i_15_n_0,
   I1 => SIGMA_LCASE_1339_out_30,
   I2 => W_22_31_i_17_n_0,
   I3 => M_reg_15_30,
   I4 => SIGMA_LCASE_0335_out_30,
   I5 => M_reg_6_30,
   O => W_22_31_i_5_n_0
);
W_22_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_22_31_i_2_n_0,
   I1 => W_22_31_i_19_n_0,
   I2 => x113_out_15,
   I3 => x113_out_17,
   I4 => W_22_31_i_15_n_0,
   O => W_22_31_i_6_n_0
);
W_22_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x113_out_14,
   I1 => x113_out_16,
   I2 => W_22_31_i_9_n_0,
   I3 => W_22_31_i_10_n_0,
   I4 => W_22_31_i_3_n_0,
   O => W_22_31_i_7_n_0
);
W_22_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x113_out_13,
   I1 => x113_out_15,
   I2 => W_22_31_i_11_n_0,
   I3 => W_22_31_i_12_n_0,
   I4 => W_22_31_i_4_n_0,
   O => W_22_31_i_8_n_0
);
W_22_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => M_reg_6_29,
   I1 => M_reg_15_29,
   I2 => M_reg_7_15,
   I3 => M_reg_7_4,
   O => W_22_31_i_9_n_0
);
W_22_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_6_2,
   I1 => M_reg_15_2,
   I2 => M_reg_7_20,
   I3 => M_reg_7_9,
   I4 => M_reg_7_5,
   O => W_22_3_i_10_n_0
);
W_22_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_15_1,
   I1 => M_reg_7_4,
   I2 => M_reg_7_8,
   I3 => M_reg_7_19,
   I4 => M_reg_6_1,
   O => W_22_3_i_11_n_0
);
W_22_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => M_reg_7_19,
   I1 => M_reg_7_8,
   I2 => M_reg_7_4,
   O => SIGMA_LCASE_0335_out_1
);
W_22_3_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_6_1,
   I1 => M_reg_15_1,
   I2 => M_reg_7_19,
   I3 => M_reg_7_8,
   I4 => M_reg_7_4,
   O => W_22_3_i_13_n_0
);
W_22_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x113_out_12,
   I1 => x113_out_19,
   I2 => x113_out_21,
   I3 => W_22_3_i_10_n_0,
   I4 => W_22_3_i_11_n_0,
   O => W_22_3_i_2_n_0
);
W_22_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_22_3_i_11_n_0,
   I1 => x113_out_21,
   I2 => x113_out_19,
   I3 => x113_out_12,
   I4 => W_22_3_i_10_n_0,
   O => W_22_3_i_3_n_0
);
W_22_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_0335_out_1,
   I1 => M_reg_15_1,
   I2 => M_reg_6_1,
   I3 => x113_out_11,
   I4 => x113_out_18,
   I5 => x113_out_20,
   O => W_22_3_i_4_n_0
);
W_22_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_6_0,
   I1 => M_reg_15_0,
   I2 => M_reg_7_18,
   I3 => M_reg_7_7,
   I4 => M_reg_7_3,
   O => W_22_3_i_5_n_0
);
W_22_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_22_3_i_2_n_0,
   I1 => W_22_7_i_16_n_0,
   I2 => x113_out_13,
   I3 => x113_out_20,
   I4 => x113_out_22,
   I5 => W_22_7_i_17_n_0,
   O => W_22_3_i_6_n_0
);
W_22_3_i_7 : LUT5
  generic map(
   INIT => X"6aa6a66a"
  )
 port map (
   I0 => W_22_3_i_3_n_0,
   I1 => W_22_3_i_13_n_0,
   I2 => x113_out_20,
   I3 => x113_out_18,
   I4 => x113_out_11,
   O => W_22_3_i_7_n_0
);
W_22_3_i_8 : LUT6
  generic map(
   INIT => X"566565566aa6a66a"
  )
 port map (
   I0 => W_22_3_i_4_n_0,
   I1 => M_reg_6_0,
   I2 => M_reg_7_18,
   I3 => M_reg_7_7,
   I4 => M_reg_7_3,
   I5 => M_reg_15_0,
   O => W_22_3_i_8_n_0
);
W_22_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_22_3_i_5_n_0,
   I1 => x113_out_10,
   I2 => x113_out_17,
   I3 => x113_out_19,
   O => W_22_3_i_9_n_0
);
W_22_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_6_6,
   I1 => M_reg_15_6,
   I2 => M_reg_7_24,
   I3 => M_reg_7_13,
   I4 => M_reg_7_9,
   O => W_22_7_i_10_n_0
);
W_22_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_15_5,
   I1 => M_reg_7_8,
   I2 => M_reg_7_12,
   I3 => M_reg_7_23,
   I4 => M_reg_6_5,
   O => W_22_7_i_11_n_0
);
W_22_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_6_5,
   I1 => M_reg_15_5,
   I2 => M_reg_7_23,
   I3 => M_reg_7_12,
   I4 => M_reg_7_8,
   O => W_22_7_i_12_n_0
);
W_22_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_15_4,
   I1 => M_reg_7_7,
   I2 => M_reg_7_11,
   I3 => M_reg_7_22,
   I4 => M_reg_6_4,
   O => W_22_7_i_13_n_0
);
W_22_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_6_4,
   I1 => M_reg_15_4,
   I2 => M_reg_7_22,
   I3 => M_reg_7_11,
   I4 => M_reg_7_7,
   O => W_22_7_i_14_n_0
);
W_22_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_15_3,
   I1 => M_reg_7_6,
   I2 => M_reg_7_10,
   I3 => M_reg_7_21,
   I4 => M_reg_6_3,
   O => W_22_7_i_15_n_0
);
W_22_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_6_3,
   I1 => M_reg_15_3,
   I2 => M_reg_7_21,
   I3 => M_reg_7_10,
   I4 => M_reg_7_6,
   O => W_22_7_i_16_n_0
);
W_22_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => M_reg_15_2,
   I1 => M_reg_7_5,
   I2 => M_reg_7_9,
   I3 => M_reg_7_20,
   I4 => M_reg_6_2,
   O => W_22_7_i_17_n_0
);
W_22_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x113_out_16,
   I1 => x113_out_23,
   I2 => x113_out_25,
   I3 => W_22_7_i_10_n_0,
   I4 => W_22_7_i_11_n_0,
   O => W_22_7_i_2_n_0
);
W_22_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x113_out_15,
   I1 => x113_out_22,
   I2 => x113_out_24,
   I3 => W_22_7_i_12_n_0,
   I4 => W_22_7_i_13_n_0,
   O => W_22_7_i_3_n_0
);
W_22_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x113_out_14,
   I1 => x113_out_21,
   I2 => x113_out_23,
   I3 => W_22_7_i_14_n_0,
   I4 => W_22_7_i_15_n_0,
   O => W_22_7_i_4_n_0
);
W_22_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x113_out_13,
   I1 => x113_out_20,
   I2 => x113_out_22,
   I3 => W_22_7_i_16_n_0,
   I4 => W_22_7_i_17_n_0,
   O => W_22_7_i_5_n_0
);
W_22_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_22_7_i_2_n_0,
   I1 => W_22_11_i_16_n_0,
   I2 => x113_out_17,
   I3 => x113_out_24,
   I4 => x113_out_26,
   I5 => W_22_11_i_17_n_0,
   O => W_22_7_i_6_n_0
);
W_22_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_22_7_i_3_n_0,
   I1 => W_22_7_i_10_n_0,
   I2 => x113_out_16,
   I3 => x113_out_23,
   I4 => x113_out_25,
   I5 => W_22_7_i_11_n_0,
   O => W_22_7_i_7_n_0
);
W_22_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_22_7_i_4_n_0,
   I1 => W_22_7_i_12_n_0,
   I2 => x113_out_15,
   I3 => x113_out_22,
   I4 => x113_out_24,
   I5 => W_22_7_i_13_n_0,
   O => W_22_7_i_8_n_0
);
W_22_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_22_7_i_5_n_0,
   I1 => W_22_7_i_14_n_0,
   I2 => x113_out_14,
   I3 => x113_out_21,
   I4 => x113_out_23,
   I5 => W_22_7_i_15_n_0,
   O => W_22_7_i_9_n_0
);
W_23_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_7_10,
   I1 => x117_out_10,
   I2 => M_reg_8_28,
   I3 => M_reg_8_17,
   I4 => M_reg_8_13,
   O => W_23_11_i_10_n_0
);
W_23_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x117_out_9,
   I1 => M_reg_8_12,
   I2 => M_reg_8_16,
   I3 => M_reg_8_27,
   I4 => M_reg_7_9,
   O => W_23_11_i_11_n_0
);
W_23_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_7_9,
   I1 => x117_out_9,
   I2 => M_reg_8_27,
   I3 => M_reg_8_16,
   I4 => M_reg_8_12,
   O => W_23_11_i_12_n_0
);
W_23_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x117_out_8,
   I1 => M_reg_8_11,
   I2 => M_reg_8_15,
   I3 => M_reg_8_26,
   I4 => M_reg_7_8,
   O => W_23_11_i_13_n_0
);
W_23_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_7_8,
   I1 => x117_out_8,
   I2 => M_reg_8_26,
   I3 => M_reg_8_15,
   I4 => M_reg_8_11,
   O => W_23_11_i_14_n_0
);
W_23_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x117_out_7,
   I1 => M_reg_8_10,
   I2 => M_reg_8_14,
   I3 => M_reg_8_25,
   I4 => M_reg_7_7,
   O => W_23_11_i_15_n_0
);
W_23_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_7_7,
   I1 => x117_out_7,
   I2 => M_reg_8_25,
   I3 => M_reg_8_14,
   I4 => M_reg_8_10,
   O => W_23_11_i_16_n_0
);
W_23_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x117_out_6,
   I1 => M_reg_8_9,
   I2 => M_reg_8_13,
   I3 => M_reg_8_24,
   I4 => M_reg_7_6,
   O => W_23_11_i_17_n_0
);
W_23_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x112_out_20,
   I1 => x112_out_27,
   I2 => x112_out_29,
   I3 => W_23_11_i_10_n_0,
   I4 => W_23_11_i_11_n_0,
   O => W_23_11_i_2_n_0
);
W_23_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x112_out_19,
   I1 => x112_out_26,
   I2 => x112_out_28,
   I3 => W_23_11_i_12_n_0,
   I4 => W_23_11_i_13_n_0,
   O => W_23_11_i_3_n_0
);
W_23_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x112_out_18,
   I1 => x112_out_25,
   I2 => x112_out_27,
   I3 => W_23_11_i_14_n_0,
   I4 => W_23_11_i_15_n_0,
   O => W_23_11_i_4_n_0
);
W_23_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x112_out_17,
   I1 => x112_out_24,
   I2 => x112_out_26,
   I3 => W_23_11_i_16_n_0,
   I4 => W_23_11_i_17_n_0,
   O => W_23_11_i_5_n_0
);
W_23_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_23_11_i_2_n_0,
   I1 => W_23_15_i_16_n_0,
   I2 => x112_out_21,
   I3 => x112_out_28,
   I4 => x112_out_30,
   I5 => W_23_15_i_17_n_0,
   O => W_23_11_i_6_n_0
);
W_23_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_23_11_i_3_n_0,
   I1 => W_23_11_i_10_n_0,
   I2 => x112_out_20,
   I3 => x112_out_27,
   I4 => x112_out_29,
   I5 => W_23_11_i_11_n_0,
   O => W_23_11_i_7_n_0
);
W_23_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_23_11_i_4_n_0,
   I1 => W_23_11_i_12_n_0,
   I2 => x112_out_19,
   I3 => x112_out_26,
   I4 => x112_out_28,
   I5 => W_23_11_i_13_n_0,
   O => W_23_11_i_8_n_0
);
W_23_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_23_11_i_5_n_0,
   I1 => W_23_11_i_14_n_0,
   I2 => x112_out_18,
   I3 => x112_out_25,
   I4 => x112_out_27,
   I5 => W_23_11_i_15_n_0,
   O => W_23_11_i_9_n_0
);
W_23_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_7_14,
   I1 => x117_out_14,
   I2 => M_reg_8_0,
   I3 => M_reg_8_21,
   I4 => M_reg_8_17,
   O => W_23_15_i_10_n_0
);
W_23_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x117_out_13,
   I1 => M_reg_8_16,
   I2 => M_reg_8_20,
   I3 => M_reg_8_31,
   I4 => M_reg_7_13,
   O => W_23_15_i_11_n_0
);
W_23_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_7_13,
   I1 => x117_out_13,
   I2 => M_reg_8_31,
   I3 => M_reg_8_20,
   I4 => M_reg_8_16,
   O => W_23_15_i_12_n_0
);
W_23_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x117_out_12,
   I1 => M_reg_8_15,
   I2 => M_reg_8_19,
   I3 => M_reg_8_30,
   I4 => M_reg_7_12,
   O => W_23_15_i_13_n_0
);
W_23_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_7_12,
   I1 => x117_out_12,
   I2 => M_reg_8_30,
   I3 => M_reg_8_19,
   I4 => M_reg_8_15,
   O => W_23_15_i_14_n_0
);
W_23_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x117_out_11,
   I1 => M_reg_8_14,
   I2 => M_reg_8_18,
   I3 => M_reg_8_29,
   I4 => M_reg_7_11,
   O => W_23_15_i_15_n_0
);
W_23_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_7_11,
   I1 => x117_out_11,
   I2 => M_reg_8_29,
   I3 => M_reg_8_18,
   I4 => M_reg_8_14,
   O => W_23_15_i_16_n_0
);
W_23_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x117_out_10,
   I1 => M_reg_8_13,
   I2 => M_reg_8_17,
   I3 => M_reg_8_28,
   I4 => M_reg_7_10,
   O => W_23_15_i_17_n_0
);
W_23_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x112_out_24,
   I1 => x112_out_31,
   I2 => x112_out_1,
   I3 => W_23_15_i_10_n_0,
   I4 => W_23_15_i_11_n_0,
   O => W_23_15_i_2_n_0
);
W_23_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x112_out_23,
   I1 => x112_out_30,
   I2 => x112_out_0,
   I3 => W_23_15_i_12_n_0,
   I4 => W_23_15_i_13_n_0,
   O => W_23_15_i_3_n_0
);
W_23_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x112_out_22,
   I1 => x112_out_29,
   I2 => x112_out_31,
   I3 => W_23_15_i_14_n_0,
   I4 => W_23_15_i_15_n_0,
   O => W_23_15_i_4_n_0
);
W_23_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x112_out_21,
   I1 => x112_out_28,
   I2 => x112_out_30,
   I3 => W_23_15_i_16_n_0,
   I4 => W_23_15_i_17_n_0,
   O => W_23_15_i_5_n_0
);
W_23_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_23_15_i_2_n_0,
   I1 => W_23_19_i_16_n_0,
   I2 => x112_out_25,
   I3 => x112_out_0,
   I4 => x112_out_2,
   I5 => W_23_19_i_17_n_0,
   O => W_23_15_i_6_n_0
);
W_23_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_23_15_i_3_n_0,
   I1 => W_23_15_i_10_n_0,
   I2 => x112_out_24,
   I3 => x112_out_31,
   I4 => x112_out_1,
   I5 => W_23_15_i_11_n_0,
   O => W_23_15_i_7_n_0
);
W_23_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_23_15_i_4_n_0,
   I1 => W_23_15_i_12_n_0,
   I2 => x112_out_23,
   I3 => x112_out_30,
   I4 => x112_out_0,
   I5 => W_23_15_i_13_n_0,
   O => W_23_15_i_8_n_0
);
W_23_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_23_15_i_5_n_0,
   I1 => W_23_15_i_14_n_0,
   I2 => x112_out_22,
   I3 => x112_out_29,
   I4 => x112_out_31,
   I5 => W_23_15_i_15_n_0,
   O => W_23_15_i_9_n_0
);
W_23_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_7_18,
   I1 => x117_out_18,
   I2 => M_reg_8_4,
   I3 => M_reg_8_25,
   I4 => M_reg_8_21,
   O => W_23_19_i_10_n_0
);
W_23_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x117_out_17,
   I1 => M_reg_8_20,
   I2 => M_reg_8_24,
   I3 => M_reg_8_3,
   I4 => M_reg_7_17,
   O => W_23_19_i_11_n_0
);
W_23_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_7_17,
   I1 => x117_out_17,
   I2 => M_reg_8_3,
   I3 => M_reg_8_24,
   I4 => M_reg_8_20,
   O => W_23_19_i_12_n_0
);
W_23_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x117_out_16,
   I1 => M_reg_8_19,
   I2 => M_reg_8_23,
   I3 => M_reg_8_2,
   I4 => M_reg_7_16,
   O => W_23_19_i_13_n_0
);
W_23_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_7_16,
   I1 => x117_out_16,
   I2 => M_reg_8_2,
   I3 => M_reg_8_23,
   I4 => M_reg_8_19,
   O => W_23_19_i_14_n_0
);
W_23_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x117_out_15,
   I1 => M_reg_8_18,
   I2 => M_reg_8_22,
   I3 => M_reg_8_1,
   I4 => M_reg_7_15,
   O => W_23_19_i_15_n_0
);
W_23_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_7_15,
   I1 => x117_out_15,
   I2 => M_reg_8_1,
   I3 => M_reg_8_22,
   I4 => M_reg_8_18,
   O => W_23_19_i_16_n_0
);
W_23_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x117_out_14,
   I1 => M_reg_8_17,
   I2 => M_reg_8_21,
   I3 => M_reg_8_0,
   I4 => M_reg_7_14,
   O => W_23_19_i_17_n_0
);
W_23_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x112_out_28,
   I1 => x112_out_3,
   I2 => x112_out_5,
   I3 => W_23_19_i_10_n_0,
   I4 => W_23_19_i_11_n_0,
   O => W_23_19_i_2_n_0
);
W_23_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x112_out_27,
   I1 => x112_out_2,
   I2 => x112_out_4,
   I3 => W_23_19_i_12_n_0,
   I4 => W_23_19_i_13_n_0,
   O => W_23_19_i_3_n_0
);
W_23_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x112_out_26,
   I1 => x112_out_1,
   I2 => x112_out_3,
   I3 => W_23_19_i_14_n_0,
   I4 => W_23_19_i_15_n_0,
   O => W_23_19_i_4_n_0
);
W_23_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x112_out_25,
   I1 => x112_out_0,
   I2 => x112_out_2,
   I3 => W_23_19_i_16_n_0,
   I4 => W_23_19_i_17_n_0,
   O => W_23_19_i_5_n_0
);
W_23_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_23_19_i_2_n_0,
   I1 => W_23_23_i_16_n_0,
   I2 => x112_out_29,
   I3 => x112_out_4,
   I4 => x112_out_6,
   I5 => W_23_23_i_17_n_0,
   O => W_23_19_i_6_n_0
);
W_23_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_23_19_i_3_n_0,
   I1 => W_23_19_i_10_n_0,
   I2 => x112_out_28,
   I3 => x112_out_3,
   I4 => x112_out_5,
   I5 => W_23_19_i_11_n_0,
   O => W_23_19_i_7_n_0
);
W_23_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_23_19_i_4_n_0,
   I1 => W_23_19_i_12_n_0,
   I2 => x112_out_27,
   I3 => x112_out_2,
   I4 => x112_out_4,
   I5 => W_23_19_i_13_n_0,
   O => W_23_19_i_8_n_0
);
W_23_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_23_19_i_5_n_0,
   I1 => W_23_19_i_14_n_0,
   I2 => x112_out_26,
   I3 => x112_out_1,
   I4 => x112_out_3,
   I5 => W_23_19_i_15_n_0,
   O => W_23_19_i_9_n_0
);
W_23_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_7_22,
   I1 => x117_out_22,
   I2 => M_reg_8_8,
   I3 => M_reg_8_29,
   I4 => M_reg_8_25,
   O => W_23_23_i_10_n_0
);
W_23_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x117_out_21,
   I1 => M_reg_8_24,
   I2 => M_reg_8_28,
   I3 => M_reg_8_7,
   I4 => M_reg_7_21,
   O => W_23_23_i_11_n_0
);
W_23_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_7_21,
   I1 => x117_out_21,
   I2 => M_reg_8_7,
   I3 => M_reg_8_28,
   I4 => M_reg_8_24,
   O => W_23_23_i_12_n_0
);
W_23_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x117_out_20,
   I1 => M_reg_8_23,
   I2 => M_reg_8_27,
   I3 => M_reg_8_6,
   I4 => M_reg_7_20,
   O => W_23_23_i_13_n_0
);
W_23_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_7_20,
   I1 => x117_out_20,
   I2 => M_reg_8_6,
   I3 => M_reg_8_27,
   I4 => M_reg_8_23,
   O => W_23_23_i_14_n_0
);
W_23_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x117_out_19,
   I1 => M_reg_8_22,
   I2 => M_reg_8_26,
   I3 => M_reg_8_5,
   I4 => M_reg_7_19,
   O => W_23_23_i_15_n_0
);
W_23_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_7_19,
   I1 => x117_out_19,
   I2 => M_reg_8_5,
   I3 => M_reg_8_26,
   I4 => M_reg_8_22,
   O => W_23_23_i_16_n_0
);
W_23_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x117_out_18,
   I1 => M_reg_8_21,
   I2 => M_reg_8_25,
   I3 => M_reg_8_4,
   I4 => M_reg_7_18,
   O => W_23_23_i_17_n_0
);
W_23_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x112_out_7,
   I1 => x112_out_9,
   I2 => W_23_23_i_10_n_0,
   I3 => W_23_23_i_11_n_0,
   O => W_23_23_i_2_n_0
);
W_23_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x112_out_31,
   I1 => x112_out_6,
   I2 => x112_out_8,
   I3 => W_23_23_i_12_n_0,
   I4 => W_23_23_i_13_n_0,
   O => W_23_23_i_3_n_0
);
W_23_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x112_out_30,
   I1 => x112_out_5,
   I2 => x112_out_7,
   I3 => W_23_23_i_14_n_0,
   I4 => W_23_23_i_15_n_0,
   O => W_23_23_i_4_n_0
);
W_23_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x112_out_29,
   I1 => x112_out_4,
   I2 => x112_out_6,
   I3 => W_23_23_i_16_n_0,
   I4 => W_23_23_i_17_n_0,
   O => W_23_23_i_5_n_0
);
W_23_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x112_out_8,
   I1 => x112_out_10,
   I2 => W_23_27_i_16_n_0,
   I3 => W_23_27_i_17_n_0,
   I4 => W_23_23_i_2_n_0,
   O => W_23_23_i_6_n_0
);
W_23_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x112_out_7,
   I1 => x112_out_9,
   I2 => W_23_23_i_10_n_0,
   I3 => W_23_23_i_11_n_0,
   I4 => W_23_23_i_3_n_0,
   O => W_23_23_i_7_n_0
);
W_23_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_23_23_i_4_n_0,
   I1 => W_23_23_i_12_n_0,
   I2 => x112_out_31,
   I3 => x112_out_6,
   I4 => x112_out_8,
   I5 => W_23_23_i_13_n_0,
   O => W_23_23_i_8_n_0
);
W_23_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_23_23_i_5_n_0,
   I1 => W_23_23_i_14_n_0,
   I2 => x112_out_30,
   I3 => x112_out_5,
   I4 => x112_out_7,
   I5 => W_23_23_i_15_n_0,
   O => W_23_23_i_9_n_0
);
W_23_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_7_26,
   I1 => x117_out_26,
   I2 => M_reg_8_12,
   I3 => M_reg_8_1,
   I4 => M_reg_8_29,
   O => W_23_27_i_10_n_0
);
W_23_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x117_out_25,
   I1 => M_reg_8_28,
   I2 => M_reg_8_0,
   I3 => M_reg_8_11,
   I4 => M_reg_7_25,
   O => W_23_27_i_11_n_0
);
W_23_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_7_25,
   I1 => x117_out_25,
   I2 => M_reg_8_11,
   I3 => M_reg_8_0,
   I4 => M_reg_8_28,
   O => W_23_27_i_12_n_0
);
W_23_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x117_out_24,
   I1 => M_reg_8_27,
   I2 => M_reg_8_31,
   I3 => M_reg_8_10,
   I4 => M_reg_7_24,
   O => W_23_27_i_13_n_0
);
W_23_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_7_24,
   I1 => x117_out_24,
   I2 => M_reg_8_10,
   I3 => M_reg_8_31,
   I4 => M_reg_8_27,
   O => W_23_27_i_14_n_0
);
W_23_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x117_out_23,
   I1 => M_reg_8_26,
   I2 => M_reg_8_30,
   I3 => M_reg_8_9,
   I4 => M_reg_7_23,
   O => W_23_27_i_15_n_0
);
W_23_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_7_23,
   I1 => x117_out_23,
   I2 => M_reg_8_9,
   I3 => M_reg_8_30,
   I4 => M_reg_8_26,
   O => W_23_27_i_16_n_0
);
W_23_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x117_out_22,
   I1 => M_reg_8_25,
   I2 => M_reg_8_29,
   I3 => M_reg_8_8,
   I4 => M_reg_7_22,
   O => W_23_27_i_17_n_0
);
W_23_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x112_out_11,
   I1 => x112_out_13,
   I2 => W_23_27_i_10_n_0,
   I3 => W_23_27_i_11_n_0,
   O => W_23_27_i_2_n_0
);
W_23_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x112_out_10,
   I1 => x112_out_12,
   I2 => W_23_27_i_12_n_0,
   I3 => W_23_27_i_13_n_0,
   O => W_23_27_i_3_n_0
);
W_23_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x112_out_9,
   I1 => x112_out_11,
   I2 => W_23_27_i_14_n_0,
   I3 => W_23_27_i_15_n_0,
   O => W_23_27_i_4_n_0
);
W_23_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x112_out_8,
   I1 => x112_out_10,
   I2 => W_23_27_i_16_n_0,
   I3 => W_23_27_i_17_n_0,
   O => W_23_27_i_5_n_0
);
W_23_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x112_out_12,
   I1 => x112_out_14,
   I2 => W_23_31_i_13_n_0,
   I3 => W_23_31_i_14_n_0,
   I4 => W_23_27_i_2_n_0,
   O => W_23_27_i_6_n_0
);
W_23_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x112_out_11,
   I1 => x112_out_13,
   I2 => W_23_27_i_10_n_0,
   I3 => W_23_27_i_11_n_0,
   I4 => W_23_27_i_3_n_0,
   O => W_23_27_i_7_n_0
);
W_23_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x112_out_10,
   I1 => x112_out_12,
   I2 => W_23_27_i_12_n_0,
   I3 => W_23_27_i_13_n_0,
   I4 => W_23_27_i_4_n_0,
   O => W_23_27_i_8_n_0
);
W_23_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x112_out_9,
   I1 => x112_out_11,
   I2 => W_23_27_i_14_n_0,
   I3 => W_23_27_i_15_n_0,
   I4 => W_23_27_i_5_n_0,
   O => W_23_27_i_9_n_0
);
W_23_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x117_out_28,
   I1 => M_reg_8_31,
   I2 => M_reg_8_3,
   I3 => M_reg_8_14,
   I4 => M_reg_7_28,
   O => W_23_31_i_10_n_0
);
W_23_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_7_28,
   I1 => x117_out_28,
   I2 => M_reg_8_14,
   I3 => M_reg_8_3,
   I4 => M_reg_8_31,
   O => W_23_31_i_11_n_0
);
W_23_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x117_out_27,
   I1 => M_reg_8_30,
   I2 => M_reg_8_2,
   I3 => M_reg_8_13,
   I4 => M_reg_7_27,
   O => W_23_31_i_12_n_0
);
W_23_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_7_27,
   I1 => x117_out_27,
   I2 => M_reg_8_13,
   I3 => M_reg_8_2,
   I4 => M_reg_8_30,
   O => W_23_31_i_13_n_0
);
W_23_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x117_out_26,
   I1 => M_reg_8_29,
   I2 => M_reg_8_1,
   I3 => M_reg_8_12,
   I4 => M_reg_7_26,
   O => W_23_31_i_14_n_0
);
W_23_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x117_out_29,
   I1 => M_reg_8_4,
   I2 => M_reg_8_15,
   I3 => M_reg_7_29,
   O => W_23_31_i_15_n_0
);
W_23_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x112_out_17,
   I1 => x112_out_15,
   O => SIGMA_LCASE_1331_out_0_30
);
W_23_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => M_reg_8_6,
   I1 => M_reg_8_17,
   I2 => x117_out_31,
   I3 => M_reg_7_31,
   I4 => x112_out_16,
   I5 => x112_out_18,
   O => W_23_31_i_17_n_0
);
W_23_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => M_reg_8_16,
   I1 => M_reg_8_5,
   O => SIGMA_LCASE_0327_out_30
);
W_23_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => M_reg_7_30,
   I1 => x117_out_30,
   I2 => M_reg_8_16,
   I3 => M_reg_8_5,
   O => W_23_31_i_19_n_0
);
W_23_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x112_out_14,
   I1 => x112_out_16,
   I2 => W_23_31_i_9_n_0,
   I3 => W_23_31_i_10_n_0,
   O => W_23_31_i_2_n_0
);
W_23_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x112_out_13,
   I1 => x112_out_15,
   I2 => W_23_31_i_11_n_0,
   I3 => W_23_31_i_12_n_0,
   O => W_23_31_i_3_n_0
);
W_23_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x112_out_12,
   I1 => x112_out_14,
   I2 => W_23_31_i_13_n_0,
   I3 => W_23_31_i_14_n_0,
   O => W_23_31_i_4_n_0
);
W_23_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_23_31_i_15_n_0,
   I1 => SIGMA_LCASE_1331_out_0_30,
   I2 => W_23_31_i_17_n_0,
   I3 => x117_out_30,
   I4 => SIGMA_LCASE_0327_out_30,
   I5 => M_reg_7_30,
   O => W_23_31_i_5_n_0
);
W_23_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_23_31_i_2_n_0,
   I1 => W_23_31_i_19_n_0,
   I2 => x112_out_15,
   I3 => x112_out_17,
   I4 => W_23_31_i_15_n_0,
   O => W_23_31_i_6_n_0
);
W_23_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x112_out_14,
   I1 => x112_out_16,
   I2 => W_23_31_i_9_n_0,
   I3 => W_23_31_i_10_n_0,
   I4 => W_23_31_i_3_n_0,
   O => W_23_31_i_7_n_0
);
W_23_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x112_out_13,
   I1 => x112_out_15,
   I2 => W_23_31_i_11_n_0,
   I3 => W_23_31_i_12_n_0,
   I4 => W_23_31_i_4_n_0,
   O => W_23_31_i_8_n_0
);
W_23_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => M_reg_7_29,
   I1 => x117_out_29,
   I2 => M_reg_8_15,
   I3 => M_reg_8_4,
   O => W_23_31_i_9_n_0
);
W_23_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_7_2,
   I1 => x117_out_2,
   I2 => M_reg_8_20,
   I3 => M_reg_8_9,
   I4 => M_reg_8_5,
   O => W_23_3_i_10_n_0
);
W_23_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x117_out_1,
   I1 => M_reg_8_4,
   I2 => M_reg_8_8,
   I3 => M_reg_8_19,
   I4 => M_reg_7_1,
   O => W_23_3_i_11_n_0
);
W_23_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => M_reg_8_19,
   I1 => M_reg_8_8,
   I2 => M_reg_8_4,
   O => SIGMA_LCASE_0327_out_1
);
W_23_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x112_out_21,
   I1 => x112_out_19,
   I2 => x112_out_12,
   O => SIGMA_LCASE_1331_out_0_2
);
W_23_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x112_out_20,
   I1 => x112_out_18,
   I2 => x112_out_11,
   O => SIGMA_LCASE_1331_out_1
);
W_23_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x112_out_12,
   I1 => x112_out_19,
   I2 => x112_out_21,
   I3 => W_23_3_i_10_n_0,
   I4 => W_23_3_i_11_n_0,
   O => W_23_3_i_2_n_0
);
W_23_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_23_3_i_11_n_0,
   I1 => x112_out_21,
   I2 => x112_out_19,
   I3 => x112_out_12,
   I4 => W_23_3_i_10_n_0,
   O => W_23_3_i_3_n_0
);
W_23_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_0327_out_1,
   I1 => x117_out_1,
   I2 => M_reg_7_1,
   I3 => x112_out_11,
   I4 => x112_out_18,
   I5 => x112_out_20,
   O => W_23_3_i_4_n_0
);
W_23_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_7_0,
   I1 => x117_out_0,
   I2 => M_reg_8_18,
   I3 => M_reg_8_7,
   I4 => M_reg_8_3,
   O => W_23_3_i_5_n_0
);
W_23_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_23_3_i_2_n_0,
   I1 => W_23_7_i_16_n_0,
   I2 => x112_out_13,
   I3 => x112_out_20,
   I4 => x112_out_22,
   I5 => W_23_7_i_17_n_0,
   O => W_23_3_i_6_n_0
);
W_23_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_23_3_i_10_n_0,
   I1 => SIGMA_LCASE_1331_out_0_2,
   I2 => M_reg_7_1,
   I3 => x117_out_1,
   I4 => SIGMA_LCASE_0327_out_1,
   I5 => SIGMA_LCASE_1331_out_1,
   O => W_23_3_i_7_n_0
);
W_23_3_i_8 : LUT6
  generic map(
   INIT => X"566565566aa6a66a"
  )
 port map (
   I0 => W_23_3_i_4_n_0,
   I1 => M_reg_7_0,
   I2 => M_reg_8_18,
   I3 => M_reg_8_7,
   I4 => M_reg_8_3,
   I5 => x117_out_0,
   O => W_23_3_i_8_n_0
);
W_23_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_23_3_i_5_n_0,
   I1 => x112_out_10,
   I2 => x112_out_17,
   I3 => x112_out_19,
   O => W_23_3_i_9_n_0
);
W_23_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_7_6,
   I1 => x117_out_6,
   I2 => M_reg_8_24,
   I3 => M_reg_8_13,
   I4 => M_reg_8_9,
   O => W_23_7_i_10_n_0
);
W_23_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x117_out_5,
   I1 => M_reg_8_8,
   I2 => M_reg_8_12,
   I3 => M_reg_8_23,
   I4 => M_reg_7_5,
   O => W_23_7_i_11_n_0
);
W_23_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_7_5,
   I1 => x117_out_5,
   I2 => M_reg_8_23,
   I3 => M_reg_8_12,
   I4 => M_reg_8_8,
   O => W_23_7_i_12_n_0
);
W_23_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x117_out_4,
   I1 => M_reg_8_7,
   I2 => M_reg_8_11,
   I3 => M_reg_8_22,
   I4 => M_reg_7_4,
   O => W_23_7_i_13_n_0
);
W_23_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_7_4,
   I1 => x117_out_4,
   I2 => M_reg_8_22,
   I3 => M_reg_8_11,
   I4 => M_reg_8_7,
   O => W_23_7_i_14_n_0
);
W_23_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x117_out_3,
   I1 => M_reg_8_6,
   I2 => M_reg_8_10,
   I3 => M_reg_8_21,
   I4 => M_reg_7_3,
   O => W_23_7_i_15_n_0
);
W_23_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_7_3,
   I1 => x117_out_3,
   I2 => M_reg_8_21,
   I3 => M_reg_8_10,
   I4 => M_reg_8_6,
   O => W_23_7_i_16_n_0
);
W_23_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x117_out_2,
   I1 => M_reg_8_5,
   I2 => M_reg_8_9,
   I3 => M_reg_8_20,
   I4 => M_reg_7_2,
   O => W_23_7_i_17_n_0
);
W_23_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x112_out_16,
   I1 => x112_out_23,
   I2 => x112_out_25,
   I3 => W_23_7_i_10_n_0,
   I4 => W_23_7_i_11_n_0,
   O => W_23_7_i_2_n_0
);
W_23_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x112_out_15,
   I1 => x112_out_22,
   I2 => x112_out_24,
   I3 => W_23_7_i_12_n_0,
   I4 => W_23_7_i_13_n_0,
   O => W_23_7_i_3_n_0
);
W_23_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x112_out_14,
   I1 => x112_out_21,
   I2 => x112_out_23,
   I3 => W_23_7_i_14_n_0,
   I4 => W_23_7_i_15_n_0,
   O => W_23_7_i_4_n_0
);
W_23_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x112_out_13,
   I1 => x112_out_20,
   I2 => x112_out_22,
   I3 => W_23_7_i_16_n_0,
   I4 => W_23_7_i_17_n_0,
   O => W_23_7_i_5_n_0
);
W_23_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_23_7_i_2_n_0,
   I1 => W_23_11_i_16_n_0,
   I2 => x112_out_17,
   I3 => x112_out_24,
   I4 => x112_out_26,
   I5 => W_23_11_i_17_n_0,
   O => W_23_7_i_6_n_0
);
W_23_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_23_7_i_3_n_0,
   I1 => W_23_7_i_10_n_0,
   I2 => x112_out_16,
   I3 => x112_out_23,
   I4 => x112_out_25,
   I5 => W_23_7_i_11_n_0,
   O => W_23_7_i_7_n_0
);
W_23_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_23_7_i_4_n_0,
   I1 => W_23_7_i_12_n_0,
   I2 => x112_out_15,
   I3 => x112_out_22,
   I4 => x112_out_24,
   I5 => W_23_7_i_13_n_0,
   O => W_23_7_i_8_n_0
);
W_23_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_23_7_i_5_n_0,
   I1 => W_23_7_i_14_n_0,
   I2 => x112_out_14,
   I3 => x112_out_21,
   I4 => x112_out_23,
   I5 => W_23_7_i_15_n_0,
   O => W_23_7_i_9_n_0
);
W_24_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_8_10,
   I1 => x116_out_10,
   I2 => M_reg_9_28,
   I3 => M_reg_9_17,
   I4 => M_reg_9_13,
   O => W_24_11_i_10_n_0
);
W_24_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x116_out_9,
   I1 => M_reg_9_12,
   I2 => M_reg_9_16,
   I3 => M_reg_9_27,
   I4 => M_reg_8_9,
   O => W_24_11_i_11_n_0
);
W_24_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_8_9,
   I1 => x116_out_9,
   I2 => M_reg_9_27,
   I3 => M_reg_9_16,
   I4 => M_reg_9_12,
   O => W_24_11_i_12_n_0
);
W_24_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x116_out_8,
   I1 => M_reg_9_11,
   I2 => M_reg_9_15,
   I3 => M_reg_9_26,
   I4 => M_reg_8_8,
   O => W_24_11_i_13_n_0
);
W_24_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_8_8,
   I1 => x116_out_8,
   I2 => M_reg_9_26,
   I3 => M_reg_9_15,
   I4 => M_reg_9_11,
   O => W_24_11_i_14_n_0
);
W_24_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x116_out_7,
   I1 => M_reg_9_10,
   I2 => M_reg_9_14,
   I3 => M_reg_9_25,
   I4 => M_reg_8_7,
   O => W_24_11_i_15_n_0
);
W_24_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_8_7,
   I1 => x116_out_7,
   I2 => M_reg_9_25,
   I3 => M_reg_9_14,
   I4 => M_reg_9_10,
   O => W_24_11_i_16_n_0
);
W_24_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x116_out_6,
   I1 => M_reg_9_9,
   I2 => M_reg_9_13,
   I3 => M_reg_9_24,
   I4 => M_reg_8_6,
   O => W_24_11_i_17_n_0
);
W_24_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x111_out_20,
   I1 => x111_out_27,
   I2 => x111_out_29,
   I3 => W_24_11_i_10_n_0,
   I4 => W_24_11_i_11_n_0,
   O => W_24_11_i_2_n_0
);
W_24_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x111_out_19,
   I1 => x111_out_26,
   I2 => x111_out_28,
   I3 => W_24_11_i_12_n_0,
   I4 => W_24_11_i_13_n_0,
   O => W_24_11_i_3_n_0
);
W_24_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x111_out_18,
   I1 => x111_out_25,
   I2 => x111_out_27,
   I3 => W_24_11_i_14_n_0,
   I4 => W_24_11_i_15_n_0,
   O => W_24_11_i_4_n_0
);
W_24_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x111_out_17,
   I1 => x111_out_24,
   I2 => x111_out_26,
   I3 => W_24_11_i_16_n_0,
   I4 => W_24_11_i_17_n_0,
   O => W_24_11_i_5_n_0
);
W_24_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_24_11_i_2_n_0,
   I1 => W_24_15_i_16_n_0,
   I2 => x111_out_21,
   I3 => x111_out_28,
   I4 => x111_out_30,
   I5 => W_24_15_i_17_n_0,
   O => W_24_11_i_6_n_0
);
W_24_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_24_11_i_3_n_0,
   I1 => W_24_11_i_10_n_0,
   I2 => x111_out_20,
   I3 => x111_out_27,
   I4 => x111_out_29,
   I5 => W_24_11_i_11_n_0,
   O => W_24_11_i_7_n_0
);
W_24_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_24_11_i_4_n_0,
   I1 => W_24_11_i_12_n_0,
   I2 => x111_out_19,
   I3 => x111_out_26,
   I4 => x111_out_28,
   I5 => W_24_11_i_13_n_0,
   O => W_24_11_i_8_n_0
);
W_24_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_24_11_i_5_n_0,
   I1 => W_24_11_i_14_n_0,
   I2 => x111_out_18,
   I3 => x111_out_25,
   I4 => x111_out_27,
   I5 => W_24_11_i_15_n_0,
   O => W_24_11_i_9_n_0
);
W_24_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_8_14,
   I1 => x116_out_14,
   I2 => M_reg_9_0,
   I3 => M_reg_9_21,
   I4 => M_reg_9_17,
   O => W_24_15_i_10_n_0
);
W_24_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x116_out_13,
   I1 => M_reg_9_16,
   I2 => M_reg_9_20,
   I3 => M_reg_9_31,
   I4 => M_reg_8_13,
   O => W_24_15_i_11_n_0
);
W_24_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_8_13,
   I1 => x116_out_13,
   I2 => M_reg_9_31,
   I3 => M_reg_9_20,
   I4 => M_reg_9_16,
   O => W_24_15_i_12_n_0
);
W_24_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x116_out_12,
   I1 => M_reg_9_15,
   I2 => M_reg_9_19,
   I3 => M_reg_9_30,
   I4 => M_reg_8_12,
   O => W_24_15_i_13_n_0
);
W_24_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_8_12,
   I1 => x116_out_12,
   I2 => M_reg_9_30,
   I3 => M_reg_9_19,
   I4 => M_reg_9_15,
   O => W_24_15_i_14_n_0
);
W_24_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x116_out_11,
   I1 => M_reg_9_14,
   I2 => M_reg_9_18,
   I3 => M_reg_9_29,
   I4 => M_reg_8_11,
   O => W_24_15_i_15_n_0
);
W_24_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_8_11,
   I1 => x116_out_11,
   I2 => M_reg_9_29,
   I3 => M_reg_9_18,
   I4 => M_reg_9_14,
   O => W_24_15_i_16_n_0
);
W_24_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x116_out_10,
   I1 => M_reg_9_13,
   I2 => M_reg_9_17,
   I3 => M_reg_9_28,
   I4 => M_reg_8_10,
   O => W_24_15_i_17_n_0
);
W_24_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x111_out_24,
   I1 => x111_out_31,
   I2 => x111_out_1,
   I3 => W_24_15_i_10_n_0,
   I4 => W_24_15_i_11_n_0,
   O => W_24_15_i_2_n_0
);
W_24_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x111_out_23,
   I1 => x111_out_30,
   I2 => x111_out_0,
   I3 => W_24_15_i_12_n_0,
   I4 => W_24_15_i_13_n_0,
   O => W_24_15_i_3_n_0
);
W_24_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x111_out_22,
   I1 => x111_out_29,
   I2 => x111_out_31,
   I3 => W_24_15_i_14_n_0,
   I4 => W_24_15_i_15_n_0,
   O => W_24_15_i_4_n_0
);
W_24_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x111_out_21,
   I1 => x111_out_28,
   I2 => x111_out_30,
   I3 => W_24_15_i_16_n_0,
   I4 => W_24_15_i_17_n_0,
   O => W_24_15_i_5_n_0
);
W_24_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_24_15_i_2_n_0,
   I1 => W_24_19_i_16_n_0,
   I2 => x111_out_25,
   I3 => x111_out_0,
   I4 => x111_out_2,
   I5 => W_24_19_i_17_n_0,
   O => W_24_15_i_6_n_0
);
W_24_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_24_15_i_3_n_0,
   I1 => W_24_15_i_10_n_0,
   I2 => x111_out_24,
   I3 => x111_out_31,
   I4 => x111_out_1,
   I5 => W_24_15_i_11_n_0,
   O => W_24_15_i_7_n_0
);
W_24_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_24_15_i_4_n_0,
   I1 => W_24_15_i_12_n_0,
   I2 => x111_out_23,
   I3 => x111_out_30,
   I4 => x111_out_0,
   I5 => W_24_15_i_13_n_0,
   O => W_24_15_i_8_n_0
);
W_24_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_24_15_i_5_n_0,
   I1 => W_24_15_i_14_n_0,
   I2 => x111_out_22,
   I3 => x111_out_29,
   I4 => x111_out_31,
   I5 => W_24_15_i_15_n_0,
   O => W_24_15_i_9_n_0
);
W_24_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_8_18,
   I1 => x116_out_18,
   I2 => M_reg_9_4,
   I3 => M_reg_9_25,
   I4 => M_reg_9_21,
   O => W_24_19_i_10_n_0
);
W_24_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x116_out_17,
   I1 => M_reg_9_20,
   I2 => M_reg_9_24,
   I3 => M_reg_9_3,
   I4 => M_reg_8_17,
   O => W_24_19_i_11_n_0
);
W_24_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_8_17,
   I1 => x116_out_17,
   I2 => M_reg_9_3,
   I3 => M_reg_9_24,
   I4 => M_reg_9_20,
   O => W_24_19_i_12_n_0
);
W_24_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x116_out_16,
   I1 => M_reg_9_19,
   I2 => M_reg_9_23,
   I3 => M_reg_9_2,
   I4 => M_reg_8_16,
   O => W_24_19_i_13_n_0
);
W_24_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_8_16,
   I1 => x116_out_16,
   I2 => M_reg_9_2,
   I3 => M_reg_9_23,
   I4 => M_reg_9_19,
   O => W_24_19_i_14_n_0
);
W_24_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x116_out_15,
   I1 => M_reg_9_18,
   I2 => M_reg_9_22,
   I3 => M_reg_9_1,
   I4 => M_reg_8_15,
   O => W_24_19_i_15_n_0
);
W_24_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_8_15,
   I1 => x116_out_15,
   I2 => M_reg_9_1,
   I3 => M_reg_9_22,
   I4 => M_reg_9_18,
   O => W_24_19_i_16_n_0
);
W_24_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x116_out_14,
   I1 => M_reg_9_17,
   I2 => M_reg_9_21,
   I3 => M_reg_9_0,
   I4 => M_reg_8_14,
   O => W_24_19_i_17_n_0
);
W_24_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x111_out_28,
   I1 => x111_out_3,
   I2 => x111_out_5,
   I3 => W_24_19_i_10_n_0,
   I4 => W_24_19_i_11_n_0,
   O => W_24_19_i_2_n_0
);
W_24_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x111_out_27,
   I1 => x111_out_2,
   I2 => x111_out_4,
   I3 => W_24_19_i_12_n_0,
   I4 => W_24_19_i_13_n_0,
   O => W_24_19_i_3_n_0
);
W_24_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x111_out_26,
   I1 => x111_out_1,
   I2 => x111_out_3,
   I3 => W_24_19_i_14_n_0,
   I4 => W_24_19_i_15_n_0,
   O => W_24_19_i_4_n_0
);
W_24_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x111_out_25,
   I1 => x111_out_0,
   I2 => x111_out_2,
   I3 => W_24_19_i_16_n_0,
   I4 => W_24_19_i_17_n_0,
   O => W_24_19_i_5_n_0
);
W_24_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_24_19_i_2_n_0,
   I1 => W_24_23_i_16_n_0,
   I2 => x111_out_29,
   I3 => x111_out_4,
   I4 => x111_out_6,
   I5 => W_24_23_i_17_n_0,
   O => W_24_19_i_6_n_0
);
W_24_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_24_19_i_3_n_0,
   I1 => W_24_19_i_10_n_0,
   I2 => x111_out_28,
   I3 => x111_out_3,
   I4 => x111_out_5,
   I5 => W_24_19_i_11_n_0,
   O => W_24_19_i_7_n_0
);
W_24_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_24_19_i_4_n_0,
   I1 => W_24_19_i_12_n_0,
   I2 => x111_out_27,
   I3 => x111_out_2,
   I4 => x111_out_4,
   I5 => W_24_19_i_13_n_0,
   O => W_24_19_i_8_n_0
);
W_24_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_24_19_i_5_n_0,
   I1 => W_24_19_i_14_n_0,
   I2 => x111_out_26,
   I3 => x111_out_1,
   I4 => x111_out_3,
   I5 => W_24_19_i_15_n_0,
   O => W_24_19_i_9_n_0
);
W_24_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_8_22,
   I1 => x116_out_22,
   I2 => M_reg_9_8,
   I3 => M_reg_9_29,
   I4 => M_reg_9_25,
   O => W_24_23_i_10_n_0
);
W_24_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x116_out_21,
   I1 => M_reg_9_24,
   I2 => M_reg_9_28,
   I3 => M_reg_9_7,
   I4 => M_reg_8_21,
   O => W_24_23_i_11_n_0
);
W_24_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_8_21,
   I1 => x116_out_21,
   I2 => M_reg_9_7,
   I3 => M_reg_9_28,
   I4 => M_reg_9_24,
   O => W_24_23_i_12_n_0
);
W_24_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x116_out_20,
   I1 => M_reg_9_23,
   I2 => M_reg_9_27,
   I3 => M_reg_9_6,
   I4 => M_reg_8_20,
   O => W_24_23_i_13_n_0
);
W_24_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_8_20,
   I1 => x116_out_20,
   I2 => M_reg_9_6,
   I3 => M_reg_9_27,
   I4 => M_reg_9_23,
   O => W_24_23_i_14_n_0
);
W_24_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x116_out_19,
   I1 => M_reg_9_22,
   I2 => M_reg_9_26,
   I3 => M_reg_9_5,
   I4 => M_reg_8_19,
   O => W_24_23_i_15_n_0
);
W_24_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_8_19,
   I1 => x116_out_19,
   I2 => M_reg_9_5,
   I3 => M_reg_9_26,
   I4 => M_reg_9_22,
   O => W_24_23_i_16_n_0
);
W_24_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x116_out_18,
   I1 => M_reg_9_21,
   I2 => M_reg_9_25,
   I3 => M_reg_9_4,
   I4 => M_reg_8_18,
   O => W_24_23_i_17_n_0
);
W_24_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x111_out_7,
   I1 => x111_out_9,
   I2 => W_24_23_i_10_n_0,
   I3 => W_24_23_i_11_n_0,
   O => W_24_23_i_2_n_0
);
W_24_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x111_out_31,
   I1 => x111_out_6,
   I2 => x111_out_8,
   I3 => W_24_23_i_12_n_0,
   I4 => W_24_23_i_13_n_0,
   O => W_24_23_i_3_n_0
);
W_24_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x111_out_30,
   I1 => x111_out_5,
   I2 => x111_out_7,
   I3 => W_24_23_i_14_n_0,
   I4 => W_24_23_i_15_n_0,
   O => W_24_23_i_4_n_0
);
W_24_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x111_out_29,
   I1 => x111_out_4,
   I2 => x111_out_6,
   I3 => W_24_23_i_16_n_0,
   I4 => W_24_23_i_17_n_0,
   O => W_24_23_i_5_n_0
);
W_24_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x111_out_8,
   I1 => x111_out_10,
   I2 => W_24_27_i_16_n_0,
   I3 => W_24_27_i_17_n_0,
   I4 => W_24_23_i_2_n_0,
   O => W_24_23_i_6_n_0
);
W_24_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x111_out_7,
   I1 => x111_out_9,
   I2 => W_24_23_i_10_n_0,
   I3 => W_24_23_i_11_n_0,
   I4 => W_24_23_i_3_n_0,
   O => W_24_23_i_7_n_0
);
W_24_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_24_23_i_4_n_0,
   I1 => W_24_23_i_12_n_0,
   I2 => x111_out_31,
   I3 => x111_out_6,
   I4 => x111_out_8,
   I5 => W_24_23_i_13_n_0,
   O => W_24_23_i_8_n_0
);
W_24_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_24_23_i_5_n_0,
   I1 => W_24_23_i_14_n_0,
   I2 => x111_out_30,
   I3 => x111_out_5,
   I4 => x111_out_7,
   I5 => W_24_23_i_15_n_0,
   O => W_24_23_i_9_n_0
);
W_24_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_8_26,
   I1 => x116_out_26,
   I2 => M_reg_9_12,
   I3 => M_reg_9_1,
   I4 => M_reg_9_29,
   O => W_24_27_i_10_n_0
);
W_24_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x116_out_25,
   I1 => M_reg_9_28,
   I2 => M_reg_9_0,
   I3 => M_reg_9_11,
   I4 => M_reg_8_25,
   O => W_24_27_i_11_n_0
);
W_24_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_8_25,
   I1 => x116_out_25,
   I2 => M_reg_9_11,
   I3 => M_reg_9_0,
   I4 => M_reg_9_28,
   O => W_24_27_i_12_n_0
);
W_24_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x116_out_24,
   I1 => M_reg_9_27,
   I2 => M_reg_9_31,
   I3 => M_reg_9_10,
   I4 => M_reg_8_24,
   O => W_24_27_i_13_n_0
);
W_24_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_8_24,
   I1 => x116_out_24,
   I2 => M_reg_9_10,
   I3 => M_reg_9_31,
   I4 => M_reg_9_27,
   O => W_24_27_i_14_n_0
);
W_24_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x116_out_23,
   I1 => M_reg_9_26,
   I2 => M_reg_9_30,
   I3 => M_reg_9_9,
   I4 => M_reg_8_23,
   O => W_24_27_i_15_n_0
);
W_24_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_8_23,
   I1 => x116_out_23,
   I2 => M_reg_9_9,
   I3 => M_reg_9_30,
   I4 => M_reg_9_26,
   O => W_24_27_i_16_n_0
);
W_24_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x116_out_22,
   I1 => M_reg_9_25,
   I2 => M_reg_9_29,
   I3 => M_reg_9_8,
   I4 => M_reg_8_22,
   O => W_24_27_i_17_n_0
);
W_24_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x111_out_11,
   I1 => x111_out_13,
   I2 => W_24_27_i_10_n_0,
   I3 => W_24_27_i_11_n_0,
   O => W_24_27_i_2_n_0
);
W_24_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x111_out_10,
   I1 => x111_out_12,
   I2 => W_24_27_i_12_n_0,
   I3 => W_24_27_i_13_n_0,
   O => W_24_27_i_3_n_0
);
W_24_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x111_out_9,
   I1 => x111_out_11,
   I2 => W_24_27_i_14_n_0,
   I3 => W_24_27_i_15_n_0,
   O => W_24_27_i_4_n_0
);
W_24_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x111_out_8,
   I1 => x111_out_10,
   I2 => W_24_27_i_16_n_0,
   I3 => W_24_27_i_17_n_0,
   O => W_24_27_i_5_n_0
);
W_24_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x111_out_12,
   I1 => x111_out_14,
   I2 => W_24_31_i_13_n_0,
   I3 => W_24_31_i_14_n_0,
   I4 => W_24_27_i_2_n_0,
   O => W_24_27_i_6_n_0
);
W_24_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x111_out_11,
   I1 => x111_out_13,
   I2 => W_24_27_i_10_n_0,
   I3 => W_24_27_i_11_n_0,
   I4 => W_24_27_i_3_n_0,
   O => W_24_27_i_7_n_0
);
W_24_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x111_out_10,
   I1 => x111_out_12,
   I2 => W_24_27_i_12_n_0,
   I3 => W_24_27_i_13_n_0,
   I4 => W_24_27_i_4_n_0,
   O => W_24_27_i_8_n_0
);
W_24_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x111_out_9,
   I1 => x111_out_11,
   I2 => W_24_27_i_14_n_0,
   I3 => W_24_27_i_15_n_0,
   I4 => W_24_27_i_5_n_0,
   O => W_24_27_i_9_n_0
);
W_24_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x116_out_28,
   I1 => M_reg_9_31,
   I2 => M_reg_9_3,
   I3 => M_reg_9_14,
   I4 => M_reg_8_28,
   O => W_24_31_i_10_n_0
);
W_24_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_8_28,
   I1 => x116_out_28,
   I2 => M_reg_9_14,
   I3 => M_reg_9_3,
   I4 => M_reg_9_31,
   O => W_24_31_i_11_n_0
);
W_24_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x116_out_27,
   I1 => M_reg_9_30,
   I2 => M_reg_9_2,
   I3 => M_reg_9_13,
   I4 => M_reg_8_27,
   O => W_24_31_i_12_n_0
);
W_24_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_8_27,
   I1 => x116_out_27,
   I2 => M_reg_9_13,
   I3 => M_reg_9_2,
   I4 => M_reg_9_30,
   O => W_24_31_i_13_n_0
);
W_24_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x116_out_26,
   I1 => M_reg_9_29,
   I2 => M_reg_9_1,
   I3 => M_reg_9_12,
   I4 => M_reg_8_26,
   O => W_24_31_i_14_n_0
);
W_24_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x116_out_29,
   I1 => M_reg_9_4,
   I2 => M_reg_9_15,
   I3 => M_reg_8_29,
   O => W_24_31_i_15_n_0
);
W_24_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x111_out_17,
   I1 => x111_out_15,
   O => SIGMA_LCASE_1323_out_0_30
);
W_24_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => M_reg_9_6,
   I1 => M_reg_9_17,
   I2 => x116_out_31,
   I3 => M_reg_8_31,
   I4 => x111_out_16,
   I5 => x111_out_18,
   O => W_24_31_i_17_n_0
);
W_24_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => M_reg_9_16,
   I1 => M_reg_9_5,
   O => SIGMA_LCASE_0319_out_30
);
W_24_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => M_reg_8_30,
   I1 => x116_out_30,
   I2 => M_reg_9_16,
   I3 => M_reg_9_5,
   O => W_24_31_i_19_n_0
);
W_24_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x111_out_14,
   I1 => x111_out_16,
   I2 => W_24_31_i_9_n_0,
   I3 => W_24_31_i_10_n_0,
   O => W_24_31_i_2_n_0
);
W_24_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x111_out_13,
   I1 => x111_out_15,
   I2 => W_24_31_i_11_n_0,
   I3 => W_24_31_i_12_n_0,
   O => W_24_31_i_3_n_0
);
W_24_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x111_out_12,
   I1 => x111_out_14,
   I2 => W_24_31_i_13_n_0,
   I3 => W_24_31_i_14_n_0,
   O => W_24_31_i_4_n_0
);
W_24_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_24_31_i_15_n_0,
   I1 => SIGMA_LCASE_1323_out_0_30,
   I2 => W_24_31_i_17_n_0,
   I3 => x116_out_30,
   I4 => SIGMA_LCASE_0319_out_30,
   I5 => M_reg_8_30,
   O => W_24_31_i_5_n_0
);
W_24_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_24_31_i_2_n_0,
   I1 => W_24_31_i_19_n_0,
   I2 => x111_out_15,
   I3 => x111_out_17,
   I4 => W_24_31_i_15_n_0,
   O => W_24_31_i_6_n_0
);
W_24_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x111_out_14,
   I1 => x111_out_16,
   I2 => W_24_31_i_9_n_0,
   I3 => W_24_31_i_10_n_0,
   I4 => W_24_31_i_3_n_0,
   O => W_24_31_i_7_n_0
);
W_24_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x111_out_13,
   I1 => x111_out_15,
   I2 => W_24_31_i_11_n_0,
   I3 => W_24_31_i_12_n_0,
   I4 => W_24_31_i_4_n_0,
   O => W_24_31_i_8_n_0
);
W_24_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => M_reg_8_29,
   I1 => x116_out_29,
   I2 => M_reg_9_15,
   I3 => M_reg_9_4,
   O => W_24_31_i_9_n_0
);
W_24_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_8_2,
   I1 => x116_out_2,
   I2 => M_reg_9_20,
   I3 => M_reg_9_9,
   I4 => M_reg_9_5,
   O => W_24_3_i_10_n_0
);
W_24_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x116_out_1,
   I1 => M_reg_9_4,
   I2 => M_reg_9_8,
   I3 => M_reg_9_19,
   I4 => M_reg_8_1,
   O => W_24_3_i_11_n_0
);
W_24_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => M_reg_9_19,
   I1 => M_reg_9_8,
   I2 => M_reg_9_4,
   O => SIGMA_LCASE_0319_out_1
);
W_24_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x111_out_21,
   I1 => x111_out_19,
   I2 => x111_out_12,
   O => SIGMA_LCASE_1323_out_0_2
);
W_24_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x111_out_20,
   I1 => x111_out_18,
   I2 => x111_out_11,
   O => SIGMA_LCASE_1323_out_1
);
W_24_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x111_out_12,
   I1 => x111_out_19,
   I2 => x111_out_21,
   I3 => W_24_3_i_10_n_0,
   I4 => W_24_3_i_11_n_0,
   O => W_24_3_i_2_n_0
);
W_24_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_24_3_i_11_n_0,
   I1 => x111_out_21,
   I2 => x111_out_19,
   I3 => x111_out_12,
   I4 => W_24_3_i_10_n_0,
   O => W_24_3_i_3_n_0
);
W_24_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_0319_out_1,
   I1 => x116_out_1,
   I2 => M_reg_8_1,
   I3 => x111_out_11,
   I4 => x111_out_18,
   I5 => x111_out_20,
   O => W_24_3_i_4_n_0
);
W_24_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_8_0,
   I1 => x116_out_0,
   I2 => M_reg_9_18,
   I3 => M_reg_9_7,
   I4 => M_reg_9_3,
   O => W_24_3_i_5_n_0
);
W_24_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_24_3_i_2_n_0,
   I1 => W_24_7_i_16_n_0,
   I2 => x111_out_13,
   I3 => x111_out_20,
   I4 => x111_out_22,
   I5 => W_24_7_i_17_n_0,
   O => W_24_3_i_6_n_0
);
W_24_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_24_3_i_10_n_0,
   I1 => SIGMA_LCASE_1323_out_0_2,
   I2 => M_reg_8_1,
   I3 => x116_out_1,
   I4 => SIGMA_LCASE_0319_out_1,
   I5 => SIGMA_LCASE_1323_out_1,
   O => W_24_3_i_7_n_0
);
W_24_3_i_8 : LUT6
  generic map(
   INIT => X"566565566aa6a66a"
  )
 port map (
   I0 => W_24_3_i_4_n_0,
   I1 => M_reg_8_0,
   I2 => M_reg_9_18,
   I3 => M_reg_9_7,
   I4 => M_reg_9_3,
   I5 => x116_out_0,
   O => W_24_3_i_8_n_0
);
W_24_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_24_3_i_5_n_0,
   I1 => x111_out_10,
   I2 => x111_out_17,
   I3 => x111_out_19,
   O => W_24_3_i_9_n_0
);
W_24_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_8_6,
   I1 => x116_out_6,
   I2 => M_reg_9_24,
   I3 => M_reg_9_13,
   I4 => M_reg_9_9,
   O => W_24_7_i_10_n_0
);
W_24_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x116_out_5,
   I1 => M_reg_9_8,
   I2 => M_reg_9_12,
   I3 => M_reg_9_23,
   I4 => M_reg_8_5,
   O => W_24_7_i_11_n_0
);
W_24_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_8_5,
   I1 => x116_out_5,
   I2 => M_reg_9_23,
   I3 => M_reg_9_12,
   I4 => M_reg_9_8,
   O => W_24_7_i_12_n_0
);
W_24_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x116_out_4,
   I1 => M_reg_9_7,
   I2 => M_reg_9_11,
   I3 => M_reg_9_22,
   I4 => M_reg_8_4,
   O => W_24_7_i_13_n_0
);
W_24_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_8_4,
   I1 => x116_out_4,
   I2 => M_reg_9_22,
   I3 => M_reg_9_11,
   I4 => M_reg_9_7,
   O => W_24_7_i_14_n_0
);
W_24_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x116_out_3,
   I1 => M_reg_9_6,
   I2 => M_reg_9_10,
   I3 => M_reg_9_21,
   I4 => M_reg_8_3,
   O => W_24_7_i_15_n_0
);
W_24_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_8_3,
   I1 => x116_out_3,
   I2 => M_reg_9_21,
   I3 => M_reg_9_10,
   I4 => M_reg_9_6,
   O => W_24_7_i_16_n_0
);
W_24_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x116_out_2,
   I1 => M_reg_9_5,
   I2 => M_reg_9_9,
   I3 => M_reg_9_20,
   I4 => M_reg_8_2,
   O => W_24_7_i_17_n_0
);
W_24_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x111_out_16,
   I1 => x111_out_23,
   I2 => x111_out_25,
   I3 => W_24_7_i_10_n_0,
   I4 => W_24_7_i_11_n_0,
   O => W_24_7_i_2_n_0
);
W_24_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x111_out_15,
   I1 => x111_out_22,
   I2 => x111_out_24,
   I3 => W_24_7_i_12_n_0,
   I4 => W_24_7_i_13_n_0,
   O => W_24_7_i_3_n_0
);
W_24_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x111_out_14,
   I1 => x111_out_21,
   I2 => x111_out_23,
   I3 => W_24_7_i_14_n_0,
   I4 => W_24_7_i_15_n_0,
   O => W_24_7_i_4_n_0
);
W_24_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x111_out_13,
   I1 => x111_out_20,
   I2 => x111_out_22,
   I3 => W_24_7_i_16_n_0,
   I4 => W_24_7_i_17_n_0,
   O => W_24_7_i_5_n_0
);
W_24_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_24_7_i_2_n_0,
   I1 => W_24_11_i_16_n_0,
   I2 => x111_out_17,
   I3 => x111_out_24,
   I4 => x111_out_26,
   I5 => W_24_11_i_17_n_0,
   O => W_24_7_i_6_n_0
);
W_24_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_24_7_i_3_n_0,
   I1 => W_24_7_i_10_n_0,
   I2 => x111_out_16,
   I3 => x111_out_23,
   I4 => x111_out_25,
   I5 => W_24_7_i_11_n_0,
   O => W_24_7_i_7_n_0
);
W_24_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_24_7_i_4_n_0,
   I1 => W_24_7_i_12_n_0,
   I2 => x111_out_15,
   I3 => x111_out_22,
   I4 => x111_out_24,
   I5 => W_24_7_i_13_n_0,
   O => W_24_7_i_8_n_0
);
W_24_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_24_7_i_5_n_0,
   I1 => W_24_7_i_14_n_0,
   I2 => x111_out_14,
   I3 => x111_out_21,
   I4 => x111_out_23,
   I5 => W_24_7_i_15_n_0,
   O => W_24_7_i_9_n_0
);
W_25_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_9_10,
   I1 => x115_out_10,
   I2 => M_reg_10_28,
   I3 => M_reg_10_17,
   I4 => M_reg_10_13,
   O => W_25_11_i_10_n_0
);
W_25_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x115_out_9,
   I1 => M_reg_10_12,
   I2 => M_reg_10_16,
   I3 => M_reg_10_27,
   I4 => M_reg_9_9,
   O => W_25_11_i_11_n_0
);
W_25_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_9_9,
   I1 => x115_out_9,
   I2 => M_reg_10_27,
   I3 => M_reg_10_16,
   I4 => M_reg_10_12,
   O => W_25_11_i_12_n_0
);
W_25_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x115_out_8,
   I1 => M_reg_10_11,
   I2 => M_reg_10_15,
   I3 => M_reg_10_26,
   I4 => M_reg_9_8,
   O => W_25_11_i_13_n_0
);
W_25_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_9_8,
   I1 => x115_out_8,
   I2 => M_reg_10_26,
   I3 => M_reg_10_15,
   I4 => M_reg_10_11,
   O => W_25_11_i_14_n_0
);
W_25_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x115_out_7,
   I1 => M_reg_10_10,
   I2 => M_reg_10_14,
   I3 => M_reg_10_25,
   I4 => M_reg_9_7,
   O => W_25_11_i_15_n_0
);
W_25_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_9_7,
   I1 => x115_out_7,
   I2 => M_reg_10_25,
   I3 => M_reg_10_14,
   I4 => M_reg_10_10,
   O => W_25_11_i_16_n_0
);
W_25_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x115_out_6,
   I1 => M_reg_10_9,
   I2 => M_reg_10_13,
   I3 => M_reg_10_24,
   I4 => M_reg_9_6,
   O => W_25_11_i_17_n_0
);
W_25_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x110_out_20,
   I1 => x110_out_27,
   I2 => x110_out_29,
   I3 => W_25_11_i_10_n_0,
   I4 => W_25_11_i_11_n_0,
   O => W_25_11_i_2_n_0
);
W_25_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x110_out_19,
   I1 => x110_out_26,
   I2 => x110_out_28,
   I3 => W_25_11_i_12_n_0,
   I4 => W_25_11_i_13_n_0,
   O => W_25_11_i_3_n_0
);
W_25_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x110_out_18,
   I1 => x110_out_25,
   I2 => x110_out_27,
   I3 => W_25_11_i_14_n_0,
   I4 => W_25_11_i_15_n_0,
   O => W_25_11_i_4_n_0
);
W_25_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x110_out_17,
   I1 => x110_out_24,
   I2 => x110_out_26,
   I3 => W_25_11_i_16_n_0,
   I4 => W_25_11_i_17_n_0,
   O => W_25_11_i_5_n_0
);
W_25_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_25_11_i_2_n_0,
   I1 => W_25_15_i_16_n_0,
   I2 => x110_out_21,
   I3 => x110_out_28,
   I4 => x110_out_30,
   I5 => W_25_15_i_17_n_0,
   O => W_25_11_i_6_n_0
);
W_25_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_25_11_i_3_n_0,
   I1 => W_25_11_i_10_n_0,
   I2 => x110_out_20,
   I3 => x110_out_27,
   I4 => x110_out_29,
   I5 => W_25_11_i_11_n_0,
   O => W_25_11_i_7_n_0
);
W_25_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_25_11_i_4_n_0,
   I1 => W_25_11_i_12_n_0,
   I2 => x110_out_19,
   I3 => x110_out_26,
   I4 => x110_out_28,
   I5 => W_25_11_i_13_n_0,
   O => W_25_11_i_8_n_0
);
W_25_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_25_11_i_5_n_0,
   I1 => W_25_11_i_14_n_0,
   I2 => x110_out_18,
   I3 => x110_out_25,
   I4 => x110_out_27,
   I5 => W_25_11_i_15_n_0,
   O => W_25_11_i_9_n_0
);
W_25_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_9_14,
   I1 => x115_out_14,
   I2 => M_reg_10_0,
   I3 => M_reg_10_21,
   I4 => M_reg_10_17,
   O => W_25_15_i_10_n_0
);
W_25_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x115_out_13,
   I1 => M_reg_10_16,
   I2 => M_reg_10_20,
   I3 => M_reg_10_31,
   I4 => M_reg_9_13,
   O => W_25_15_i_11_n_0
);
W_25_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_9_13,
   I1 => x115_out_13,
   I2 => M_reg_10_31,
   I3 => M_reg_10_20,
   I4 => M_reg_10_16,
   O => W_25_15_i_12_n_0
);
W_25_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x115_out_12,
   I1 => M_reg_10_15,
   I2 => M_reg_10_19,
   I3 => M_reg_10_30,
   I4 => M_reg_9_12,
   O => W_25_15_i_13_n_0
);
W_25_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_9_12,
   I1 => x115_out_12,
   I2 => M_reg_10_30,
   I3 => M_reg_10_19,
   I4 => M_reg_10_15,
   O => W_25_15_i_14_n_0
);
W_25_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x115_out_11,
   I1 => M_reg_10_14,
   I2 => M_reg_10_18,
   I3 => M_reg_10_29,
   I4 => M_reg_9_11,
   O => W_25_15_i_15_n_0
);
W_25_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_9_11,
   I1 => x115_out_11,
   I2 => M_reg_10_29,
   I3 => M_reg_10_18,
   I4 => M_reg_10_14,
   O => W_25_15_i_16_n_0
);
W_25_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x115_out_10,
   I1 => M_reg_10_13,
   I2 => M_reg_10_17,
   I3 => M_reg_10_28,
   I4 => M_reg_9_10,
   O => W_25_15_i_17_n_0
);
W_25_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x110_out_24,
   I1 => x110_out_31,
   I2 => x110_out_1,
   I3 => W_25_15_i_10_n_0,
   I4 => W_25_15_i_11_n_0,
   O => W_25_15_i_2_n_0
);
W_25_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x110_out_23,
   I1 => x110_out_30,
   I2 => x110_out_0,
   I3 => W_25_15_i_12_n_0,
   I4 => W_25_15_i_13_n_0,
   O => W_25_15_i_3_n_0
);
W_25_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x110_out_22,
   I1 => x110_out_29,
   I2 => x110_out_31,
   I3 => W_25_15_i_14_n_0,
   I4 => W_25_15_i_15_n_0,
   O => W_25_15_i_4_n_0
);
W_25_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x110_out_21,
   I1 => x110_out_28,
   I2 => x110_out_30,
   I3 => W_25_15_i_16_n_0,
   I4 => W_25_15_i_17_n_0,
   O => W_25_15_i_5_n_0
);
W_25_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_25_15_i_2_n_0,
   I1 => W_25_19_i_16_n_0,
   I2 => x110_out_25,
   I3 => x110_out_0,
   I4 => x110_out_2,
   I5 => W_25_19_i_17_n_0,
   O => W_25_15_i_6_n_0
);
W_25_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_25_15_i_3_n_0,
   I1 => W_25_15_i_10_n_0,
   I2 => x110_out_24,
   I3 => x110_out_31,
   I4 => x110_out_1,
   I5 => W_25_15_i_11_n_0,
   O => W_25_15_i_7_n_0
);
W_25_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_25_15_i_4_n_0,
   I1 => W_25_15_i_12_n_0,
   I2 => x110_out_23,
   I3 => x110_out_30,
   I4 => x110_out_0,
   I5 => W_25_15_i_13_n_0,
   O => W_25_15_i_8_n_0
);
W_25_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_25_15_i_5_n_0,
   I1 => W_25_15_i_14_n_0,
   I2 => x110_out_22,
   I3 => x110_out_29,
   I4 => x110_out_31,
   I5 => W_25_15_i_15_n_0,
   O => W_25_15_i_9_n_0
);
W_25_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_9_18,
   I1 => x115_out_18,
   I2 => M_reg_10_4,
   I3 => M_reg_10_25,
   I4 => M_reg_10_21,
   O => W_25_19_i_10_n_0
);
W_25_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x115_out_17,
   I1 => M_reg_10_20,
   I2 => M_reg_10_24,
   I3 => M_reg_10_3,
   I4 => M_reg_9_17,
   O => W_25_19_i_11_n_0
);
W_25_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_9_17,
   I1 => x115_out_17,
   I2 => M_reg_10_3,
   I3 => M_reg_10_24,
   I4 => M_reg_10_20,
   O => W_25_19_i_12_n_0
);
W_25_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x115_out_16,
   I1 => M_reg_10_19,
   I2 => M_reg_10_23,
   I3 => M_reg_10_2,
   I4 => M_reg_9_16,
   O => W_25_19_i_13_n_0
);
W_25_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_9_16,
   I1 => x115_out_16,
   I2 => M_reg_10_2,
   I3 => M_reg_10_23,
   I4 => M_reg_10_19,
   O => W_25_19_i_14_n_0
);
W_25_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x115_out_15,
   I1 => M_reg_10_18,
   I2 => M_reg_10_22,
   I3 => M_reg_10_1,
   I4 => M_reg_9_15,
   O => W_25_19_i_15_n_0
);
W_25_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_9_15,
   I1 => x115_out_15,
   I2 => M_reg_10_1,
   I3 => M_reg_10_22,
   I4 => M_reg_10_18,
   O => W_25_19_i_16_n_0
);
W_25_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x115_out_14,
   I1 => M_reg_10_17,
   I2 => M_reg_10_21,
   I3 => M_reg_10_0,
   I4 => M_reg_9_14,
   O => W_25_19_i_17_n_0
);
W_25_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x110_out_28,
   I1 => x110_out_3,
   I2 => x110_out_5,
   I3 => W_25_19_i_10_n_0,
   I4 => W_25_19_i_11_n_0,
   O => W_25_19_i_2_n_0
);
W_25_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x110_out_27,
   I1 => x110_out_2,
   I2 => x110_out_4,
   I3 => W_25_19_i_12_n_0,
   I4 => W_25_19_i_13_n_0,
   O => W_25_19_i_3_n_0
);
W_25_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x110_out_26,
   I1 => x110_out_1,
   I2 => x110_out_3,
   I3 => W_25_19_i_14_n_0,
   I4 => W_25_19_i_15_n_0,
   O => W_25_19_i_4_n_0
);
W_25_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x110_out_25,
   I1 => x110_out_0,
   I2 => x110_out_2,
   I3 => W_25_19_i_16_n_0,
   I4 => W_25_19_i_17_n_0,
   O => W_25_19_i_5_n_0
);
W_25_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_25_19_i_2_n_0,
   I1 => W_25_23_i_16_n_0,
   I2 => x110_out_29,
   I3 => x110_out_4,
   I4 => x110_out_6,
   I5 => W_25_23_i_17_n_0,
   O => W_25_19_i_6_n_0
);
W_25_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_25_19_i_3_n_0,
   I1 => W_25_19_i_10_n_0,
   I2 => x110_out_28,
   I3 => x110_out_3,
   I4 => x110_out_5,
   I5 => W_25_19_i_11_n_0,
   O => W_25_19_i_7_n_0
);
W_25_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_25_19_i_4_n_0,
   I1 => W_25_19_i_12_n_0,
   I2 => x110_out_27,
   I3 => x110_out_2,
   I4 => x110_out_4,
   I5 => W_25_19_i_13_n_0,
   O => W_25_19_i_8_n_0
);
W_25_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_25_19_i_5_n_0,
   I1 => W_25_19_i_14_n_0,
   I2 => x110_out_26,
   I3 => x110_out_1,
   I4 => x110_out_3,
   I5 => W_25_19_i_15_n_0,
   O => W_25_19_i_9_n_0
);
W_25_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_9_22,
   I1 => x115_out_22,
   I2 => M_reg_10_8,
   I3 => M_reg_10_29,
   I4 => M_reg_10_25,
   O => W_25_23_i_10_n_0
);
W_25_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x115_out_21,
   I1 => M_reg_10_24,
   I2 => M_reg_10_28,
   I3 => M_reg_10_7,
   I4 => M_reg_9_21,
   O => W_25_23_i_11_n_0
);
W_25_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_9_21,
   I1 => x115_out_21,
   I2 => M_reg_10_7,
   I3 => M_reg_10_28,
   I4 => M_reg_10_24,
   O => W_25_23_i_12_n_0
);
W_25_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x115_out_20,
   I1 => M_reg_10_23,
   I2 => M_reg_10_27,
   I3 => M_reg_10_6,
   I4 => M_reg_9_20,
   O => W_25_23_i_13_n_0
);
W_25_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_9_20,
   I1 => x115_out_20,
   I2 => M_reg_10_6,
   I3 => M_reg_10_27,
   I4 => M_reg_10_23,
   O => W_25_23_i_14_n_0
);
W_25_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x115_out_19,
   I1 => M_reg_10_22,
   I2 => M_reg_10_26,
   I3 => M_reg_10_5,
   I4 => M_reg_9_19,
   O => W_25_23_i_15_n_0
);
W_25_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_9_19,
   I1 => x115_out_19,
   I2 => M_reg_10_5,
   I3 => M_reg_10_26,
   I4 => M_reg_10_22,
   O => W_25_23_i_16_n_0
);
W_25_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x115_out_18,
   I1 => M_reg_10_21,
   I2 => M_reg_10_25,
   I3 => M_reg_10_4,
   I4 => M_reg_9_18,
   O => W_25_23_i_17_n_0
);
W_25_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x110_out_7,
   I1 => x110_out_9,
   I2 => W_25_23_i_10_n_0,
   I3 => W_25_23_i_11_n_0,
   O => W_25_23_i_2_n_0
);
W_25_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x110_out_31,
   I1 => x110_out_6,
   I2 => x110_out_8,
   I3 => W_25_23_i_12_n_0,
   I4 => W_25_23_i_13_n_0,
   O => W_25_23_i_3_n_0
);
W_25_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x110_out_30,
   I1 => x110_out_5,
   I2 => x110_out_7,
   I3 => W_25_23_i_14_n_0,
   I4 => W_25_23_i_15_n_0,
   O => W_25_23_i_4_n_0
);
W_25_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x110_out_29,
   I1 => x110_out_4,
   I2 => x110_out_6,
   I3 => W_25_23_i_16_n_0,
   I4 => W_25_23_i_17_n_0,
   O => W_25_23_i_5_n_0
);
W_25_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x110_out_8,
   I1 => x110_out_10,
   I2 => W_25_27_i_16_n_0,
   I3 => W_25_27_i_17_n_0,
   I4 => W_25_23_i_2_n_0,
   O => W_25_23_i_6_n_0
);
W_25_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x110_out_7,
   I1 => x110_out_9,
   I2 => W_25_23_i_10_n_0,
   I3 => W_25_23_i_11_n_0,
   I4 => W_25_23_i_3_n_0,
   O => W_25_23_i_7_n_0
);
W_25_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_25_23_i_4_n_0,
   I1 => W_25_23_i_12_n_0,
   I2 => x110_out_31,
   I3 => x110_out_6,
   I4 => x110_out_8,
   I5 => W_25_23_i_13_n_0,
   O => W_25_23_i_8_n_0
);
W_25_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_25_23_i_5_n_0,
   I1 => W_25_23_i_14_n_0,
   I2 => x110_out_30,
   I3 => x110_out_5,
   I4 => x110_out_7,
   I5 => W_25_23_i_15_n_0,
   O => W_25_23_i_9_n_0
);
W_25_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_9_26,
   I1 => x115_out_26,
   I2 => M_reg_10_12,
   I3 => M_reg_10_1,
   I4 => M_reg_10_29,
   O => W_25_27_i_10_n_0
);
W_25_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x115_out_25,
   I1 => M_reg_10_28,
   I2 => M_reg_10_0,
   I3 => M_reg_10_11,
   I4 => M_reg_9_25,
   O => W_25_27_i_11_n_0
);
W_25_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_9_25,
   I1 => x115_out_25,
   I2 => M_reg_10_11,
   I3 => M_reg_10_0,
   I4 => M_reg_10_28,
   O => W_25_27_i_12_n_0
);
W_25_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x115_out_24,
   I1 => M_reg_10_27,
   I2 => M_reg_10_31,
   I3 => M_reg_10_10,
   I4 => M_reg_9_24,
   O => W_25_27_i_13_n_0
);
W_25_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_9_24,
   I1 => x115_out_24,
   I2 => M_reg_10_10,
   I3 => M_reg_10_31,
   I4 => M_reg_10_27,
   O => W_25_27_i_14_n_0
);
W_25_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x115_out_23,
   I1 => M_reg_10_26,
   I2 => M_reg_10_30,
   I3 => M_reg_10_9,
   I4 => M_reg_9_23,
   O => W_25_27_i_15_n_0
);
W_25_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_9_23,
   I1 => x115_out_23,
   I2 => M_reg_10_9,
   I3 => M_reg_10_30,
   I4 => M_reg_10_26,
   O => W_25_27_i_16_n_0
);
W_25_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x115_out_22,
   I1 => M_reg_10_25,
   I2 => M_reg_10_29,
   I3 => M_reg_10_8,
   I4 => M_reg_9_22,
   O => W_25_27_i_17_n_0
);
W_25_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x110_out_11,
   I1 => x110_out_13,
   I2 => W_25_27_i_10_n_0,
   I3 => W_25_27_i_11_n_0,
   O => W_25_27_i_2_n_0
);
W_25_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x110_out_10,
   I1 => x110_out_12,
   I2 => W_25_27_i_12_n_0,
   I3 => W_25_27_i_13_n_0,
   O => W_25_27_i_3_n_0
);
W_25_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x110_out_9,
   I1 => x110_out_11,
   I2 => W_25_27_i_14_n_0,
   I3 => W_25_27_i_15_n_0,
   O => W_25_27_i_4_n_0
);
W_25_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x110_out_8,
   I1 => x110_out_10,
   I2 => W_25_27_i_16_n_0,
   I3 => W_25_27_i_17_n_0,
   O => W_25_27_i_5_n_0
);
W_25_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x110_out_12,
   I1 => x110_out_14,
   I2 => W_25_31_i_13_n_0,
   I3 => W_25_31_i_14_n_0,
   I4 => W_25_27_i_2_n_0,
   O => W_25_27_i_6_n_0
);
W_25_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x110_out_11,
   I1 => x110_out_13,
   I2 => W_25_27_i_10_n_0,
   I3 => W_25_27_i_11_n_0,
   I4 => W_25_27_i_3_n_0,
   O => W_25_27_i_7_n_0
);
W_25_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x110_out_10,
   I1 => x110_out_12,
   I2 => W_25_27_i_12_n_0,
   I3 => W_25_27_i_13_n_0,
   I4 => W_25_27_i_4_n_0,
   O => W_25_27_i_8_n_0
);
W_25_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x110_out_9,
   I1 => x110_out_11,
   I2 => W_25_27_i_14_n_0,
   I3 => W_25_27_i_15_n_0,
   I4 => W_25_27_i_5_n_0,
   O => W_25_27_i_9_n_0
);
W_25_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x115_out_28,
   I1 => M_reg_10_31,
   I2 => M_reg_10_3,
   I3 => M_reg_10_14,
   I4 => M_reg_9_28,
   O => W_25_31_i_10_n_0
);
W_25_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_9_28,
   I1 => x115_out_28,
   I2 => M_reg_10_14,
   I3 => M_reg_10_3,
   I4 => M_reg_10_31,
   O => W_25_31_i_11_n_0
);
W_25_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x115_out_27,
   I1 => M_reg_10_30,
   I2 => M_reg_10_2,
   I3 => M_reg_10_13,
   I4 => M_reg_9_27,
   O => W_25_31_i_12_n_0
);
W_25_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_9_27,
   I1 => x115_out_27,
   I2 => M_reg_10_13,
   I3 => M_reg_10_2,
   I4 => M_reg_10_30,
   O => W_25_31_i_13_n_0
);
W_25_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x115_out_26,
   I1 => M_reg_10_29,
   I2 => M_reg_10_1,
   I3 => M_reg_10_12,
   I4 => M_reg_9_26,
   O => W_25_31_i_14_n_0
);
W_25_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x115_out_29,
   I1 => M_reg_10_4,
   I2 => M_reg_10_15,
   I3 => M_reg_9_29,
   O => W_25_31_i_15_n_0
);
W_25_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x110_out_17,
   I1 => x110_out_15,
   O => SIGMA_LCASE_1315_out_0_30
);
W_25_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => M_reg_10_6,
   I1 => M_reg_10_17,
   I2 => x115_out_31,
   I3 => M_reg_9_31,
   I4 => x110_out_16,
   I5 => x110_out_18,
   O => W_25_31_i_17_n_0
);
W_25_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => M_reg_10_16,
   I1 => M_reg_10_5,
   O => SIGMA_LCASE_0311_out_30
);
W_25_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => M_reg_9_30,
   I1 => x115_out_30,
   I2 => M_reg_10_16,
   I3 => M_reg_10_5,
   O => W_25_31_i_19_n_0
);
W_25_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x110_out_14,
   I1 => x110_out_16,
   I2 => W_25_31_i_9_n_0,
   I3 => W_25_31_i_10_n_0,
   O => W_25_31_i_2_n_0
);
W_25_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x110_out_13,
   I1 => x110_out_15,
   I2 => W_25_31_i_11_n_0,
   I3 => W_25_31_i_12_n_0,
   O => W_25_31_i_3_n_0
);
W_25_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x110_out_12,
   I1 => x110_out_14,
   I2 => W_25_31_i_13_n_0,
   I3 => W_25_31_i_14_n_0,
   O => W_25_31_i_4_n_0
);
W_25_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_25_31_i_15_n_0,
   I1 => SIGMA_LCASE_1315_out_0_30,
   I2 => W_25_31_i_17_n_0,
   I3 => x115_out_30,
   I4 => SIGMA_LCASE_0311_out_30,
   I5 => M_reg_9_30,
   O => W_25_31_i_5_n_0
);
W_25_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_25_31_i_2_n_0,
   I1 => W_25_31_i_19_n_0,
   I2 => x110_out_15,
   I3 => x110_out_17,
   I4 => W_25_31_i_15_n_0,
   O => W_25_31_i_6_n_0
);
W_25_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x110_out_14,
   I1 => x110_out_16,
   I2 => W_25_31_i_9_n_0,
   I3 => W_25_31_i_10_n_0,
   I4 => W_25_31_i_3_n_0,
   O => W_25_31_i_7_n_0
);
W_25_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x110_out_13,
   I1 => x110_out_15,
   I2 => W_25_31_i_11_n_0,
   I3 => W_25_31_i_12_n_0,
   I4 => W_25_31_i_4_n_0,
   O => W_25_31_i_8_n_0
);
W_25_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => M_reg_9_29,
   I1 => x115_out_29,
   I2 => M_reg_10_15,
   I3 => M_reg_10_4,
   O => W_25_31_i_9_n_0
);
W_25_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_9_2,
   I1 => x115_out_2,
   I2 => M_reg_10_20,
   I3 => M_reg_10_9,
   I4 => M_reg_10_5,
   O => W_25_3_i_10_n_0
);
W_25_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x115_out_1,
   I1 => M_reg_10_4,
   I2 => M_reg_10_8,
   I3 => M_reg_10_19,
   I4 => M_reg_9_1,
   O => W_25_3_i_11_n_0
);
W_25_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => M_reg_10_19,
   I1 => M_reg_10_8,
   I2 => M_reg_10_4,
   O => SIGMA_LCASE_0311_out_1
);
W_25_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x110_out_21,
   I1 => x110_out_19,
   I2 => x110_out_12,
   O => SIGMA_LCASE_1315_out_0_2
);
W_25_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x110_out_20,
   I1 => x110_out_18,
   I2 => x110_out_11,
   O => SIGMA_LCASE_1315_out_1
);
W_25_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x110_out_12,
   I1 => x110_out_19,
   I2 => x110_out_21,
   I3 => W_25_3_i_10_n_0,
   I4 => W_25_3_i_11_n_0,
   O => W_25_3_i_2_n_0
);
W_25_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_25_3_i_11_n_0,
   I1 => x110_out_21,
   I2 => x110_out_19,
   I3 => x110_out_12,
   I4 => W_25_3_i_10_n_0,
   O => W_25_3_i_3_n_0
);
W_25_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_0311_out_1,
   I1 => x115_out_1,
   I2 => M_reg_9_1,
   I3 => x110_out_11,
   I4 => x110_out_18,
   I5 => x110_out_20,
   O => W_25_3_i_4_n_0
);
W_25_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_9_0,
   I1 => x115_out_0,
   I2 => M_reg_10_18,
   I3 => M_reg_10_7,
   I4 => M_reg_10_3,
   O => W_25_3_i_5_n_0
);
W_25_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_25_3_i_2_n_0,
   I1 => W_25_7_i_16_n_0,
   I2 => x110_out_13,
   I3 => x110_out_20,
   I4 => x110_out_22,
   I5 => W_25_7_i_17_n_0,
   O => W_25_3_i_6_n_0
);
W_25_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_25_3_i_10_n_0,
   I1 => SIGMA_LCASE_1315_out_0_2,
   I2 => M_reg_9_1,
   I3 => x115_out_1,
   I4 => SIGMA_LCASE_0311_out_1,
   I5 => SIGMA_LCASE_1315_out_1,
   O => W_25_3_i_7_n_0
);
W_25_3_i_8 : LUT6
  generic map(
   INIT => X"566565566aa6a66a"
  )
 port map (
   I0 => W_25_3_i_4_n_0,
   I1 => M_reg_9_0,
   I2 => M_reg_10_18,
   I3 => M_reg_10_7,
   I4 => M_reg_10_3,
   I5 => x115_out_0,
   O => W_25_3_i_8_n_0
);
W_25_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_25_3_i_5_n_0,
   I1 => x110_out_10,
   I2 => x110_out_17,
   I3 => x110_out_19,
   O => W_25_3_i_9_n_0
);
W_25_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_9_6,
   I1 => x115_out_6,
   I2 => M_reg_10_24,
   I3 => M_reg_10_13,
   I4 => M_reg_10_9,
   O => W_25_7_i_10_n_0
);
W_25_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x115_out_5,
   I1 => M_reg_10_8,
   I2 => M_reg_10_12,
   I3 => M_reg_10_23,
   I4 => M_reg_9_5,
   O => W_25_7_i_11_n_0
);
W_25_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_9_5,
   I1 => x115_out_5,
   I2 => M_reg_10_23,
   I3 => M_reg_10_12,
   I4 => M_reg_10_8,
   O => W_25_7_i_12_n_0
);
W_25_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x115_out_4,
   I1 => M_reg_10_7,
   I2 => M_reg_10_11,
   I3 => M_reg_10_22,
   I4 => M_reg_9_4,
   O => W_25_7_i_13_n_0
);
W_25_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_9_4,
   I1 => x115_out_4,
   I2 => M_reg_10_22,
   I3 => M_reg_10_11,
   I4 => M_reg_10_7,
   O => W_25_7_i_14_n_0
);
W_25_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x115_out_3,
   I1 => M_reg_10_6,
   I2 => M_reg_10_10,
   I3 => M_reg_10_21,
   I4 => M_reg_9_3,
   O => W_25_7_i_15_n_0
);
W_25_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_9_3,
   I1 => x115_out_3,
   I2 => M_reg_10_21,
   I3 => M_reg_10_10,
   I4 => M_reg_10_6,
   O => W_25_7_i_16_n_0
);
W_25_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x115_out_2,
   I1 => M_reg_10_5,
   I2 => M_reg_10_9,
   I3 => M_reg_10_20,
   I4 => M_reg_9_2,
   O => W_25_7_i_17_n_0
);
W_25_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x110_out_16,
   I1 => x110_out_23,
   I2 => x110_out_25,
   I3 => W_25_7_i_10_n_0,
   I4 => W_25_7_i_11_n_0,
   O => W_25_7_i_2_n_0
);
W_25_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x110_out_15,
   I1 => x110_out_22,
   I2 => x110_out_24,
   I3 => W_25_7_i_12_n_0,
   I4 => W_25_7_i_13_n_0,
   O => W_25_7_i_3_n_0
);
W_25_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x110_out_14,
   I1 => x110_out_21,
   I2 => x110_out_23,
   I3 => W_25_7_i_14_n_0,
   I4 => W_25_7_i_15_n_0,
   O => W_25_7_i_4_n_0
);
W_25_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x110_out_13,
   I1 => x110_out_20,
   I2 => x110_out_22,
   I3 => W_25_7_i_16_n_0,
   I4 => W_25_7_i_17_n_0,
   O => W_25_7_i_5_n_0
);
W_25_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_25_7_i_2_n_0,
   I1 => W_25_11_i_16_n_0,
   I2 => x110_out_17,
   I3 => x110_out_24,
   I4 => x110_out_26,
   I5 => W_25_11_i_17_n_0,
   O => W_25_7_i_6_n_0
);
W_25_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_25_7_i_3_n_0,
   I1 => W_25_7_i_10_n_0,
   I2 => x110_out_16,
   I3 => x110_out_23,
   I4 => x110_out_25,
   I5 => W_25_7_i_11_n_0,
   O => W_25_7_i_7_n_0
);
W_25_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_25_7_i_4_n_0,
   I1 => W_25_7_i_12_n_0,
   I2 => x110_out_15,
   I3 => x110_out_22,
   I4 => x110_out_24,
   I5 => W_25_7_i_13_n_0,
   O => W_25_7_i_8_n_0
);
W_25_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_25_7_i_5_n_0,
   I1 => W_25_7_i_14_n_0,
   I2 => x110_out_14,
   I3 => x110_out_21,
   I4 => x110_out_23,
   I5 => W_25_7_i_15_n_0,
   O => W_25_7_i_9_n_0
);
W_26_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_10_10,
   I1 => x114_out_10,
   I2 => M_reg_11_28,
   I3 => M_reg_11_17,
   I4 => M_reg_11_13,
   O => W_26_11_i_10_n_0
);
W_26_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x114_out_9,
   I1 => M_reg_11_12,
   I2 => M_reg_11_16,
   I3 => M_reg_11_27,
   I4 => M_reg_10_9,
   O => W_26_11_i_11_n_0
);
W_26_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_10_9,
   I1 => x114_out_9,
   I2 => M_reg_11_27,
   I3 => M_reg_11_16,
   I4 => M_reg_11_12,
   O => W_26_11_i_12_n_0
);
W_26_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x114_out_8,
   I1 => M_reg_11_11,
   I2 => M_reg_11_15,
   I3 => M_reg_11_26,
   I4 => M_reg_10_8,
   O => W_26_11_i_13_n_0
);
W_26_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_10_8,
   I1 => x114_out_8,
   I2 => M_reg_11_26,
   I3 => M_reg_11_15,
   I4 => M_reg_11_11,
   O => W_26_11_i_14_n_0
);
W_26_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x114_out_7,
   I1 => M_reg_11_10,
   I2 => M_reg_11_14,
   I3 => M_reg_11_25,
   I4 => M_reg_10_7,
   O => W_26_11_i_15_n_0
);
W_26_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_10_7,
   I1 => x114_out_7,
   I2 => M_reg_11_25,
   I3 => M_reg_11_14,
   I4 => M_reg_11_10,
   O => W_26_11_i_16_n_0
);
W_26_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x114_out_6,
   I1 => M_reg_11_9,
   I2 => M_reg_11_13,
   I3 => M_reg_11_24,
   I4 => M_reg_10_6,
   O => W_26_11_i_17_n_0
);
W_26_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x108_out_20,
   I1 => x108_out_27,
   I2 => x108_out_29,
   I3 => W_26_11_i_10_n_0,
   I4 => W_26_11_i_11_n_0,
   O => W_26_11_i_2_n_0
);
W_26_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x108_out_19,
   I1 => x108_out_26,
   I2 => x108_out_28,
   I3 => W_26_11_i_12_n_0,
   I4 => W_26_11_i_13_n_0,
   O => W_26_11_i_3_n_0
);
W_26_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x108_out_18,
   I1 => x108_out_25,
   I2 => x108_out_27,
   I3 => W_26_11_i_14_n_0,
   I4 => W_26_11_i_15_n_0,
   O => W_26_11_i_4_n_0
);
W_26_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x108_out_17,
   I1 => x108_out_24,
   I2 => x108_out_26,
   I3 => W_26_11_i_16_n_0,
   I4 => W_26_11_i_17_n_0,
   O => W_26_11_i_5_n_0
);
W_26_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_26_11_i_2_n_0,
   I1 => W_26_15_i_16_n_0,
   I2 => x108_out_21,
   I3 => x108_out_28,
   I4 => x108_out_30,
   I5 => W_26_15_i_17_n_0,
   O => W_26_11_i_6_n_0
);
W_26_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_26_11_i_3_n_0,
   I1 => W_26_11_i_10_n_0,
   I2 => x108_out_20,
   I3 => x108_out_27,
   I4 => x108_out_29,
   I5 => W_26_11_i_11_n_0,
   O => W_26_11_i_7_n_0
);
W_26_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_26_11_i_4_n_0,
   I1 => W_26_11_i_12_n_0,
   I2 => x108_out_19,
   I3 => x108_out_26,
   I4 => x108_out_28,
   I5 => W_26_11_i_13_n_0,
   O => W_26_11_i_8_n_0
);
W_26_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_26_11_i_5_n_0,
   I1 => W_26_11_i_14_n_0,
   I2 => x108_out_18,
   I3 => x108_out_25,
   I4 => x108_out_27,
   I5 => W_26_11_i_15_n_0,
   O => W_26_11_i_9_n_0
);
W_26_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_10_14,
   I1 => x114_out_14,
   I2 => M_reg_11_0,
   I3 => M_reg_11_21,
   I4 => M_reg_11_17,
   O => W_26_15_i_10_n_0
);
W_26_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x114_out_13,
   I1 => M_reg_11_16,
   I2 => M_reg_11_20,
   I3 => M_reg_11_31,
   I4 => M_reg_10_13,
   O => W_26_15_i_11_n_0
);
W_26_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_10_13,
   I1 => x114_out_13,
   I2 => M_reg_11_31,
   I3 => M_reg_11_20,
   I4 => M_reg_11_16,
   O => W_26_15_i_12_n_0
);
W_26_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x114_out_12,
   I1 => M_reg_11_15,
   I2 => M_reg_11_19,
   I3 => M_reg_11_30,
   I4 => M_reg_10_12,
   O => W_26_15_i_13_n_0
);
W_26_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_10_12,
   I1 => x114_out_12,
   I2 => M_reg_11_30,
   I3 => M_reg_11_19,
   I4 => M_reg_11_15,
   O => W_26_15_i_14_n_0
);
W_26_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x114_out_11,
   I1 => M_reg_11_14,
   I2 => M_reg_11_18,
   I3 => M_reg_11_29,
   I4 => M_reg_10_11,
   O => W_26_15_i_15_n_0
);
W_26_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_10_11,
   I1 => x114_out_11,
   I2 => M_reg_11_29,
   I3 => M_reg_11_18,
   I4 => M_reg_11_14,
   O => W_26_15_i_16_n_0
);
W_26_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x114_out_10,
   I1 => M_reg_11_13,
   I2 => M_reg_11_17,
   I3 => M_reg_11_28,
   I4 => M_reg_10_10,
   O => W_26_15_i_17_n_0
);
W_26_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x108_out_24,
   I1 => x108_out_31,
   I2 => x108_out_1,
   I3 => W_26_15_i_10_n_0,
   I4 => W_26_15_i_11_n_0,
   O => W_26_15_i_2_n_0
);
W_26_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x108_out_23,
   I1 => x108_out_30,
   I2 => x108_out_0,
   I3 => W_26_15_i_12_n_0,
   I4 => W_26_15_i_13_n_0,
   O => W_26_15_i_3_n_0
);
W_26_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x108_out_22,
   I1 => x108_out_29,
   I2 => x108_out_31,
   I3 => W_26_15_i_14_n_0,
   I4 => W_26_15_i_15_n_0,
   O => W_26_15_i_4_n_0
);
W_26_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x108_out_21,
   I1 => x108_out_28,
   I2 => x108_out_30,
   I3 => W_26_15_i_16_n_0,
   I4 => W_26_15_i_17_n_0,
   O => W_26_15_i_5_n_0
);
W_26_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_26_15_i_2_n_0,
   I1 => W_26_19_i_16_n_0,
   I2 => x108_out_25,
   I3 => x108_out_0,
   I4 => x108_out_2,
   I5 => W_26_19_i_17_n_0,
   O => W_26_15_i_6_n_0
);
W_26_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_26_15_i_3_n_0,
   I1 => W_26_15_i_10_n_0,
   I2 => x108_out_24,
   I3 => x108_out_31,
   I4 => x108_out_1,
   I5 => W_26_15_i_11_n_0,
   O => W_26_15_i_7_n_0
);
W_26_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_26_15_i_4_n_0,
   I1 => W_26_15_i_12_n_0,
   I2 => x108_out_23,
   I3 => x108_out_30,
   I4 => x108_out_0,
   I5 => W_26_15_i_13_n_0,
   O => W_26_15_i_8_n_0
);
W_26_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_26_15_i_5_n_0,
   I1 => W_26_15_i_14_n_0,
   I2 => x108_out_22,
   I3 => x108_out_29,
   I4 => x108_out_31,
   I5 => W_26_15_i_15_n_0,
   O => W_26_15_i_9_n_0
);
W_26_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_10_18,
   I1 => x114_out_18,
   I2 => M_reg_11_4,
   I3 => M_reg_11_25,
   I4 => M_reg_11_21,
   O => W_26_19_i_10_n_0
);
W_26_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x114_out_17,
   I1 => M_reg_11_20,
   I2 => M_reg_11_24,
   I3 => M_reg_11_3,
   I4 => M_reg_10_17,
   O => W_26_19_i_11_n_0
);
W_26_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_10_17,
   I1 => x114_out_17,
   I2 => M_reg_11_3,
   I3 => M_reg_11_24,
   I4 => M_reg_11_20,
   O => W_26_19_i_12_n_0
);
W_26_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x114_out_16,
   I1 => M_reg_11_19,
   I2 => M_reg_11_23,
   I3 => M_reg_11_2,
   I4 => M_reg_10_16,
   O => W_26_19_i_13_n_0
);
W_26_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_10_16,
   I1 => x114_out_16,
   I2 => M_reg_11_2,
   I3 => M_reg_11_23,
   I4 => M_reg_11_19,
   O => W_26_19_i_14_n_0
);
W_26_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x114_out_15,
   I1 => M_reg_11_18,
   I2 => M_reg_11_22,
   I3 => M_reg_11_1,
   I4 => M_reg_10_15,
   O => W_26_19_i_15_n_0
);
W_26_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_10_15,
   I1 => x114_out_15,
   I2 => M_reg_11_1,
   I3 => M_reg_11_22,
   I4 => M_reg_11_18,
   O => W_26_19_i_16_n_0
);
W_26_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x114_out_14,
   I1 => M_reg_11_17,
   I2 => M_reg_11_21,
   I3 => M_reg_11_0,
   I4 => M_reg_10_14,
   O => W_26_19_i_17_n_0
);
W_26_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x108_out_28,
   I1 => x108_out_3,
   I2 => x108_out_5,
   I3 => W_26_19_i_10_n_0,
   I4 => W_26_19_i_11_n_0,
   O => W_26_19_i_2_n_0
);
W_26_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x108_out_27,
   I1 => x108_out_2,
   I2 => x108_out_4,
   I3 => W_26_19_i_12_n_0,
   I4 => W_26_19_i_13_n_0,
   O => W_26_19_i_3_n_0
);
W_26_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x108_out_26,
   I1 => x108_out_1,
   I2 => x108_out_3,
   I3 => W_26_19_i_14_n_0,
   I4 => W_26_19_i_15_n_0,
   O => W_26_19_i_4_n_0
);
W_26_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x108_out_25,
   I1 => x108_out_0,
   I2 => x108_out_2,
   I3 => W_26_19_i_16_n_0,
   I4 => W_26_19_i_17_n_0,
   O => W_26_19_i_5_n_0
);
W_26_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_26_19_i_2_n_0,
   I1 => W_26_23_i_16_n_0,
   I2 => x108_out_29,
   I3 => x108_out_4,
   I4 => x108_out_6,
   I5 => W_26_23_i_17_n_0,
   O => W_26_19_i_6_n_0
);
W_26_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_26_19_i_3_n_0,
   I1 => W_26_19_i_10_n_0,
   I2 => x108_out_28,
   I3 => x108_out_3,
   I4 => x108_out_5,
   I5 => W_26_19_i_11_n_0,
   O => W_26_19_i_7_n_0
);
W_26_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_26_19_i_4_n_0,
   I1 => W_26_19_i_12_n_0,
   I2 => x108_out_27,
   I3 => x108_out_2,
   I4 => x108_out_4,
   I5 => W_26_19_i_13_n_0,
   O => W_26_19_i_8_n_0
);
W_26_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_26_19_i_5_n_0,
   I1 => W_26_19_i_14_n_0,
   I2 => x108_out_26,
   I3 => x108_out_1,
   I4 => x108_out_3,
   I5 => W_26_19_i_15_n_0,
   O => W_26_19_i_9_n_0
);
W_26_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_10_22,
   I1 => x114_out_22,
   I2 => M_reg_11_8,
   I3 => M_reg_11_29,
   I4 => M_reg_11_25,
   O => W_26_23_i_10_n_0
);
W_26_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x114_out_21,
   I1 => M_reg_11_24,
   I2 => M_reg_11_28,
   I3 => M_reg_11_7,
   I4 => M_reg_10_21,
   O => W_26_23_i_11_n_0
);
W_26_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_10_21,
   I1 => x114_out_21,
   I2 => M_reg_11_7,
   I3 => M_reg_11_28,
   I4 => M_reg_11_24,
   O => W_26_23_i_12_n_0
);
W_26_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x114_out_20,
   I1 => M_reg_11_23,
   I2 => M_reg_11_27,
   I3 => M_reg_11_6,
   I4 => M_reg_10_20,
   O => W_26_23_i_13_n_0
);
W_26_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_10_20,
   I1 => x114_out_20,
   I2 => M_reg_11_6,
   I3 => M_reg_11_27,
   I4 => M_reg_11_23,
   O => W_26_23_i_14_n_0
);
W_26_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x114_out_19,
   I1 => M_reg_11_22,
   I2 => M_reg_11_26,
   I3 => M_reg_11_5,
   I4 => M_reg_10_19,
   O => W_26_23_i_15_n_0
);
W_26_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_10_19,
   I1 => x114_out_19,
   I2 => M_reg_11_5,
   I3 => M_reg_11_26,
   I4 => M_reg_11_22,
   O => W_26_23_i_16_n_0
);
W_26_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x114_out_18,
   I1 => M_reg_11_21,
   I2 => M_reg_11_25,
   I3 => M_reg_11_4,
   I4 => M_reg_10_18,
   O => W_26_23_i_17_n_0
);
W_26_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x108_out_7,
   I1 => x108_out_9,
   I2 => W_26_23_i_10_n_0,
   I3 => W_26_23_i_11_n_0,
   O => W_26_23_i_2_n_0
);
W_26_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x108_out_31,
   I1 => x108_out_6,
   I2 => x108_out_8,
   I3 => W_26_23_i_12_n_0,
   I4 => W_26_23_i_13_n_0,
   O => W_26_23_i_3_n_0
);
W_26_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x108_out_30,
   I1 => x108_out_5,
   I2 => x108_out_7,
   I3 => W_26_23_i_14_n_0,
   I4 => W_26_23_i_15_n_0,
   O => W_26_23_i_4_n_0
);
W_26_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x108_out_29,
   I1 => x108_out_4,
   I2 => x108_out_6,
   I3 => W_26_23_i_16_n_0,
   I4 => W_26_23_i_17_n_0,
   O => W_26_23_i_5_n_0
);
W_26_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x108_out_8,
   I1 => x108_out_10,
   I2 => W_26_27_i_16_n_0,
   I3 => W_26_27_i_17_n_0,
   I4 => W_26_23_i_2_n_0,
   O => W_26_23_i_6_n_0
);
W_26_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x108_out_7,
   I1 => x108_out_9,
   I2 => W_26_23_i_10_n_0,
   I3 => W_26_23_i_11_n_0,
   I4 => W_26_23_i_3_n_0,
   O => W_26_23_i_7_n_0
);
W_26_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_26_23_i_4_n_0,
   I1 => W_26_23_i_12_n_0,
   I2 => x108_out_31,
   I3 => x108_out_6,
   I4 => x108_out_8,
   I5 => W_26_23_i_13_n_0,
   O => W_26_23_i_8_n_0
);
W_26_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_26_23_i_5_n_0,
   I1 => W_26_23_i_14_n_0,
   I2 => x108_out_30,
   I3 => x108_out_5,
   I4 => x108_out_7,
   I5 => W_26_23_i_15_n_0,
   O => W_26_23_i_9_n_0
);
W_26_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_10_26,
   I1 => x114_out_26,
   I2 => M_reg_11_12,
   I3 => M_reg_11_1,
   I4 => M_reg_11_29,
   O => W_26_27_i_10_n_0
);
W_26_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x114_out_25,
   I1 => M_reg_11_28,
   I2 => M_reg_11_0,
   I3 => M_reg_11_11,
   I4 => M_reg_10_25,
   O => W_26_27_i_11_n_0
);
W_26_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_10_25,
   I1 => x114_out_25,
   I2 => M_reg_11_11,
   I3 => M_reg_11_0,
   I4 => M_reg_11_28,
   O => W_26_27_i_12_n_0
);
W_26_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x114_out_24,
   I1 => M_reg_11_27,
   I2 => M_reg_11_31,
   I3 => M_reg_11_10,
   I4 => M_reg_10_24,
   O => W_26_27_i_13_n_0
);
W_26_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_10_24,
   I1 => x114_out_24,
   I2 => M_reg_11_10,
   I3 => M_reg_11_31,
   I4 => M_reg_11_27,
   O => W_26_27_i_14_n_0
);
W_26_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x114_out_23,
   I1 => M_reg_11_26,
   I2 => M_reg_11_30,
   I3 => M_reg_11_9,
   I4 => M_reg_10_23,
   O => W_26_27_i_15_n_0
);
W_26_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_10_23,
   I1 => x114_out_23,
   I2 => M_reg_11_9,
   I3 => M_reg_11_30,
   I4 => M_reg_11_26,
   O => W_26_27_i_16_n_0
);
W_26_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x114_out_22,
   I1 => M_reg_11_25,
   I2 => M_reg_11_29,
   I3 => M_reg_11_8,
   I4 => M_reg_10_22,
   O => W_26_27_i_17_n_0
);
W_26_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x108_out_11,
   I1 => x108_out_13,
   I2 => W_26_27_i_10_n_0,
   I3 => W_26_27_i_11_n_0,
   O => W_26_27_i_2_n_0
);
W_26_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x108_out_10,
   I1 => x108_out_12,
   I2 => W_26_27_i_12_n_0,
   I3 => W_26_27_i_13_n_0,
   O => W_26_27_i_3_n_0
);
W_26_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x108_out_9,
   I1 => x108_out_11,
   I2 => W_26_27_i_14_n_0,
   I3 => W_26_27_i_15_n_0,
   O => W_26_27_i_4_n_0
);
W_26_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x108_out_8,
   I1 => x108_out_10,
   I2 => W_26_27_i_16_n_0,
   I3 => W_26_27_i_17_n_0,
   O => W_26_27_i_5_n_0
);
W_26_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x108_out_12,
   I1 => x108_out_14,
   I2 => W_26_31_i_13_n_0,
   I3 => W_26_31_i_14_n_0,
   I4 => W_26_27_i_2_n_0,
   O => W_26_27_i_6_n_0
);
W_26_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x108_out_11,
   I1 => x108_out_13,
   I2 => W_26_27_i_10_n_0,
   I3 => W_26_27_i_11_n_0,
   I4 => W_26_27_i_3_n_0,
   O => W_26_27_i_7_n_0
);
W_26_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x108_out_10,
   I1 => x108_out_12,
   I2 => W_26_27_i_12_n_0,
   I3 => W_26_27_i_13_n_0,
   I4 => W_26_27_i_4_n_0,
   O => W_26_27_i_8_n_0
);
W_26_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x108_out_9,
   I1 => x108_out_11,
   I2 => W_26_27_i_14_n_0,
   I3 => W_26_27_i_15_n_0,
   I4 => W_26_27_i_5_n_0,
   O => W_26_27_i_9_n_0
);
W_26_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x114_out_28,
   I1 => M_reg_11_31,
   I2 => M_reg_11_3,
   I3 => M_reg_11_14,
   I4 => M_reg_10_28,
   O => W_26_31_i_10_n_0
);
W_26_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_10_28,
   I1 => x114_out_28,
   I2 => M_reg_11_14,
   I3 => M_reg_11_3,
   I4 => M_reg_11_31,
   O => W_26_31_i_11_n_0
);
W_26_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x114_out_27,
   I1 => M_reg_11_30,
   I2 => M_reg_11_2,
   I3 => M_reg_11_13,
   I4 => M_reg_10_27,
   O => W_26_31_i_12_n_0
);
W_26_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_10_27,
   I1 => x114_out_27,
   I2 => M_reg_11_13,
   I3 => M_reg_11_2,
   I4 => M_reg_11_30,
   O => W_26_31_i_13_n_0
);
W_26_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x114_out_26,
   I1 => M_reg_11_29,
   I2 => M_reg_11_1,
   I3 => M_reg_11_12,
   I4 => M_reg_10_26,
   O => W_26_31_i_14_n_0
);
W_26_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x114_out_29,
   I1 => M_reg_11_4,
   I2 => M_reg_11_15,
   I3 => M_reg_10_29,
   O => W_26_31_i_15_n_0
);
W_26_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x108_out_17,
   I1 => x108_out_15,
   O => SIGMA_LCASE_1307_out_0_30
);
W_26_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => M_reg_11_6,
   I1 => M_reg_11_17,
   I2 => x114_out_31,
   I3 => M_reg_10_31,
   I4 => x108_out_16,
   I5 => x108_out_18,
   O => W_26_31_i_17_n_0
);
W_26_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => M_reg_11_16,
   I1 => M_reg_11_5,
   O => SIGMA_LCASE_0303_out_30
);
W_26_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => M_reg_10_30,
   I1 => x114_out_30,
   I2 => M_reg_11_16,
   I3 => M_reg_11_5,
   O => W_26_31_i_19_n_0
);
W_26_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x108_out_14,
   I1 => x108_out_16,
   I2 => W_26_31_i_9_n_0,
   I3 => W_26_31_i_10_n_0,
   O => W_26_31_i_2_n_0
);
W_26_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x108_out_13,
   I1 => x108_out_15,
   I2 => W_26_31_i_11_n_0,
   I3 => W_26_31_i_12_n_0,
   O => W_26_31_i_3_n_0
);
W_26_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x108_out_12,
   I1 => x108_out_14,
   I2 => W_26_31_i_13_n_0,
   I3 => W_26_31_i_14_n_0,
   O => W_26_31_i_4_n_0
);
W_26_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_26_31_i_15_n_0,
   I1 => SIGMA_LCASE_1307_out_0_30,
   I2 => W_26_31_i_17_n_0,
   I3 => x114_out_30,
   I4 => SIGMA_LCASE_0303_out_30,
   I5 => M_reg_10_30,
   O => W_26_31_i_5_n_0
);
W_26_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_26_31_i_2_n_0,
   I1 => W_26_31_i_19_n_0,
   I2 => x108_out_15,
   I3 => x108_out_17,
   I4 => W_26_31_i_15_n_0,
   O => W_26_31_i_6_n_0
);
W_26_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x108_out_14,
   I1 => x108_out_16,
   I2 => W_26_31_i_9_n_0,
   I3 => W_26_31_i_10_n_0,
   I4 => W_26_31_i_3_n_0,
   O => W_26_31_i_7_n_0
);
W_26_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x108_out_13,
   I1 => x108_out_15,
   I2 => W_26_31_i_11_n_0,
   I3 => W_26_31_i_12_n_0,
   I4 => W_26_31_i_4_n_0,
   O => W_26_31_i_8_n_0
);
W_26_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => M_reg_10_29,
   I1 => x114_out_29,
   I2 => M_reg_11_15,
   I3 => M_reg_11_4,
   O => W_26_31_i_9_n_0
);
W_26_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_10_2,
   I1 => x114_out_2,
   I2 => M_reg_11_20,
   I3 => M_reg_11_9,
   I4 => M_reg_11_5,
   O => W_26_3_i_10_n_0
);
W_26_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x114_out_1,
   I1 => M_reg_11_4,
   I2 => M_reg_11_8,
   I3 => M_reg_11_19,
   I4 => M_reg_10_1,
   O => W_26_3_i_11_n_0
);
W_26_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => M_reg_11_19,
   I1 => M_reg_11_8,
   I2 => M_reg_11_4,
   O => SIGMA_LCASE_0303_out_1
);
W_26_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x108_out_21,
   I1 => x108_out_19,
   I2 => x108_out_12,
   O => SIGMA_LCASE_1307_out_0_2
);
W_26_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x108_out_20,
   I1 => x108_out_18,
   I2 => x108_out_11,
   O => SIGMA_LCASE_1307_out_1
);
W_26_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x108_out_12,
   I1 => x108_out_19,
   I2 => x108_out_21,
   I3 => W_26_3_i_10_n_0,
   I4 => W_26_3_i_11_n_0,
   O => W_26_3_i_2_n_0
);
W_26_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_26_3_i_11_n_0,
   I1 => x108_out_21,
   I2 => x108_out_19,
   I3 => x108_out_12,
   I4 => W_26_3_i_10_n_0,
   O => W_26_3_i_3_n_0
);
W_26_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_0303_out_1,
   I1 => x114_out_1,
   I2 => M_reg_10_1,
   I3 => x108_out_11,
   I4 => x108_out_18,
   I5 => x108_out_20,
   O => W_26_3_i_4_n_0
);
W_26_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_10_0,
   I1 => x114_out_0,
   I2 => M_reg_11_18,
   I3 => M_reg_11_7,
   I4 => M_reg_11_3,
   O => W_26_3_i_5_n_0
);
W_26_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_26_3_i_2_n_0,
   I1 => W_26_7_i_16_n_0,
   I2 => x108_out_13,
   I3 => x108_out_20,
   I4 => x108_out_22,
   I5 => W_26_7_i_17_n_0,
   O => W_26_3_i_6_n_0
);
W_26_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_26_3_i_10_n_0,
   I1 => SIGMA_LCASE_1307_out_0_2,
   I2 => M_reg_10_1,
   I3 => x114_out_1,
   I4 => SIGMA_LCASE_0303_out_1,
   I5 => SIGMA_LCASE_1307_out_1,
   O => W_26_3_i_7_n_0
);
W_26_3_i_8 : LUT6
  generic map(
   INIT => X"566565566aa6a66a"
  )
 port map (
   I0 => W_26_3_i_4_n_0,
   I1 => M_reg_10_0,
   I2 => M_reg_11_18,
   I3 => M_reg_11_7,
   I4 => M_reg_11_3,
   I5 => x114_out_0,
   O => W_26_3_i_8_n_0
);
W_26_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_26_3_i_5_n_0,
   I1 => x108_out_10,
   I2 => x108_out_17,
   I3 => x108_out_19,
   O => W_26_3_i_9_n_0
);
W_26_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_10_6,
   I1 => x114_out_6,
   I2 => M_reg_11_24,
   I3 => M_reg_11_13,
   I4 => M_reg_11_9,
   O => W_26_7_i_10_n_0
);
W_26_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x114_out_5,
   I1 => M_reg_11_8,
   I2 => M_reg_11_12,
   I3 => M_reg_11_23,
   I4 => M_reg_10_5,
   O => W_26_7_i_11_n_0
);
W_26_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_10_5,
   I1 => x114_out_5,
   I2 => M_reg_11_23,
   I3 => M_reg_11_12,
   I4 => M_reg_11_8,
   O => W_26_7_i_12_n_0
);
W_26_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x114_out_4,
   I1 => M_reg_11_7,
   I2 => M_reg_11_11,
   I3 => M_reg_11_22,
   I4 => M_reg_10_4,
   O => W_26_7_i_13_n_0
);
W_26_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_10_4,
   I1 => x114_out_4,
   I2 => M_reg_11_22,
   I3 => M_reg_11_11,
   I4 => M_reg_11_7,
   O => W_26_7_i_14_n_0
);
W_26_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x114_out_3,
   I1 => M_reg_11_6,
   I2 => M_reg_11_10,
   I3 => M_reg_11_21,
   I4 => M_reg_10_3,
   O => W_26_7_i_15_n_0
);
W_26_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_10_3,
   I1 => x114_out_3,
   I2 => M_reg_11_21,
   I3 => M_reg_11_10,
   I4 => M_reg_11_6,
   O => W_26_7_i_16_n_0
);
W_26_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x114_out_2,
   I1 => M_reg_11_5,
   I2 => M_reg_11_9,
   I3 => M_reg_11_20,
   I4 => M_reg_10_2,
   O => W_26_7_i_17_n_0
);
W_26_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x108_out_16,
   I1 => x108_out_23,
   I2 => x108_out_25,
   I3 => W_26_7_i_10_n_0,
   I4 => W_26_7_i_11_n_0,
   O => W_26_7_i_2_n_0
);
W_26_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x108_out_15,
   I1 => x108_out_22,
   I2 => x108_out_24,
   I3 => W_26_7_i_12_n_0,
   I4 => W_26_7_i_13_n_0,
   O => W_26_7_i_3_n_0
);
W_26_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x108_out_14,
   I1 => x108_out_21,
   I2 => x108_out_23,
   I3 => W_26_7_i_14_n_0,
   I4 => W_26_7_i_15_n_0,
   O => W_26_7_i_4_n_0
);
W_26_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x108_out_13,
   I1 => x108_out_20,
   I2 => x108_out_22,
   I3 => W_26_7_i_16_n_0,
   I4 => W_26_7_i_17_n_0,
   O => W_26_7_i_5_n_0
);
W_26_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_26_7_i_2_n_0,
   I1 => W_26_11_i_16_n_0,
   I2 => x108_out_17,
   I3 => x108_out_24,
   I4 => x108_out_26,
   I5 => W_26_11_i_17_n_0,
   O => W_26_7_i_6_n_0
);
W_26_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_26_7_i_3_n_0,
   I1 => W_26_7_i_10_n_0,
   I2 => x108_out_16,
   I3 => x108_out_23,
   I4 => x108_out_25,
   I5 => W_26_7_i_11_n_0,
   O => W_26_7_i_7_n_0
);
W_26_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_26_7_i_4_n_0,
   I1 => W_26_7_i_12_n_0,
   I2 => x108_out_15,
   I3 => x108_out_22,
   I4 => x108_out_24,
   I5 => W_26_7_i_13_n_0,
   O => W_26_7_i_8_n_0
);
W_26_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_26_7_i_5_n_0,
   I1 => W_26_7_i_14_n_0,
   I2 => x108_out_14,
   I3 => x108_out_21,
   I4 => x108_out_23,
   I5 => W_26_7_i_15_n_0,
   O => W_26_7_i_9_n_0
);
W_27_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_11_10,
   I1 => x113_out_10,
   I2 => M_reg_12_28,
   I3 => M_reg_12_17,
   I4 => M_reg_12_13,
   O => W_27_11_i_10_n_0
);
W_27_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x113_out_9,
   I1 => M_reg_12_12,
   I2 => M_reg_12_16,
   I3 => M_reg_12_27,
   I4 => M_reg_11_9,
   O => W_27_11_i_11_n_0
);
W_27_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_11_9,
   I1 => x113_out_9,
   I2 => M_reg_12_27,
   I3 => M_reg_12_16,
   I4 => M_reg_12_12,
   O => W_27_11_i_12_n_0
);
W_27_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x113_out_8,
   I1 => M_reg_12_11,
   I2 => M_reg_12_15,
   I3 => M_reg_12_26,
   I4 => M_reg_11_8,
   O => W_27_11_i_13_n_0
);
W_27_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_11_8,
   I1 => x113_out_8,
   I2 => M_reg_12_26,
   I3 => M_reg_12_15,
   I4 => M_reg_12_11,
   O => W_27_11_i_14_n_0
);
W_27_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x113_out_7,
   I1 => M_reg_12_10,
   I2 => M_reg_12_14,
   I3 => M_reg_12_25,
   I4 => M_reg_11_7,
   O => W_27_11_i_15_n_0
);
W_27_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_11_7,
   I1 => x113_out_7,
   I2 => M_reg_12_25,
   I3 => M_reg_12_14,
   I4 => M_reg_12_10,
   O => W_27_11_i_16_n_0
);
W_27_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x113_out_6,
   I1 => M_reg_12_9,
   I2 => M_reg_12_13,
   I3 => M_reg_12_24,
   I4 => M_reg_11_6,
   O => W_27_11_i_17_n_0
);
W_27_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x106_out_20,
   I1 => x106_out_27,
   I2 => x106_out_29,
   I3 => W_27_11_i_10_n_0,
   I4 => W_27_11_i_11_n_0,
   O => W_27_11_i_2_n_0
);
W_27_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x106_out_19,
   I1 => x106_out_26,
   I2 => x106_out_28,
   I3 => W_27_11_i_12_n_0,
   I4 => W_27_11_i_13_n_0,
   O => W_27_11_i_3_n_0
);
W_27_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x106_out_18,
   I1 => x106_out_25,
   I2 => x106_out_27,
   I3 => W_27_11_i_14_n_0,
   I4 => W_27_11_i_15_n_0,
   O => W_27_11_i_4_n_0
);
W_27_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x106_out_17,
   I1 => x106_out_24,
   I2 => x106_out_26,
   I3 => W_27_11_i_16_n_0,
   I4 => W_27_11_i_17_n_0,
   O => W_27_11_i_5_n_0
);
W_27_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_27_11_i_2_n_0,
   I1 => W_27_15_i_16_n_0,
   I2 => x106_out_21,
   I3 => x106_out_28,
   I4 => x106_out_30,
   I5 => W_27_15_i_17_n_0,
   O => W_27_11_i_6_n_0
);
W_27_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_27_11_i_3_n_0,
   I1 => W_27_11_i_10_n_0,
   I2 => x106_out_20,
   I3 => x106_out_27,
   I4 => x106_out_29,
   I5 => W_27_11_i_11_n_0,
   O => W_27_11_i_7_n_0
);
W_27_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_27_11_i_4_n_0,
   I1 => W_27_11_i_12_n_0,
   I2 => x106_out_19,
   I3 => x106_out_26,
   I4 => x106_out_28,
   I5 => W_27_11_i_13_n_0,
   O => W_27_11_i_8_n_0
);
W_27_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_27_11_i_5_n_0,
   I1 => W_27_11_i_14_n_0,
   I2 => x106_out_18,
   I3 => x106_out_25,
   I4 => x106_out_27,
   I5 => W_27_11_i_15_n_0,
   O => W_27_11_i_9_n_0
);
W_27_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_11_14,
   I1 => x113_out_14,
   I2 => M_reg_12_0,
   I3 => M_reg_12_21,
   I4 => M_reg_12_17,
   O => W_27_15_i_10_n_0
);
W_27_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x113_out_13,
   I1 => M_reg_12_16,
   I2 => M_reg_12_20,
   I3 => M_reg_12_31,
   I4 => M_reg_11_13,
   O => W_27_15_i_11_n_0
);
W_27_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_11_13,
   I1 => x113_out_13,
   I2 => M_reg_12_31,
   I3 => M_reg_12_20,
   I4 => M_reg_12_16,
   O => W_27_15_i_12_n_0
);
W_27_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x113_out_12,
   I1 => M_reg_12_15,
   I2 => M_reg_12_19,
   I3 => M_reg_12_30,
   I4 => M_reg_11_12,
   O => W_27_15_i_13_n_0
);
W_27_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_11_12,
   I1 => x113_out_12,
   I2 => M_reg_12_30,
   I3 => M_reg_12_19,
   I4 => M_reg_12_15,
   O => W_27_15_i_14_n_0
);
W_27_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x113_out_11,
   I1 => M_reg_12_14,
   I2 => M_reg_12_18,
   I3 => M_reg_12_29,
   I4 => M_reg_11_11,
   O => W_27_15_i_15_n_0
);
W_27_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_11_11,
   I1 => x113_out_11,
   I2 => M_reg_12_29,
   I3 => M_reg_12_18,
   I4 => M_reg_12_14,
   O => W_27_15_i_16_n_0
);
W_27_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x113_out_10,
   I1 => M_reg_12_13,
   I2 => M_reg_12_17,
   I3 => M_reg_12_28,
   I4 => M_reg_11_10,
   O => W_27_15_i_17_n_0
);
W_27_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x106_out_24,
   I1 => x106_out_31,
   I2 => x106_out_1,
   I3 => W_27_15_i_10_n_0,
   I4 => W_27_15_i_11_n_0,
   O => W_27_15_i_2_n_0
);
W_27_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x106_out_23,
   I1 => x106_out_30,
   I2 => x106_out_0,
   I3 => W_27_15_i_12_n_0,
   I4 => W_27_15_i_13_n_0,
   O => W_27_15_i_3_n_0
);
W_27_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x106_out_22,
   I1 => x106_out_29,
   I2 => x106_out_31,
   I3 => W_27_15_i_14_n_0,
   I4 => W_27_15_i_15_n_0,
   O => W_27_15_i_4_n_0
);
W_27_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x106_out_21,
   I1 => x106_out_28,
   I2 => x106_out_30,
   I3 => W_27_15_i_16_n_0,
   I4 => W_27_15_i_17_n_0,
   O => W_27_15_i_5_n_0
);
W_27_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_27_15_i_2_n_0,
   I1 => W_27_19_i_16_n_0,
   I2 => x106_out_25,
   I3 => x106_out_0,
   I4 => x106_out_2,
   I5 => W_27_19_i_17_n_0,
   O => W_27_15_i_6_n_0
);
W_27_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_27_15_i_3_n_0,
   I1 => W_27_15_i_10_n_0,
   I2 => x106_out_24,
   I3 => x106_out_31,
   I4 => x106_out_1,
   I5 => W_27_15_i_11_n_0,
   O => W_27_15_i_7_n_0
);
W_27_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_27_15_i_4_n_0,
   I1 => W_27_15_i_12_n_0,
   I2 => x106_out_23,
   I3 => x106_out_30,
   I4 => x106_out_0,
   I5 => W_27_15_i_13_n_0,
   O => W_27_15_i_8_n_0
);
W_27_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_27_15_i_5_n_0,
   I1 => W_27_15_i_14_n_0,
   I2 => x106_out_22,
   I3 => x106_out_29,
   I4 => x106_out_31,
   I5 => W_27_15_i_15_n_0,
   O => W_27_15_i_9_n_0
);
W_27_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_11_18,
   I1 => x113_out_18,
   I2 => M_reg_12_4,
   I3 => M_reg_12_25,
   I4 => M_reg_12_21,
   O => W_27_19_i_10_n_0
);
W_27_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x113_out_17,
   I1 => M_reg_12_20,
   I2 => M_reg_12_24,
   I3 => M_reg_12_3,
   I4 => M_reg_11_17,
   O => W_27_19_i_11_n_0
);
W_27_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_11_17,
   I1 => x113_out_17,
   I2 => M_reg_12_3,
   I3 => M_reg_12_24,
   I4 => M_reg_12_20,
   O => W_27_19_i_12_n_0
);
W_27_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x113_out_16,
   I1 => M_reg_12_19,
   I2 => M_reg_12_23,
   I3 => M_reg_12_2,
   I4 => M_reg_11_16,
   O => W_27_19_i_13_n_0
);
W_27_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_11_16,
   I1 => x113_out_16,
   I2 => M_reg_12_2,
   I3 => M_reg_12_23,
   I4 => M_reg_12_19,
   O => W_27_19_i_14_n_0
);
W_27_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x113_out_15,
   I1 => M_reg_12_18,
   I2 => M_reg_12_22,
   I3 => M_reg_12_1,
   I4 => M_reg_11_15,
   O => W_27_19_i_15_n_0
);
W_27_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_11_15,
   I1 => x113_out_15,
   I2 => M_reg_12_1,
   I3 => M_reg_12_22,
   I4 => M_reg_12_18,
   O => W_27_19_i_16_n_0
);
W_27_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x113_out_14,
   I1 => M_reg_12_17,
   I2 => M_reg_12_21,
   I3 => M_reg_12_0,
   I4 => M_reg_11_14,
   O => W_27_19_i_17_n_0
);
W_27_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x106_out_28,
   I1 => x106_out_3,
   I2 => x106_out_5,
   I3 => W_27_19_i_10_n_0,
   I4 => W_27_19_i_11_n_0,
   O => W_27_19_i_2_n_0
);
W_27_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x106_out_27,
   I1 => x106_out_2,
   I2 => x106_out_4,
   I3 => W_27_19_i_12_n_0,
   I4 => W_27_19_i_13_n_0,
   O => W_27_19_i_3_n_0
);
W_27_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x106_out_26,
   I1 => x106_out_1,
   I2 => x106_out_3,
   I3 => W_27_19_i_14_n_0,
   I4 => W_27_19_i_15_n_0,
   O => W_27_19_i_4_n_0
);
W_27_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x106_out_25,
   I1 => x106_out_0,
   I2 => x106_out_2,
   I3 => W_27_19_i_16_n_0,
   I4 => W_27_19_i_17_n_0,
   O => W_27_19_i_5_n_0
);
W_27_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_27_19_i_2_n_0,
   I1 => W_27_23_i_16_n_0,
   I2 => x106_out_29,
   I3 => x106_out_4,
   I4 => x106_out_6,
   I5 => W_27_23_i_17_n_0,
   O => W_27_19_i_6_n_0
);
W_27_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_27_19_i_3_n_0,
   I1 => W_27_19_i_10_n_0,
   I2 => x106_out_28,
   I3 => x106_out_3,
   I4 => x106_out_5,
   I5 => W_27_19_i_11_n_0,
   O => W_27_19_i_7_n_0
);
W_27_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_27_19_i_4_n_0,
   I1 => W_27_19_i_12_n_0,
   I2 => x106_out_27,
   I3 => x106_out_2,
   I4 => x106_out_4,
   I5 => W_27_19_i_13_n_0,
   O => W_27_19_i_8_n_0
);
W_27_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_27_19_i_5_n_0,
   I1 => W_27_19_i_14_n_0,
   I2 => x106_out_26,
   I3 => x106_out_1,
   I4 => x106_out_3,
   I5 => W_27_19_i_15_n_0,
   O => W_27_19_i_9_n_0
);
W_27_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_11_22,
   I1 => x113_out_22,
   I2 => M_reg_12_8,
   I3 => M_reg_12_29,
   I4 => M_reg_12_25,
   O => W_27_23_i_10_n_0
);
W_27_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x113_out_21,
   I1 => M_reg_12_24,
   I2 => M_reg_12_28,
   I3 => M_reg_12_7,
   I4 => M_reg_11_21,
   O => W_27_23_i_11_n_0
);
W_27_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_11_21,
   I1 => x113_out_21,
   I2 => M_reg_12_7,
   I3 => M_reg_12_28,
   I4 => M_reg_12_24,
   O => W_27_23_i_12_n_0
);
W_27_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x113_out_20,
   I1 => M_reg_12_23,
   I2 => M_reg_12_27,
   I3 => M_reg_12_6,
   I4 => M_reg_11_20,
   O => W_27_23_i_13_n_0
);
W_27_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_11_20,
   I1 => x113_out_20,
   I2 => M_reg_12_6,
   I3 => M_reg_12_27,
   I4 => M_reg_12_23,
   O => W_27_23_i_14_n_0
);
W_27_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x113_out_19,
   I1 => M_reg_12_22,
   I2 => M_reg_12_26,
   I3 => M_reg_12_5,
   I4 => M_reg_11_19,
   O => W_27_23_i_15_n_0
);
W_27_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_11_19,
   I1 => x113_out_19,
   I2 => M_reg_12_5,
   I3 => M_reg_12_26,
   I4 => M_reg_12_22,
   O => W_27_23_i_16_n_0
);
W_27_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x113_out_18,
   I1 => M_reg_12_21,
   I2 => M_reg_12_25,
   I3 => M_reg_12_4,
   I4 => M_reg_11_18,
   O => W_27_23_i_17_n_0
);
W_27_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x106_out_7,
   I1 => x106_out_9,
   I2 => W_27_23_i_10_n_0,
   I3 => W_27_23_i_11_n_0,
   O => W_27_23_i_2_n_0
);
W_27_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x106_out_31,
   I1 => x106_out_6,
   I2 => x106_out_8,
   I3 => W_27_23_i_12_n_0,
   I4 => W_27_23_i_13_n_0,
   O => W_27_23_i_3_n_0
);
W_27_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x106_out_30,
   I1 => x106_out_5,
   I2 => x106_out_7,
   I3 => W_27_23_i_14_n_0,
   I4 => W_27_23_i_15_n_0,
   O => W_27_23_i_4_n_0
);
W_27_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x106_out_29,
   I1 => x106_out_4,
   I2 => x106_out_6,
   I3 => W_27_23_i_16_n_0,
   I4 => W_27_23_i_17_n_0,
   O => W_27_23_i_5_n_0
);
W_27_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x106_out_8,
   I1 => x106_out_10,
   I2 => W_27_27_i_16_n_0,
   I3 => W_27_27_i_17_n_0,
   I4 => W_27_23_i_2_n_0,
   O => W_27_23_i_6_n_0
);
W_27_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x106_out_7,
   I1 => x106_out_9,
   I2 => W_27_23_i_10_n_0,
   I3 => W_27_23_i_11_n_0,
   I4 => W_27_23_i_3_n_0,
   O => W_27_23_i_7_n_0
);
W_27_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_27_23_i_4_n_0,
   I1 => W_27_23_i_12_n_0,
   I2 => x106_out_31,
   I3 => x106_out_6,
   I4 => x106_out_8,
   I5 => W_27_23_i_13_n_0,
   O => W_27_23_i_8_n_0
);
W_27_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_27_23_i_5_n_0,
   I1 => W_27_23_i_14_n_0,
   I2 => x106_out_30,
   I3 => x106_out_5,
   I4 => x106_out_7,
   I5 => W_27_23_i_15_n_0,
   O => W_27_23_i_9_n_0
);
W_27_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_11_26,
   I1 => x113_out_26,
   I2 => M_reg_12_12,
   I3 => M_reg_12_1,
   I4 => M_reg_12_29,
   O => W_27_27_i_10_n_0
);
W_27_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x113_out_25,
   I1 => M_reg_12_28,
   I2 => M_reg_12_0,
   I3 => M_reg_12_11,
   I4 => M_reg_11_25,
   O => W_27_27_i_11_n_0
);
W_27_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_11_25,
   I1 => x113_out_25,
   I2 => M_reg_12_11,
   I3 => M_reg_12_0,
   I4 => M_reg_12_28,
   O => W_27_27_i_12_n_0
);
W_27_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x113_out_24,
   I1 => M_reg_12_27,
   I2 => M_reg_12_31,
   I3 => M_reg_12_10,
   I4 => M_reg_11_24,
   O => W_27_27_i_13_n_0
);
W_27_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_11_24,
   I1 => x113_out_24,
   I2 => M_reg_12_10,
   I3 => M_reg_12_31,
   I4 => M_reg_12_27,
   O => W_27_27_i_14_n_0
);
W_27_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x113_out_23,
   I1 => M_reg_12_26,
   I2 => M_reg_12_30,
   I3 => M_reg_12_9,
   I4 => M_reg_11_23,
   O => W_27_27_i_15_n_0
);
W_27_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_11_23,
   I1 => x113_out_23,
   I2 => M_reg_12_9,
   I3 => M_reg_12_30,
   I4 => M_reg_12_26,
   O => W_27_27_i_16_n_0
);
W_27_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x113_out_22,
   I1 => M_reg_12_25,
   I2 => M_reg_12_29,
   I3 => M_reg_12_8,
   I4 => M_reg_11_22,
   O => W_27_27_i_17_n_0
);
W_27_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x106_out_11,
   I1 => x106_out_13,
   I2 => W_27_27_i_10_n_0,
   I3 => W_27_27_i_11_n_0,
   O => W_27_27_i_2_n_0
);
W_27_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x106_out_10,
   I1 => x106_out_12,
   I2 => W_27_27_i_12_n_0,
   I3 => W_27_27_i_13_n_0,
   O => W_27_27_i_3_n_0
);
W_27_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x106_out_9,
   I1 => x106_out_11,
   I2 => W_27_27_i_14_n_0,
   I3 => W_27_27_i_15_n_0,
   O => W_27_27_i_4_n_0
);
W_27_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x106_out_8,
   I1 => x106_out_10,
   I2 => W_27_27_i_16_n_0,
   I3 => W_27_27_i_17_n_0,
   O => W_27_27_i_5_n_0
);
W_27_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x106_out_12,
   I1 => x106_out_14,
   I2 => W_27_31_i_13_n_0,
   I3 => W_27_31_i_14_n_0,
   I4 => W_27_27_i_2_n_0,
   O => W_27_27_i_6_n_0
);
W_27_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x106_out_11,
   I1 => x106_out_13,
   I2 => W_27_27_i_10_n_0,
   I3 => W_27_27_i_11_n_0,
   I4 => W_27_27_i_3_n_0,
   O => W_27_27_i_7_n_0
);
W_27_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x106_out_10,
   I1 => x106_out_12,
   I2 => W_27_27_i_12_n_0,
   I3 => W_27_27_i_13_n_0,
   I4 => W_27_27_i_4_n_0,
   O => W_27_27_i_8_n_0
);
W_27_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x106_out_9,
   I1 => x106_out_11,
   I2 => W_27_27_i_14_n_0,
   I3 => W_27_27_i_15_n_0,
   I4 => W_27_27_i_5_n_0,
   O => W_27_27_i_9_n_0
);
W_27_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x113_out_28,
   I1 => M_reg_12_31,
   I2 => M_reg_12_3,
   I3 => M_reg_12_14,
   I4 => M_reg_11_28,
   O => W_27_31_i_10_n_0
);
W_27_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_11_28,
   I1 => x113_out_28,
   I2 => M_reg_12_14,
   I3 => M_reg_12_3,
   I4 => M_reg_12_31,
   O => W_27_31_i_11_n_0
);
W_27_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x113_out_27,
   I1 => M_reg_12_30,
   I2 => M_reg_12_2,
   I3 => M_reg_12_13,
   I4 => M_reg_11_27,
   O => W_27_31_i_12_n_0
);
W_27_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_11_27,
   I1 => x113_out_27,
   I2 => M_reg_12_13,
   I3 => M_reg_12_2,
   I4 => M_reg_12_30,
   O => W_27_31_i_13_n_0
);
W_27_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x113_out_26,
   I1 => M_reg_12_29,
   I2 => M_reg_12_1,
   I3 => M_reg_12_12,
   I4 => M_reg_11_26,
   O => W_27_31_i_14_n_0
);
W_27_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x113_out_29,
   I1 => M_reg_12_4,
   I2 => M_reg_12_15,
   I3 => M_reg_11_29,
   O => W_27_31_i_15_n_0
);
W_27_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x106_out_17,
   I1 => x106_out_15,
   O => SIGMA_LCASE_1299_out_0_30
);
W_27_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => M_reg_12_6,
   I1 => M_reg_12_17,
   I2 => x113_out_31,
   I3 => M_reg_11_31,
   I4 => x106_out_16,
   I5 => x106_out_18,
   O => W_27_31_i_17_n_0
);
W_27_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => M_reg_12_16,
   I1 => M_reg_12_5,
   O => SIGMA_LCASE_0295_out_30
);
W_27_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => M_reg_11_30,
   I1 => x113_out_30,
   I2 => M_reg_12_16,
   I3 => M_reg_12_5,
   O => W_27_31_i_19_n_0
);
W_27_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x106_out_14,
   I1 => x106_out_16,
   I2 => W_27_31_i_9_n_0,
   I3 => W_27_31_i_10_n_0,
   O => W_27_31_i_2_n_0
);
W_27_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x106_out_13,
   I1 => x106_out_15,
   I2 => W_27_31_i_11_n_0,
   I3 => W_27_31_i_12_n_0,
   O => W_27_31_i_3_n_0
);
W_27_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x106_out_12,
   I1 => x106_out_14,
   I2 => W_27_31_i_13_n_0,
   I3 => W_27_31_i_14_n_0,
   O => W_27_31_i_4_n_0
);
W_27_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_27_31_i_15_n_0,
   I1 => SIGMA_LCASE_1299_out_0_30,
   I2 => W_27_31_i_17_n_0,
   I3 => x113_out_30,
   I4 => SIGMA_LCASE_0295_out_30,
   I5 => M_reg_11_30,
   O => W_27_31_i_5_n_0
);
W_27_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_27_31_i_2_n_0,
   I1 => W_27_31_i_19_n_0,
   I2 => x106_out_15,
   I3 => x106_out_17,
   I4 => W_27_31_i_15_n_0,
   O => W_27_31_i_6_n_0
);
W_27_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x106_out_14,
   I1 => x106_out_16,
   I2 => W_27_31_i_9_n_0,
   I3 => W_27_31_i_10_n_0,
   I4 => W_27_31_i_3_n_0,
   O => W_27_31_i_7_n_0
);
W_27_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x106_out_13,
   I1 => x106_out_15,
   I2 => W_27_31_i_11_n_0,
   I3 => W_27_31_i_12_n_0,
   I4 => W_27_31_i_4_n_0,
   O => W_27_31_i_8_n_0
);
W_27_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => M_reg_11_29,
   I1 => x113_out_29,
   I2 => M_reg_12_15,
   I3 => M_reg_12_4,
   O => W_27_31_i_9_n_0
);
W_27_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_11_2,
   I1 => x113_out_2,
   I2 => M_reg_12_20,
   I3 => M_reg_12_9,
   I4 => M_reg_12_5,
   O => W_27_3_i_10_n_0
);
W_27_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x113_out_1,
   I1 => M_reg_12_4,
   I2 => M_reg_12_8,
   I3 => M_reg_12_19,
   I4 => M_reg_11_1,
   O => W_27_3_i_11_n_0
);
W_27_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => M_reg_12_19,
   I1 => M_reg_12_8,
   I2 => M_reg_12_4,
   O => SIGMA_LCASE_0295_out_1
);
W_27_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x106_out_21,
   I1 => x106_out_19,
   I2 => x106_out_12,
   O => SIGMA_LCASE_1299_out_0_2
);
W_27_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x106_out_20,
   I1 => x106_out_18,
   I2 => x106_out_11,
   O => SIGMA_LCASE_1299_out_1
);
W_27_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x106_out_12,
   I1 => x106_out_19,
   I2 => x106_out_21,
   I3 => W_27_3_i_10_n_0,
   I4 => W_27_3_i_11_n_0,
   O => W_27_3_i_2_n_0
);
W_27_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_27_3_i_11_n_0,
   I1 => x106_out_21,
   I2 => x106_out_19,
   I3 => x106_out_12,
   I4 => W_27_3_i_10_n_0,
   O => W_27_3_i_3_n_0
);
W_27_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_0295_out_1,
   I1 => x113_out_1,
   I2 => M_reg_11_1,
   I3 => x106_out_11,
   I4 => x106_out_18,
   I5 => x106_out_20,
   O => W_27_3_i_4_n_0
);
W_27_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_11_0,
   I1 => x113_out_0,
   I2 => M_reg_12_18,
   I3 => M_reg_12_7,
   I4 => M_reg_12_3,
   O => W_27_3_i_5_n_0
);
W_27_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_27_3_i_2_n_0,
   I1 => W_27_7_i_16_n_0,
   I2 => x106_out_13,
   I3 => x106_out_20,
   I4 => x106_out_22,
   I5 => W_27_7_i_17_n_0,
   O => W_27_3_i_6_n_0
);
W_27_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_27_3_i_10_n_0,
   I1 => SIGMA_LCASE_1299_out_0_2,
   I2 => M_reg_11_1,
   I3 => x113_out_1,
   I4 => SIGMA_LCASE_0295_out_1,
   I5 => SIGMA_LCASE_1299_out_1,
   O => W_27_3_i_7_n_0
);
W_27_3_i_8 : LUT6
  generic map(
   INIT => X"566565566aa6a66a"
  )
 port map (
   I0 => W_27_3_i_4_n_0,
   I1 => M_reg_11_0,
   I2 => M_reg_12_18,
   I3 => M_reg_12_7,
   I4 => M_reg_12_3,
   I5 => x113_out_0,
   O => W_27_3_i_8_n_0
);
W_27_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_27_3_i_5_n_0,
   I1 => x106_out_10,
   I2 => x106_out_17,
   I3 => x106_out_19,
   O => W_27_3_i_9_n_0
);
W_27_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_11_6,
   I1 => x113_out_6,
   I2 => M_reg_12_24,
   I3 => M_reg_12_13,
   I4 => M_reg_12_9,
   O => W_27_7_i_10_n_0
);
W_27_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x113_out_5,
   I1 => M_reg_12_8,
   I2 => M_reg_12_12,
   I3 => M_reg_12_23,
   I4 => M_reg_11_5,
   O => W_27_7_i_11_n_0
);
W_27_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_11_5,
   I1 => x113_out_5,
   I2 => M_reg_12_23,
   I3 => M_reg_12_12,
   I4 => M_reg_12_8,
   O => W_27_7_i_12_n_0
);
W_27_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x113_out_4,
   I1 => M_reg_12_7,
   I2 => M_reg_12_11,
   I3 => M_reg_12_22,
   I4 => M_reg_11_4,
   O => W_27_7_i_13_n_0
);
W_27_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_11_4,
   I1 => x113_out_4,
   I2 => M_reg_12_22,
   I3 => M_reg_12_11,
   I4 => M_reg_12_7,
   O => W_27_7_i_14_n_0
);
W_27_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x113_out_3,
   I1 => M_reg_12_6,
   I2 => M_reg_12_10,
   I3 => M_reg_12_21,
   I4 => M_reg_11_3,
   O => W_27_7_i_15_n_0
);
W_27_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_11_3,
   I1 => x113_out_3,
   I2 => M_reg_12_21,
   I3 => M_reg_12_10,
   I4 => M_reg_12_6,
   O => W_27_7_i_16_n_0
);
W_27_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x113_out_2,
   I1 => M_reg_12_5,
   I2 => M_reg_12_9,
   I3 => M_reg_12_20,
   I4 => M_reg_11_2,
   O => W_27_7_i_17_n_0
);
W_27_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x106_out_16,
   I1 => x106_out_23,
   I2 => x106_out_25,
   I3 => W_27_7_i_10_n_0,
   I4 => W_27_7_i_11_n_0,
   O => W_27_7_i_2_n_0
);
W_27_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x106_out_15,
   I1 => x106_out_22,
   I2 => x106_out_24,
   I3 => W_27_7_i_12_n_0,
   I4 => W_27_7_i_13_n_0,
   O => W_27_7_i_3_n_0
);
W_27_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x106_out_14,
   I1 => x106_out_21,
   I2 => x106_out_23,
   I3 => W_27_7_i_14_n_0,
   I4 => W_27_7_i_15_n_0,
   O => W_27_7_i_4_n_0
);
W_27_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x106_out_13,
   I1 => x106_out_20,
   I2 => x106_out_22,
   I3 => W_27_7_i_16_n_0,
   I4 => W_27_7_i_17_n_0,
   O => W_27_7_i_5_n_0
);
W_27_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_27_7_i_2_n_0,
   I1 => W_27_11_i_16_n_0,
   I2 => x106_out_17,
   I3 => x106_out_24,
   I4 => x106_out_26,
   I5 => W_27_11_i_17_n_0,
   O => W_27_7_i_6_n_0
);
W_27_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_27_7_i_3_n_0,
   I1 => W_27_7_i_10_n_0,
   I2 => x106_out_16,
   I3 => x106_out_23,
   I4 => x106_out_25,
   I5 => W_27_7_i_11_n_0,
   O => W_27_7_i_7_n_0
);
W_27_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_27_7_i_4_n_0,
   I1 => W_27_7_i_12_n_0,
   I2 => x106_out_15,
   I3 => x106_out_22,
   I4 => x106_out_24,
   I5 => W_27_7_i_13_n_0,
   O => W_27_7_i_8_n_0
);
W_27_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_27_7_i_5_n_0,
   I1 => W_27_7_i_14_n_0,
   I2 => x106_out_14,
   I3 => x106_out_21,
   I4 => x106_out_23,
   I5 => W_27_7_i_15_n_0,
   O => W_27_7_i_9_n_0
);
W_28_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_12_10,
   I1 => x112_out_10,
   I2 => M_reg_13_28,
   I3 => M_reg_13_17,
   I4 => M_reg_13_13,
   O => W_28_11_i_10_n_0
);
W_28_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x112_out_9,
   I1 => M_reg_13_12,
   I2 => M_reg_13_16,
   I3 => M_reg_13_27,
   I4 => M_reg_12_9,
   O => W_28_11_i_11_n_0
);
W_28_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_12_9,
   I1 => x112_out_9,
   I2 => M_reg_13_27,
   I3 => M_reg_13_16,
   I4 => M_reg_13_12,
   O => W_28_11_i_12_n_0
);
W_28_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x112_out_8,
   I1 => M_reg_13_11,
   I2 => M_reg_13_15,
   I3 => M_reg_13_26,
   I4 => M_reg_12_8,
   O => W_28_11_i_13_n_0
);
W_28_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_12_8,
   I1 => x112_out_8,
   I2 => M_reg_13_26,
   I3 => M_reg_13_15,
   I4 => M_reg_13_11,
   O => W_28_11_i_14_n_0
);
W_28_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x112_out_7,
   I1 => M_reg_13_10,
   I2 => M_reg_13_14,
   I3 => M_reg_13_25,
   I4 => M_reg_12_7,
   O => W_28_11_i_15_n_0
);
W_28_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_12_7,
   I1 => x112_out_7,
   I2 => M_reg_13_25,
   I3 => M_reg_13_14,
   I4 => M_reg_13_10,
   O => W_28_11_i_16_n_0
);
W_28_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x112_out_6,
   I1 => M_reg_13_9,
   I2 => M_reg_13_13,
   I3 => M_reg_13_24,
   I4 => M_reg_12_6,
   O => W_28_11_i_17_n_0
);
W_28_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x104_out_20,
   I1 => x104_out_27,
   I2 => x104_out_29,
   I3 => W_28_11_i_10_n_0,
   I4 => W_28_11_i_11_n_0,
   O => W_28_11_i_2_n_0
);
W_28_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x104_out_19,
   I1 => x104_out_26,
   I2 => x104_out_28,
   I3 => W_28_11_i_12_n_0,
   I4 => W_28_11_i_13_n_0,
   O => W_28_11_i_3_n_0
);
W_28_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x104_out_18,
   I1 => x104_out_25,
   I2 => x104_out_27,
   I3 => W_28_11_i_14_n_0,
   I4 => W_28_11_i_15_n_0,
   O => W_28_11_i_4_n_0
);
W_28_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x104_out_17,
   I1 => x104_out_24,
   I2 => x104_out_26,
   I3 => W_28_11_i_16_n_0,
   I4 => W_28_11_i_17_n_0,
   O => W_28_11_i_5_n_0
);
W_28_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_28_11_i_2_n_0,
   I1 => W_28_15_i_16_n_0,
   I2 => x104_out_21,
   I3 => x104_out_28,
   I4 => x104_out_30,
   I5 => W_28_15_i_17_n_0,
   O => W_28_11_i_6_n_0
);
W_28_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_28_11_i_3_n_0,
   I1 => W_28_11_i_10_n_0,
   I2 => x104_out_20,
   I3 => x104_out_27,
   I4 => x104_out_29,
   I5 => W_28_11_i_11_n_0,
   O => W_28_11_i_7_n_0
);
W_28_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_28_11_i_4_n_0,
   I1 => W_28_11_i_12_n_0,
   I2 => x104_out_19,
   I3 => x104_out_26,
   I4 => x104_out_28,
   I5 => W_28_11_i_13_n_0,
   O => W_28_11_i_8_n_0
);
W_28_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_28_11_i_5_n_0,
   I1 => W_28_11_i_14_n_0,
   I2 => x104_out_18,
   I3 => x104_out_25,
   I4 => x104_out_27,
   I5 => W_28_11_i_15_n_0,
   O => W_28_11_i_9_n_0
);
W_28_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_12_14,
   I1 => x112_out_14,
   I2 => M_reg_13_0,
   I3 => M_reg_13_21,
   I4 => M_reg_13_17,
   O => W_28_15_i_10_n_0
);
W_28_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x112_out_13,
   I1 => M_reg_13_16,
   I2 => M_reg_13_20,
   I3 => M_reg_13_31,
   I4 => M_reg_12_13,
   O => W_28_15_i_11_n_0
);
W_28_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_12_13,
   I1 => x112_out_13,
   I2 => M_reg_13_31,
   I3 => M_reg_13_20,
   I4 => M_reg_13_16,
   O => W_28_15_i_12_n_0
);
W_28_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x112_out_12,
   I1 => M_reg_13_15,
   I2 => M_reg_13_19,
   I3 => M_reg_13_30,
   I4 => M_reg_12_12,
   O => W_28_15_i_13_n_0
);
W_28_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_12_12,
   I1 => x112_out_12,
   I2 => M_reg_13_30,
   I3 => M_reg_13_19,
   I4 => M_reg_13_15,
   O => W_28_15_i_14_n_0
);
W_28_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x112_out_11,
   I1 => M_reg_13_14,
   I2 => M_reg_13_18,
   I3 => M_reg_13_29,
   I4 => M_reg_12_11,
   O => W_28_15_i_15_n_0
);
W_28_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_12_11,
   I1 => x112_out_11,
   I2 => M_reg_13_29,
   I3 => M_reg_13_18,
   I4 => M_reg_13_14,
   O => W_28_15_i_16_n_0
);
W_28_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x112_out_10,
   I1 => M_reg_13_13,
   I2 => M_reg_13_17,
   I3 => M_reg_13_28,
   I4 => M_reg_12_10,
   O => W_28_15_i_17_n_0
);
W_28_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x104_out_24,
   I1 => x104_out_31,
   I2 => x104_out_1,
   I3 => W_28_15_i_10_n_0,
   I4 => W_28_15_i_11_n_0,
   O => W_28_15_i_2_n_0
);
W_28_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x104_out_23,
   I1 => x104_out_30,
   I2 => x104_out_0,
   I3 => W_28_15_i_12_n_0,
   I4 => W_28_15_i_13_n_0,
   O => W_28_15_i_3_n_0
);
W_28_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x104_out_22,
   I1 => x104_out_29,
   I2 => x104_out_31,
   I3 => W_28_15_i_14_n_0,
   I4 => W_28_15_i_15_n_0,
   O => W_28_15_i_4_n_0
);
W_28_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x104_out_21,
   I1 => x104_out_28,
   I2 => x104_out_30,
   I3 => W_28_15_i_16_n_0,
   I4 => W_28_15_i_17_n_0,
   O => W_28_15_i_5_n_0
);
W_28_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_28_15_i_2_n_0,
   I1 => W_28_19_i_16_n_0,
   I2 => x104_out_25,
   I3 => x104_out_0,
   I4 => x104_out_2,
   I5 => W_28_19_i_17_n_0,
   O => W_28_15_i_6_n_0
);
W_28_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_28_15_i_3_n_0,
   I1 => W_28_15_i_10_n_0,
   I2 => x104_out_24,
   I3 => x104_out_31,
   I4 => x104_out_1,
   I5 => W_28_15_i_11_n_0,
   O => W_28_15_i_7_n_0
);
W_28_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_28_15_i_4_n_0,
   I1 => W_28_15_i_12_n_0,
   I2 => x104_out_23,
   I3 => x104_out_30,
   I4 => x104_out_0,
   I5 => W_28_15_i_13_n_0,
   O => W_28_15_i_8_n_0
);
W_28_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_28_15_i_5_n_0,
   I1 => W_28_15_i_14_n_0,
   I2 => x104_out_22,
   I3 => x104_out_29,
   I4 => x104_out_31,
   I5 => W_28_15_i_15_n_0,
   O => W_28_15_i_9_n_0
);
W_28_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_12_18,
   I1 => x112_out_18,
   I2 => M_reg_13_4,
   I3 => M_reg_13_25,
   I4 => M_reg_13_21,
   O => W_28_19_i_10_n_0
);
W_28_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x112_out_17,
   I1 => M_reg_13_20,
   I2 => M_reg_13_24,
   I3 => M_reg_13_3,
   I4 => M_reg_12_17,
   O => W_28_19_i_11_n_0
);
W_28_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_12_17,
   I1 => x112_out_17,
   I2 => M_reg_13_3,
   I3 => M_reg_13_24,
   I4 => M_reg_13_20,
   O => W_28_19_i_12_n_0
);
W_28_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x112_out_16,
   I1 => M_reg_13_19,
   I2 => M_reg_13_23,
   I3 => M_reg_13_2,
   I4 => M_reg_12_16,
   O => W_28_19_i_13_n_0
);
W_28_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_12_16,
   I1 => x112_out_16,
   I2 => M_reg_13_2,
   I3 => M_reg_13_23,
   I4 => M_reg_13_19,
   O => W_28_19_i_14_n_0
);
W_28_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x112_out_15,
   I1 => M_reg_13_18,
   I2 => M_reg_13_22,
   I3 => M_reg_13_1,
   I4 => M_reg_12_15,
   O => W_28_19_i_15_n_0
);
W_28_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_12_15,
   I1 => x112_out_15,
   I2 => M_reg_13_1,
   I3 => M_reg_13_22,
   I4 => M_reg_13_18,
   O => W_28_19_i_16_n_0
);
W_28_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x112_out_14,
   I1 => M_reg_13_17,
   I2 => M_reg_13_21,
   I3 => M_reg_13_0,
   I4 => M_reg_12_14,
   O => W_28_19_i_17_n_0
);
W_28_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x104_out_28,
   I1 => x104_out_3,
   I2 => x104_out_5,
   I3 => W_28_19_i_10_n_0,
   I4 => W_28_19_i_11_n_0,
   O => W_28_19_i_2_n_0
);
W_28_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x104_out_27,
   I1 => x104_out_2,
   I2 => x104_out_4,
   I3 => W_28_19_i_12_n_0,
   I4 => W_28_19_i_13_n_0,
   O => W_28_19_i_3_n_0
);
W_28_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x104_out_26,
   I1 => x104_out_1,
   I2 => x104_out_3,
   I3 => W_28_19_i_14_n_0,
   I4 => W_28_19_i_15_n_0,
   O => W_28_19_i_4_n_0
);
W_28_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x104_out_25,
   I1 => x104_out_0,
   I2 => x104_out_2,
   I3 => W_28_19_i_16_n_0,
   I4 => W_28_19_i_17_n_0,
   O => W_28_19_i_5_n_0
);
W_28_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_28_19_i_2_n_0,
   I1 => W_28_23_i_16_n_0,
   I2 => x104_out_29,
   I3 => x104_out_4,
   I4 => x104_out_6,
   I5 => W_28_23_i_17_n_0,
   O => W_28_19_i_6_n_0
);
W_28_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_28_19_i_3_n_0,
   I1 => W_28_19_i_10_n_0,
   I2 => x104_out_28,
   I3 => x104_out_3,
   I4 => x104_out_5,
   I5 => W_28_19_i_11_n_0,
   O => W_28_19_i_7_n_0
);
W_28_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_28_19_i_4_n_0,
   I1 => W_28_19_i_12_n_0,
   I2 => x104_out_27,
   I3 => x104_out_2,
   I4 => x104_out_4,
   I5 => W_28_19_i_13_n_0,
   O => W_28_19_i_8_n_0
);
W_28_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_28_19_i_5_n_0,
   I1 => W_28_19_i_14_n_0,
   I2 => x104_out_26,
   I3 => x104_out_1,
   I4 => x104_out_3,
   I5 => W_28_19_i_15_n_0,
   O => W_28_19_i_9_n_0
);
W_28_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_12_22,
   I1 => x112_out_22,
   I2 => M_reg_13_8,
   I3 => M_reg_13_29,
   I4 => M_reg_13_25,
   O => W_28_23_i_10_n_0
);
W_28_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x112_out_21,
   I1 => M_reg_13_24,
   I2 => M_reg_13_28,
   I3 => M_reg_13_7,
   I4 => M_reg_12_21,
   O => W_28_23_i_11_n_0
);
W_28_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_12_21,
   I1 => x112_out_21,
   I2 => M_reg_13_7,
   I3 => M_reg_13_28,
   I4 => M_reg_13_24,
   O => W_28_23_i_12_n_0
);
W_28_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x112_out_20,
   I1 => M_reg_13_23,
   I2 => M_reg_13_27,
   I3 => M_reg_13_6,
   I4 => M_reg_12_20,
   O => W_28_23_i_13_n_0
);
W_28_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_12_20,
   I1 => x112_out_20,
   I2 => M_reg_13_6,
   I3 => M_reg_13_27,
   I4 => M_reg_13_23,
   O => W_28_23_i_14_n_0
);
W_28_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x112_out_19,
   I1 => M_reg_13_22,
   I2 => M_reg_13_26,
   I3 => M_reg_13_5,
   I4 => M_reg_12_19,
   O => W_28_23_i_15_n_0
);
W_28_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_12_19,
   I1 => x112_out_19,
   I2 => M_reg_13_5,
   I3 => M_reg_13_26,
   I4 => M_reg_13_22,
   O => W_28_23_i_16_n_0
);
W_28_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x112_out_18,
   I1 => M_reg_13_21,
   I2 => M_reg_13_25,
   I3 => M_reg_13_4,
   I4 => M_reg_12_18,
   O => W_28_23_i_17_n_0
);
W_28_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x104_out_7,
   I1 => x104_out_9,
   I2 => W_28_23_i_10_n_0,
   I3 => W_28_23_i_11_n_0,
   O => W_28_23_i_2_n_0
);
W_28_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x104_out_31,
   I1 => x104_out_6,
   I2 => x104_out_8,
   I3 => W_28_23_i_12_n_0,
   I4 => W_28_23_i_13_n_0,
   O => W_28_23_i_3_n_0
);
W_28_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x104_out_30,
   I1 => x104_out_5,
   I2 => x104_out_7,
   I3 => W_28_23_i_14_n_0,
   I4 => W_28_23_i_15_n_0,
   O => W_28_23_i_4_n_0
);
W_28_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x104_out_29,
   I1 => x104_out_4,
   I2 => x104_out_6,
   I3 => W_28_23_i_16_n_0,
   I4 => W_28_23_i_17_n_0,
   O => W_28_23_i_5_n_0
);
W_28_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x104_out_8,
   I1 => x104_out_10,
   I2 => W_28_27_i_16_n_0,
   I3 => W_28_27_i_17_n_0,
   I4 => W_28_23_i_2_n_0,
   O => W_28_23_i_6_n_0
);
W_28_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x104_out_7,
   I1 => x104_out_9,
   I2 => W_28_23_i_10_n_0,
   I3 => W_28_23_i_11_n_0,
   I4 => W_28_23_i_3_n_0,
   O => W_28_23_i_7_n_0
);
W_28_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_28_23_i_4_n_0,
   I1 => W_28_23_i_12_n_0,
   I2 => x104_out_31,
   I3 => x104_out_6,
   I4 => x104_out_8,
   I5 => W_28_23_i_13_n_0,
   O => W_28_23_i_8_n_0
);
W_28_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_28_23_i_5_n_0,
   I1 => W_28_23_i_14_n_0,
   I2 => x104_out_30,
   I3 => x104_out_5,
   I4 => x104_out_7,
   I5 => W_28_23_i_15_n_0,
   O => W_28_23_i_9_n_0
);
W_28_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_12_26,
   I1 => x112_out_26,
   I2 => M_reg_13_12,
   I3 => M_reg_13_1,
   I4 => M_reg_13_29,
   O => W_28_27_i_10_n_0
);
W_28_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x112_out_25,
   I1 => M_reg_13_28,
   I2 => M_reg_13_0,
   I3 => M_reg_13_11,
   I4 => M_reg_12_25,
   O => W_28_27_i_11_n_0
);
W_28_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_12_25,
   I1 => x112_out_25,
   I2 => M_reg_13_11,
   I3 => M_reg_13_0,
   I4 => M_reg_13_28,
   O => W_28_27_i_12_n_0
);
W_28_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x112_out_24,
   I1 => M_reg_13_27,
   I2 => M_reg_13_31,
   I3 => M_reg_13_10,
   I4 => M_reg_12_24,
   O => W_28_27_i_13_n_0
);
W_28_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_12_24,
   I1 => x112_out_24,
   I2 => M_reg_13_10,
   I3 => M_reg_13_31,
   I4 => M_reg_13_27,
   O => W_28_27_i_14_n_0
);
W_28_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x112_out_23,
   I1 => M_reg_13_26,
   I2 => M_reg_13_30,
   I3 => M_reg_13_9,
   I4 => M_reg_12_23,
   O => W_28_27_i_15_n_0
);
W_28_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_12_23,
   I1 => x112_out_23,
   I2 => M_reg_13_9,
   I3 => M_reg_13_30,
   I4 => M_reg_13_26,
   O => W_28_27_i_16_n_0
);
W_28_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x112_out_22,
   I1 => M_reg_13_25,
   I2 => M_reg_13_29,
   I3 => M_reg_13_8,
   I4 => M_reg_12_22,
   O => W_28_27_i_17_n_0
);
W_28_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x104_out_11,
   I1 => x104_out_13,
   I2 => W_28_27_i_10_n_0,
   I3 => W_28_27_i_11_n_0,
   O => W_28_27_i_2_n_0
);
W_28_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x104_out_10,
   I1 => x104_out_12,
   I2 => W_28_27_i_12_n_0,
   I3 => W_28_27_i_13_n_0,
   O => W_28_27_i_3_n_0
);
W_28_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x104_out_9,
   I1 => x104_out_11,
   I2 => W_28_27_i_14_n_0,
   I3 => W_28_27_i_15_n_0,
   O => W_28_27_i_4_n_0
);
W_28_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x104_out_8,
   I1 => x104_out_10,
   I2 => W_28_27_i_16_n_0,
   I3 => W_28_27_i_17_n_0,
   O => W_28_27_i_5_n_0
);
W_28_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x104_out_12,
   I1 => x104_out_14,
   I2 => W_28_31_i_13_n_0,
   I3 => W_28_31_i_14_n_0,
   I4 => W_28_27_i_2_n_0,
   O => W_28_27_i_6_n_0
);
W_28_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x104_out_11,
   I1 => x104_out_13,
   I2 => W_28_27_i_10_n_0,
   I3 => W_28_27_i_11_n_0,
   I4 => W_28_27_i_3_n_0,
   O => W_28_27_i_7_n_0
);
W_28_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x104_out_10,
   I1 => x104_out_12,
   I2 => W_28_27_i_12_n_0,
   I3 => W_28_27_i_13_n_0,
   I4 => W_28_27_i_4_n_0,
   O => W_28_27_i_8_n_0
);
W_28_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x104_out_9,
   I1 => x104_out_11,
   I2 => W_28_27_i_14_n_0,
   I3 => W_28_27_i_15_n_0,
   I4 => W_28_27_i_5_n_0,
   O => W_28_27_i_9_n_0
);
W_28_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x112_out_28,
   I1 => M_reg_13_31,
   I2 => M_reg_13_3,
   I3 => M_reg_13_14,
   I4 => M_reg_12_28,
   O => W_28_31_i_10_n_0
);
W_28_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_12_28,
   I1 => x112_out_28,
   I2 => M_reg_13_14,
   I3 => M_reg_13_3,
   I4 => M_reg_13_31,
   O => W_28_31_i_11_n_0
);
W_28_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x112_out_27,
   I1 => M_reg_13_30,
   I2 => M_reg_13_2,
   I3 => M_reg_13_13,
   I4 => M_reg_12_27,
   O => W_28_31_i_12_n_0
);
W_28_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_12_27,
   I1 => x112_out_27,
   I2 => M_reg_13_13,
   I3 => M_reg_13_2,
   I4 => M_reg_13_30,
   O => W_28_31_i_13_n_0
);
W_28_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x112_out_26,
   I1 => M_reg_13_29,
   I2 => M_reg_13_1,
   I3 => M_reg_13_12,
   I4 => M_reg_12_26,
   O => W_28_31_i_14_n_0
);
W_28_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x112_out_29,
   I1 => M_reg_13_4,
   I2 => M_reg_13_15,
   I3 => M_reg_12_29,
   O => W_28_31_i_15_n_0
);
W_28_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x104_out_17,
   I1 => x104_out_15,
   O => SIGMA_LCASE_1291_out_0_30
);
W_28_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => M_reg_13_6,
   I1 => M_reg_13_17,
   I2 => x112_out_31,
   I3 => M_reg_12_31,
   I4 => x104_out_16,
   I5 => x104_out_18,
   O => W_28_31_i_17_n_0
);
W_28_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => M_reg_13_16,
   I1 => M_reg_13_5,
   O => SIGMA_LCASE_0287_out_30
);
W_28_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => M_reg_12_30,
   I1 => x112_out_30,
   I2 => M_reg_13_16,
   I3 => M_reg_13_5,
   O => W_28_31_i_19_n_0
);
W_28_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x104_out_14,
   I1 => x104_out_16,
   I2 => W_28_31_i_9_n_0,
   I3 => W_28_31_i_10_n_0,
   O => W_28_31_i_2_n_0
);
W_28_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x104_out_13,
   I1 => x104_out_15,
   I2 => W_28_31_i_11_n_0,
   I3 => W_28_31_i_12_n_0,
   O => W_28_31_i_3_n_0
);
W_28_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x104_out_12,
   I1 => x104_out_14,
   I2 => W_28_31_i_13_n_0,
   I3 => W_28_31_i_14_n_0,
   O => W_28_31_i_4_n_0
);
W_28_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_28_31_i_15_n_0,
   I1 => SIGMA_LCASE_1291_out_0_30,
   I2 => W_28_31_i_17_n_0,
   I3 => x112_out_30,
   I4 => SIGMA_LCASE_0287_out_30,
   I5 => M_reg_12_30,
   O => W_28_31_i_5_n_0
);
W_28_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_28_31_i_2_n_0,
   I1 => W_28_31_i_19_n_0,
   I2 => x104_out_15,
   I3 => x104_out_17,
   I4 => W_28_31_i_15_n_0,
   O => W_28_31_i_6_n_0
);
W_28_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x104_out_14,
   I1 => x104_out_16,
   I2 => W_28_31_i_9_n_0,
   I3 => W_28_31_i_10_n_0,
   I4 => W_28_31_i_3_n_0,
   O => W_28_31_i_7_n_0
);
W_28_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x104_out_13,
   I1 => x104_out_15,
   I2 => W_28_31_i_11_n_0,
   I3 => W_28_31_i_12_n_0,
   I4 => W_28_31_i_4_n_0,
   O => W_28_31_i_8_n_0
);
W_28_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => M_reg_12_29,
   I1 => x112_out_29,
   I2 => M_reg_13_15,
   I3 => M_reg_13_4,
   O => W_28_31_i_9_n_0
);
W_28_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_12_2,
   I1 => x112_out_2,
   I2 => M_reg_13_20,
   I3 => M_reg_13_9,
   I4 => M_reg_13_5,
   O => W_28_3_i_10_n_0
);
W_28_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x112_out_1,
   I1 => M_reg_13_4,
   I2 => M_reg_13_8,
   I3 => M_reg_13_19,
   I4 => M_reg_12_1,
   O => W_28_3_i_11_n_0
);
W_28_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => M_reg_13_19,
   I1 => M_reg_13_8,
   I2 => M_reg_13_4,
   O => SIGMA_LCASE_0287_out_1
);
W_28_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x104_out_21,
   I1 => x104_out_19,
   I2 => x104_out_12,
   O => SIGMA_LCASE_1291_out_0_2
);
W_28_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x104_out_20,
   I1 => x104_out_18,
   I2 => x104_out_11,
   O => SIGMA_LCASE_1291_out_1
);
W_28_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x104_out_12,
   I1 => x104_out_19,
   I2 => x104_out_21,
   I3 => W_28_3_i_10_n_0,
   I4 => W_28_3_i_11_n_0,
   O => W_28_3_i_2_n_0
);
W_28_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_28_3_i_11_n_0,
   I1 => x104_out_21,
   I2 => x104_out_19,
   I3 => x104_out_12,
   I4 => W_28_3_i_10_n_0,
   O => W_28_3_i_3_n_0
);
W_28_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_0287_out_1,
   I1 => x112_out_1,
   I2 => M_reg_12_1,
   I3 => x104_out_11,
   I4 => x104_out_18,
   I5 => x104_out_20,
   O => W_28_3_i_4_n_0
);
W_28_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_12_0,
   I1 => x112_out_0,
   I2 => M_reg_13_18,
   I3 => M_reg_13_7,
   I4 => M_reg_13_3,
   O => W_28_3_i_5_n_0
);
W_28_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_28_3_i_2_n_0,
   I1 => W_28_7_i_16_n_0,
   I2 => x104_out_13,
   I3 => x104_out_20,
   I4 => x104_out_22,
   I5 => W_28_7_i_17_n_0,
   O => W_28_3_i_6_n_0
);
W_28_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_28_3_i_10_n_0,
   I1 => SIGMA_LCASE_1291_out_0_2,
   I2 => M_reg_12_1,
   I3 => x112_out_1,
   I4 => SIGMA_LCASE_0287_out_1,
   I5 => SIGMA_LCASE_1291_out_1,
   O => W_28_3_i_7_n_0
);
W_28_3_i_8 : LUT6
  generic map(
   INIT => X"566565566aa6a66a"
  )
 port map (
   I0 => W_28_3_i_4_n_0,
   I1 => M_reg_12_0,
   I2 => M_reg_13_18,
   I3 => M_reg_13_7,
   I4 => M_reg_13_3,
   I5 => x112_out_0,
   O => W_28_3_i_8_n_0
);
W_28_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_28_3_i_5_n_0,
   I1 => x104_out_10,
   I2 => x104_out_17,
   I3 => x104_out_19,
   O => W_28_3_i_9_n_0
);
W_28_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_12_6,
   I1 => x112_out_6,
   I2 => M_reg_13_24,
   I3 => M_reg_13_13,
   I4 => M_reg_13_9,
   O => W_28_7_i_10_n_0
);
W_28_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x112_out_5,
   I1 => M_reg_13_8,
   I2 => M_reg_13_12,
   I3 => M_reg_13_23,
   I4 => M_reg_12_5,
   O => W_28_7_i_11_n_0
);
W_28_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_12_5,
   I1 => x112_out_5,
   I2 => M_reg_13_23,
   I3 => M_reg_13_12,
   I4 => M_reg_13_8,
   O => W_28_7_i_12_n_0
);
W_28_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x112_out_4,
   I1 => M_reg_13_7,
   I2 => M_reg_13_11,
   I3 => M_reg_13_22,
   I4 => M_reg_12_4,
   O => W_28_7_i_13_n_0
);
W_28_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_12_4,
   I1 => x112_out_4,
   I2 => M_reg_13_22,
   I3 => M_reg_13_11,
   I4 => M_reg_13_7,
   O => W_28_7_i_14_n_0
);
W_28_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x112_out_3,
   I1 => M_reg_13_6,
   I2 => M_reg_13_10,
   I3 => M_reg_13_21,
   I4 => M_reg_12_3,
   O => W_28_7_i_15_n_0
);
W_28_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_12_3,
   I1 => x112_out_3,
   I2 => M_reg_13_21,
   I3 => M_reg_13_10,
   I4 => M_reg_13_6,
   O => W_28_7_i_16_n_0
);
W_28_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x112_out_2,
   I1 => M_reg_13_5,
   I2 => M_reg_13_9,
   I3 => M_reg_13_20,
   I4 => M_reg_12_2,
   O => W_28_7_i_17_n_0
);
W_28_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x104_out_16,
   I1 => x104_out_23,
   I2 => x104_out_25,
   I3 => W_28_7_i_10_n_0,
   I4 => W_28_7_i_11_n_0,
   O => W_28_7_i_2_n_0
);
W_28_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x104_out_15,
   I1 => x104_out_22,
   I2 => x104_out_24,
   I3 => W_28_7_i_12_n_0,
   I4 => W_28_7_i_13_n_0,
   O => W_28_7_i_3_n_0
);
W_28_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x104_out_14,
   I1 => x104_out_21,
   I2 => x104_out_23,
   I3 => W_28_7_i_14_n_0,
   I4 => W_28_7_i_15_n_0,
   O => W_28_7_i_4_n_0
);
W_28_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x104_out_13,
   I1 => x104_out_20,
   I2 => x104_out_22,
   I3 => W_28_7_i_16_n_0,
   I4 => W_28_7_i_17_n_0,
   O => W_28_7_i_5_n_0
);
W_28_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_28_7_i_2_n_0,
   I1 => W_28_11_i_16_n_0,
   I2 => x104_out_17,
   I3 => x104_out_24,
   I4 => x104_out_26,
   I5 => W_28_11_i_17_n_0,
   O => W_28_7_i_6_n_0
);
W_28_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_28_7_i_3_n_0,
   I1 => W_28_7_i_10_n_0,
   I2 => x104_out_16,
   I3 => x104_out_23,
   I4 => x104_out_25,
   I5 => W_28_7_i_11_n_0,
   O => W_28_7_i_7_n_0
);
W_28_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_28_7_i_4_n_0,
   I1 => W_28_7_i_12_n_0,
   I2 => x104_out_15,
   I3 => x104_out_22,
   I4 => x104_out_24,
   I5 => W_28_7_i_13_n_0,
   O => W_28_7_i_8_n_0
);
W_28_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_28_7_i_5_n_0,
   I1 => W_28_7_i_14_n_0,
   I2 => x104_out_14,
   I3 => x104_out_21,
   I4 => x104_out_23,
   I5 => W_28_7_i_15_n_0,
   O => W_28_7_i_9_n_0
);
W_29_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_13_10,
   I1 => x111_out_10,
   I2 => M_reg_14_28,
   I3 => M_reg_14_17,
   I4 => M_reg_14_13,
   O => W_29_11_i_10_n_0
);
W_29_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x111_out_9,
   I1 => M_reg_14_12,
   I2 => M_reg_14_16,
   I3 => M_reg_14_27,
   I4 => M_reg_13_9,
   O => W_29_11_i_11_n_0
);
W_29_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_13_9,
   I1 => x111_out_9,
   I2 => M_reg_14_27,
   I3 => M_reg_14_16,
   I4 => M_reg_14_12,
   O => W_29_11_i_12_n_0
);
W_29_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x111_out_8,
   I1 => M_reg_14_11,
   I2 => M_reg_14_15,
   I3 => M_reg_14_26,
   I4 => M_reg_13_8,
   O => W_29_11_i_13_n_0
);
W_29_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_13_8,
   I1 => x111_out_8,
   I2 => M_reg_14_26,
   I3 => M_reg_14_15,
   I4 => M_reg_14_11,
   O => W_29_11_i_14_n_0
);
W_29_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x111_out_7,
   I1 => M_reg_14_10,
   I2 => M_reg_14_14,
   I3 => M_reg_14_25,
   I4 => M_reg_13_7,
   O => W_29_11_i_15_n_0
);
W_29_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_13_7,
   I1 => x111_out_7,
   I2 => M_reg_14_25,
   I3 => M_reg_14_14,
   I4 => M_reg_14_10,
   O => W_29_11_i_16_n_0
);
W_29_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x111_out_6,
   I1 => M_reg_14_9,
   I2 => M_reg_14_13,
   I3 => M_reg_14_24,
   I4 => M_reg_13_6,
   O => W_29_11_i_17_n_0
);
W_29_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x102_out_20,
   I1 => x102_out_27,
   I2 => x102_out_29,
   I3 => W_29_11_i_10_n_0,
   I4 => W_29_11_i_11_n_0,
   O => W_29_11_i_2_n_0
);
W_29_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x102_out_19,
   I1 => x102_out_26,
   I2 => x102_out_28,
   I3 => W_29_11_i_12_n_0,
   I4 => W_29_11_i_13_n_0,
   O => W_29_11_i_3_n_0
);
W_29_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x102_out_18,
   I1 => x102_out_25,
   I2 => x102_out_27,
   I3 => W_29_11_i_14_n_0,
   I4 => W_29_11_i_15_n_0,
   O => W_29_11_i_4_n_0
);
W_29_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x102_out_17,
   I1 => x102_out_24,
   I2 => x102_out_26,
   I3 => W_29_11_i_16_n_0,
   I4 => W_29_11_i_17_n_0,
   O => W_29_11_i_5_n_0
);
W_29_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_29_11_i_2_n_0,
   I1 => W_29_15_i_16_n_0,
   I2 => x102_out_21,
   I3 => x102_out_28,
   I4 => x102_out_30,
   I5 => W_29_15_i_17_n_0,
   O => W_29_11_i_6_n_0
);
W_29_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_29_11_i_3_n_0,
   I1 => W_29_11_i_10_n_0,
   I2 => x102_out_20,
   I3 => x102_out_27,
   I4 => x102_out_29,
   I5 => W_29_11_i_11_n_0,
   O => W_29_11_i_7_n_0
);
W_29_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_29_11_i_4_n_0,
   I1 => W_29_11_i_12_n_0,
   I2 => x102_out_19,
   I3 => x102_out_26,
   I4 => x102_out_28,
   I5 => W_29_11_i_13_n_0,
   O => W_29_11_i_8_n_0
);
W_29_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_29_11_i_5_n_0,
   I1 => W_29_11_i_14_n_0,
   I2 => x102_out_18,
   I3 => x102_out_25,
   I4 => x102_out_27,
   I5 => W_29_11_i_15_n_0,
   O => W_29_11_i_9_n_0
);
W_29_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_13_14,
   I1 => x111_out_14,
   I2 => M_reg_14_0,
   I3 => M_reg_14_21,
   I4 => M_reg_14_17,
   O => W_29_15_i_10_n_0
);
W_29_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x111_out_13,
   I1 => M_reg_14_16,
   I2 => M_reg_14_20,
   I3 => M_reg_14_31,
   I4 => M_reg_13_13,
   O => W_29_15_i_11_n_0
);
W_29_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_13_13,
   I1 => x111_out_13,
   I2 => M_reg_14_31,
   I3 => M_reg_14_20,
   I4 => M_reg_14_16,
   O => W_29_15_i_12_n_0
);
W_29_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x111_out_12,
   I1 => M_reg_14_15,
   I2 => M_reg_14_19,
   I3 => M_reg_14_30,
   I4 => M_reg_13_12,
   O => W_29_15_i_13_n_0
);
W_29_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_13_12,
   I1 => x111_out_12,
   I2 => M_reg_14_30,
   I3 => M_reg_14_19,
   I4 => M_reg_14_15,
   O => W_29_15_i_14_n_0
);
W_29_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x111_out_11,
   I1 => M_reg_14_14,
   I2 => M_reg_14_18,
   I3 => M_reg_14_29,
   I4 => M_reg_13_11,
   O => W_29_15_i_15_n_0
);
W_29_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_13_11,
   I1 => x111_out_11,
   I2 => M_reg_14_29,
   I3 => M_reg_14_18,
   I4 => M_reg_14_14,
   O => W_29_15_i_16_n_0
);
W_29_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x111_out_10,
   I1 => M_reg_14_13,
   I2 => M_reg_14_17,
   I3 => M_reg_14_28,
   I4 => M_reg_13_10,
   O => W_29_15_i_17_n_0
);
W_29_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x102_out_24,
   I1 => x102_out_31,
   I2 => x102_out_1,
   I3 => W_29_15_i_10_n_0,
   I4 => W_29_15_i_11_n_0,
   O => W_29_15_i_2_n_0
);
W_29_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x102_out_23,
   I1 => x102_out_30,
   I2 => x102_out_0,
   I3 => W_29_15_i_12_n_0,
   I4 => W_29_15_i_13_n_0,
   O => W_29_15_i_3_n_0
);
W_29_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x102_out_22,
   I1 => x102_out_29,
   I2 => x102_out_31,
   I3 => W_29_15_i_14_n_0,
   I4 => W_29_15_i_15_n_0,
   O => W_29_15_i_4_n_0
);
W_29_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x102_out_21,
   I1 => x102_out_28,
   I2 => x102_out_30,
   I3 => W_29_15_i_16_n_0,
   I4 => W_29_15_i_17_n_0,
   O => W_29_15_i_5_n_0
);
W_29_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_29_15_i_2_n_0,
   I1 => W_29_19_i_16_n_0,
   I2 => x102_out_25,
   I3 => x102_out_0,
   I4 => x102_out_2,
   I5 => W_29_19_i_17_n_0,
   O => W_29_15_i_6_n_0
);
W_29_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_29_15_i_3_n_0,
   I1 => W_29_15_i_10_n_0,
   I2 => x102_out_24,
   I3 => x102_out_31,
   I4 => x102_out_1,
   I5 => W_29_15_i_11_n_0,
   O => W_29_15_i_7_n_0
);
W_29_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_29_15_i_4_n_0,
   I1 => W_29_15_i_12_n_0,
   I2 => x102_out_23,
   I3 => x102_out_30,
   I4 => x102_out_0,
   I5 => W_29_15_i_13_n_0,
   O => W_29_15_i_8_n_0
);
W_29_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_29_15_i_5_n_0,
   I1 => W_29_15_i_14_n_0,
   I2 => x102_out_22,
   I3 => x102_out_29,
   I4 => x102_out_31,
   I5 => W_29_15_i_15_n_0,
   O => W_29_15_i_9_n_0
);
W_29_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_13_18,
   I1 => x111_out_18,
   I2 => M_reg_14_4,
   I3 => M_reg_14_25,
   I4 => M_reg_14_21,
   O => W_29_19_i_10_n_0
);
W_29_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x111_out_17,
   I1 => M_reg_14_20,
   I2 => M_reg_14_24,
   I3 => M_reg_14_3,
   I4 => M_reg_13_17,
   O => W_29_19_i_11_n_0
);
W_29_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_13_17,
   I1 => x111_out_17,
   I2 => M_reg_14_3,
   I3 => M_reg_14_24,
   I4 => M_reg_14_20,
   O => W_29_19_i_12_n_0
);
W_29_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x111_out_16,
   I1 => M_reg_14_19,
   I2 => M_reg_14_23,
   I3 => M_reg_14_2,
   I4 => M_reg_13_16,
   O => W_29_19_i_13_n_0
);
W_29_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_13_16,
   I1 => x111_out_16,
   I2 => M_reg_14_2,
   I3 => M_reg_14_23,
   I4 => M_reg_14_19,
   O => W_29_19_i_14_n_0
);
W_29_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x111_out_15,
   I1 => M_reg_14_18,
   I2 => M_reg_14_22,
   I3 => M_reg_14_1,
   I4 => M_reg_13_15,
   O => W_29_19_i_15_n_0
);
W_29_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_13_15,
   I1 => x111_out_15,
   I2 => M_reg_14_1,
   I3 => M_reg_14_22,
   I4 => M_reg_14_18,
   O => W_29_19_i_16_n_0
);
W_29_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x111_out_14,
   I1 => M_reg_14_17,
   I2 => M_reg_14_21,
   I3 => M_reg_14_0,
   I4 => M_reg_13_14,
   O => W_29_19_i_17_n_0
);
W_29_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x102_out_28,
   I1 => x102_out_3,
   I2 => x102_out_5,
   I3 => W_29_19_i_10_n_0,
   I4 => W_29_19_i_11_n_0,
   O => W_29_19_i_2_n_0
);
W_29_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x102_out_27,
   I1 => x102_out_2,
   I2 => x102_out_4,
   I3 => W_29_19_i_12_n_0,
   I4 => W_29_19_i_13_n_0,
   O => W_29_19_i_3_n_0
);
W_29_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x102_out_26,
   I1 => x102_out_1,
   I2 => x102_out_3,
   I3 => W_29_19_i_14_n_0,
   I4 => W_29_19_i_15_n_0,
   O => W_29_19_i_4_n_0
);
W_29_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x102_out_25,
   I1 => x102_out_0,
   I2 => x102_out_2,
   I3 => W_29_19_i_16_n_0,
   I4 => W_29_19_i_17_n_0,
   O => W_29_19_i_5_n_0
);
W_29_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_29_19_i_2_n_0,
   I1 => W_29_23_i_16_n_0,
   I2 => x102_out_29,
   I3 => x102_out_4,
   I4 => x102_out_6,
   I5 => W_29_23_i_17_n_0,
   O => W_29_19_i_6_n_0
);
W_29_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_29_19_i_3_n_0,
   I1 => W_29_19_i_10_n_0,
   I2 => x102_out_28,
   I3 => x102_out_3,
   I4 => x102_out_5,
   I5 => W_29_19_i_11_n_0,
   O => W_29_19_i_7_n_0
);
W_29_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_29_19_i_4_n_0,
   I1 => W_29_19_i_12_n_0,
   I2 => x102_out_27,
   I3 => x102_out_2,
   I4 => x102_out_4,
   I5 => W_29_19_i_13_n_0,
   O => W_29_19_i_8_n_0
);
W_29_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_29_19_i_5_n_0,
   I1 => W_29_19_i_14_n_0,
   I2 => x102_out_26,
   I3 => x102_out_1,
   I4 => x102_out_3,
   I5 => W_29_19_i_15_n_0,
   O => W_29_19_i_9_n_0
);
W_29_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_13_22,
   I1 => x111_out_22,
   I2 => M_reg_14_8,
   I3 => M_reg_14_29,
   I4 => M_reg_14_25,
   O => W_29_23_i_10_n_0
);
W_29_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x111_out_21,
   I1 => M_reg_14_24,
   I2 => M_reg_14_28,
   I3 => M_reg_14_7,
   I4 => M_reg_13_21,
   O => W_29_23_i_11_n_0
);
W_29_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_13_21,
   I1 => x111_out_21,
   I2 => M_reg_14_7,
   I3 => M_reg_14_28,
   I4 => M_reg_14_24,
   O => W_29_23_i_12_n_0
);
W_29_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x111_out_20,
   I1 => M_reg_14_23,
   I2 => M_reg_14_27,
   I3 => M_reg_14_6,
   I4 => M_reg_13_20,
   O => W_29_23_i_13_n_0
);
W_29_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_13_20,
   I1 => x111_out_20,
   I2 => M_reg_14_6,
   I3 => M_reg_14_27,
   I4 => M_reg_14_23,
   O => W_29_23_i_14_n_0
);
W_29_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x111_out_19,
   I1 => M_reg_14_22,
   I2 => M_reg_14_26,
   I3 => M_reg_14_5,
   I4 => M_reg_13_19,
   O => W_29_23_i_15_n_0
);
W_29_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_13_19,
   I1 => x111_out_19,
   I2 => M_reg_14_5,
   I3 => M_reg_14_26,
   I4 => M_reg_14_22,
   O => W_29_23_i_16_n_0
);
W_29_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x111_out_18,
   I1 => M_reg_14_21,
   I2 => M_reg_14_25,
   I3 => M_reg_14_4,
   I4 => M_reg_13_18,
   O => W_29_23_i_17_n_0
);
W_29_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x102_out_7,
   I1 => x102_out_9,
   I2 => W_29_23_i_10_n_0,
   I3 => W_29_23_i_11_n_0,
   O => W_29_23_i_2_n_0
);
W_29_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x102_out_31,
   I1 => x102_out_6,
   I2 => x102_out_8,
   I3 => W_29_23_i_12_n_0,
   I4 => W_29_23_i_13_n_0,
   O => W_29_23_i_3_n_0
);
W_29_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x102_out_30,
   I1 => x102_out_5,
   I2 => x102_out_7,
   I3 => W_29_23_i_14_n_0,
   I4 => W_29_23_i_15_n_0,
   O => W_29_23_i_4_n_0
);
W_29_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x102_out_29,
   I1 => x102_out_4,
   I2 => x102_out_6,
   I3 => W_29_23_i_16_n_0,
   I4 => W_29_23_i_17_n_0,
   O => W_29_23_i_5_n_0
);
W_29_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x102_out_8,
   I1 => x102_out_10,
   I2 => W_29_27_i_16_n_0,
   I3 => W_29_27_i_17_n_0,
   I4 => W_29_23_i_2_n_0,
   O => W_29_23_i_6_n_0
);
W_29_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x102_out_7,
   I1 => x102_out_9,
   I2 => W_29_23_i_10_n_0,
   I3 => W_29_23_i_11_n_0,
   I4 => W_29_23_i_3_n_0,
   O => W_29_23_i_7_n_0
);
W_29_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_29_23_i_4_n_0,
   I1 => W_29_23_i_12_n_0,
   I2 => x102_out_31,
   I3 => x102_out_6,
   I4 => x102_out_8,
   I5 => W_29_23_i_13_n_0,
   O => W_29_23_i_8_n_0
);
W_29_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_29_23_i_5_n_0,
   I1 => W_29_23_i_14_n_0,
   I2 => x102_out_30,
   I3 => x102_out_5,
   I4 => x102_out_7,
   I5 => W_29_23_i_15_n_0,
   O => W_29_23_i_9_n_0
);
W_29_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_13_26,
   I1 => x111_out_26,
   I2 => M_reg_14_12,
   I3 => M_reg_14_1,
   I4 => M_reg_14_29,
   O => W_29_27_i_10_n_0
);
W_29_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x111_out_25,
   I1 => M_reg_14_28,
   I2 => M_reg_14_0,
   I3 => M_reg_14_11,
   I4 => M_reg_13_25,
   O => W_29_27_i_11_n_0
);
W_29_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_13_25,
   I1 => x111_out_25,
   I2 => M_reg_14_11,
   I3 => M_reg_14_0,
   I4 => M_reg_14_28,
   O => W_29_27_i_12_n_0
);
W_29_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x111_out_24,
   I1 => M_reg_14_27,
   I2 => M_reg_14_31,
   I3 => M_reg_14_10,
   I4 => M_reg_13_24,
   O => W_29_27_i_13_n_0
);
W_29_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_13_24,
   I1 => x111_out_24,
   I2 => M_reg_14_10,
   I3 => M_reg_14_31,
   I4 => M_reg_14_27,
   O => W_29_27_i_14_n_0
);
W_29_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x111_out_23,
   I1 => M_reg_14_26,
   I2 => M_reg_14_30,
   I3 => M_reg_14_9,
   I4 => M_reg_13_23,
   O => W_29_27_i_15_n_0
);
W_29_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_13_23,
   I1 => x111_out_23,
   I2 => M_reg_14_9,
   I3 => M_reg_14_30,
   I4 => M_reg_14_26,
   O => W_29_27_i_16_n_0
);
W_29_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x111_out_22,
   I1 => M_reg_14_25,
   I2 => M_reg_14_29,
   I3 => M_reg_14_8,
   I4 => M_reg_13_22,
   O => W_29_27_i_17_n_0
);
W_29_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x102_out_11,
   I1 => x102_out_13,
   I2 => W_29_27_i_10_n_0,
   I3 => W_29_27_i_11_n_0,
   O => W_29_27_i_2_n_0
);
W_29_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x102_out_10,
   I1 => x102_out_12,
   I2 => W_29_27_i_12_n_0,
   I3 => W_29_27_i_13_n_0,
   O => W_29_27_i_3_n_0
);
W_29_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x102_out_9,
   I1 => x102_out_11,
   I2 => W_29_27_i_14_n_0,
   I3 => W_29_27_i_15_n_0,
   O => W_29_27_i_4_n_0
);
W_29_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x102_out_8,
   I1 => x102_out_10,
   I2 => W_29_27_i_16_n_0,
   I3 => W_29_27_i_17_n_0,
   O => W_29_27_i_5_n_0
);
W_29_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x102_out_12,
   I1 => x102_out_14,
   I2 => W_29_31_i_13_n_0,
   I3 => W_29_31_i_14_n_0,
   I4 => W_29_27_i_2_n_0,
   O => W_29_27_i_6_n_0
);
W_29_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x102_out_11,
   I1 => x102_out_13,
   I2 => W_29_27_i_10_n_0,
   I3 => W_29_27_i_11_n_0,
   I4 => W_29_27_i_3_n_0,
   O => W_29_27_i_7_n_0
);
W_29_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x102_out_10,
   I1 => x102_out_12,
   I2 => W_29_27_i_12_n_0,
   I3 => W_29_27_i_13_n_0,
   I4 => W_29_27_i_4_n_0,
   O => W_29_27_i_8_n_0
);
W_29_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x102_out_9,
   I1 => x102_out_11,
   I2 => W_29_27_i_14_n_0,
   I3 => W_29_27_i_15_n_0,
   I4 => W_29_27_i_5_n_0,
   O => W_29_27_i_9_n_0
);
W_29_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x111_out_28,
   I1 => M_reg_14_31,
   I2 => M_reg_14_3,
   I3 => M_reg_14_14,
   I4 => M_reg_13_28,
   O => W_29_31_i_10_n_0
);
W_29_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_13_28,
   I1 => x111_out_28,
   I2 => M_reg_14_14,
   I3 => M_reg_14_3,
   I4 => M_reg_14_31,
   O => W_29_31_i_11_n_0
);
W_29_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x111_out_27,
   I1 => M_reg_14_30,
   I2 => M_reg_14_2,
   I3 => M_reg_14_13,
   I4 => M_reg_13_27,
   O => W_29_31_i_12_n_0
);
W_29_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_13_27,
   I1 => x111_out_27,
   I2 => M_reg_14_13,
   I3 => M_reg_14_2,
   I4 => M_reg_14_30,
   O => W_29_31_i_13_n_0
);
W_29_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x111_out_26,
   I1 => M_reg_14_29,
   I2 => M_reg_14_1,
   I3 => M_reg_14_12,
   I4 => M_reg_13_26,
   O => W_29_31_i_14_n_0
);
W_29_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x111_out_29,
   I1 => M_reg_14_4,
   I2 => M_reg_14_15,
   I3 => M_reg_13_29,
   O => W_29_31_i_15_n_0
);
W_29_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x102_out_17,
   I1 => x102_out_15,
   O => SIGMA_LCASE_1283_out_0_30
);
W_29_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => M_reg_14_6,
   I1 => M_reg_14_17,
   I2 => x111_out_31,
   I3 => M_reg_13_31,
   I4 => x102_out_16,
   I5 => x102_out_18,
   O => W_29_31_i_17_n_0
);
W_29_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => M_reg_14_16,
   I1 => M_reg_14_5,
   O => SIGMA_LCASE_0279_out_30
);
W_29_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => M_reg_13_30,
   I1 => x111_out_30,
   I2 => M_reg_14_16,
   I3 => M_reg_14_5,
   O => W_29_31_i_19_n_0
);
W_29_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x102_out_14,
   I1 => x102_out_16,
   I2 => W_29_31_i_9_n_0,
   I3 => W_29_31_i_10_n_0,
   O => W_29_31_i_2_n_0
);
W_29_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x102_out_13,
   I1 => x102_out_15,
   I2 => W_29_31_i_11_n_0,
   I3 => W_29_31_i_12_n_0,
   O => W_29_31_i_3_n_0
);
W_29_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x102_out_12,
   I1 => x102_out_14,
   I2 => W_29_31_i_13_n_0,
   I3 => W_29_31_i_14_n_0,
   O => W_29_31_i_4_n_0
);
W_29_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_29_31_i_15_n_0,
   I1 => SIGMA_LCASE_1283_out_0_30,
   I2 => W_29_31_i_17_n_0,
   I3 => x111_out_30,
   I4 => SIGMA_LCASE_0279_out_30,
   I5 => M_reg_13_30,
   O => W_29_31_i_5_n_0
);
W_29_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_29_31_i_2_n_0,
   I1 => W_29_31_i_19_n_0,
   I2 => x102_out_15,
   I3 => x102_out_17,
   I4 => W_29_31_i_15_n_0,
   O => W_29_31_i_6_n_0
);
W_29_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x102_out_14,
   I1 => x102_out_16,
   I2 => W_29_31_i_9_n_0,
   I3 => W_29_31_i_10_n_0,
   I4 => W_29_31_i_3_n_0,
   O => W_29_31_i_7_n_0
);
W_29_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x102_out_13,
   I1 => x102_out_15,
   I2 => W_29_31_i_11_n_0,
   I3 => W_29_31_i_12_n_0,
   I4 => W_29_31_i_4_n_0,
   O => W_29_31_i_8_n_0
);
W_29_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => M_reg_13_29,
   I1 => x111_out_29,
   I2 => M_reg_14_15,
   I3 => M_reg_14_4,
   O => W_29_31_i_9_n_0
);
W_29_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_13_2,
   I1 => x111_out_2,
   I2 => M_reg_14_20,
   I3 => M_reg_14_9,
   I4 => M_reg_14_5,
   O => W_29_3_i_10_n_0
);
W_29_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x111_out_1,
   I1 => M_reg_14_4,
   I2 => M_reg_14_8,
   I3 => M_reg_14_19,
   I4 => M_reg_13_1,
   O => W_29_3_i_11_n_0
);
W_29_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => M_reg_14_19,
   I1 => M_reg_14_8,
   I2 => M_reg_14_4,
   O => SIGMA_LCASE_0279_out_1
);
W_29_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x102_out_21,
   I1 => x102_out_19,
   I2 => x102_out_12,
   O => SIGMA_LCASE_1283_out_0_2
);
W_29_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x102_out_20,
   I1 => x102_out_18,
   I2 => x102_out_11,
   O => SIGMA_LCASE_1283_out_1
);
W_29_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x102_out_12,
   I1 => x102_out_19,
   I2 => x102_out_21,
   I3 => W_29_3_i_10_n_0,
   I4 => W_29_3_i_11_n_0,
   O => W_29_3_i_2_n_0
);
W_29_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_29_3_i_11_n_0,
   I1 => x102_out_21,
   I2 => x102_out_19,
   I3 => x102_out_12,
   I4 => W_29_3_i_10_n_0,
   O => W_29_3_i_3_n_0
);
W_29_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_0279_out_1,
   I1 => x111_out_1,
   I2 => M_reg_13_1,
   I3 => x102_out_11,
   I4 => x102_out_18,
   I5 => x102_out_20,
   O => W_29_3_i_4_n_0
);
W_29_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_13_0,
   I1 => x111_out_0,
   I2 => M_reg_14_18,
   I3 => M_reg_14_7,
   I4 => M_reg_14_3,
   O => W_29_3_i_5_n_0
);
W_29_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_29_3_i_2_n_0,
   I1 => W_29_7_i_16_n_0,
   I2 => x102_out_13,
   I3 => x102_out_20,
   I4 => x102_out_22,
   I5 => W_29_7_i_17_n_0,
   O => W_29_3_i_6_n_0
);
W_29_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_29_3_i_10_n_0,
   I1 => SIGMA_LCASE_1283_out_0_2,
   I2 => M_reg_13_1,
   I3 => x111_out_1,
   I4 => SIGMA_LCASE_0279_out_1,
   I5 => SIGMA_LCASE_1283_out_1,
   O => W_29_3_i_7_n_0
);
W_29_3_i_8 : LUT6
  generic map(
   INIT => X"566565566aa6a66a"
  )
 port map (
   I0 => W_29_3_i_4_n_0,
   I1 => M_reg_13_0,
   I2 => M_reg_14_18,
   I3 => M_reg_14_7,
   I4 => M_reg_14_3,
   I5 => x111_out_0,
   O => W_29_3_i_8_n_0
);
W_29_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_29_3_i_5_n_0,
   I1 => x102_out_10,
   I2 => x102_out_17,
   I3 => x102_out_19,
   O => W_29_3_i_9_n_0
);
W_29_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_13_6,
   I1 => x111_out_6,
   I2 => M_reg_14_24,
   I3 => M_reg_14_13,
   I4 => M_reg_14_9,
   O => W_29_7_i_10_n_0
);
W_29_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x111_out_5,
   I1 => M_reg_14_8,
   I2 => M_reg_14_12,
   I3 => M_reg_14_23,
   I4 => M_reg_13_5,
   O => W_29_7_i_11_n_0
);
W_29_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_13_5,
   I1 => x111_out_5,
   I2 => M_reg_14_23,
   I3 => M_reg_14_12,
   I4 => M_reg_14_8,
   O => W_29_7_i_12_n_0
);
W_29_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x111_out_4,
   I1 => M_reg_14_7,
   I2 => M_reg_14_11,
   I3 => M_reg_14_22,
   I4 => M_reg_13_4,
   O => W_29_7_i_13_n_0
);
W_29_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_13_4,
   I1 => x111_out_4,
   I2 => M_reg_14_22,
   I3 => M_reg_14_11,
   I4 => M_reg_14_7,
   O => W_29_7_i_14_n_0
);
W_29_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x111_out_3,
   I1 => M_reg_14_6,
   I2 => M_reg_14_10,
   I3 => M_reg_14_21,
   I4 => M_reg_13_3,
   O => W_29_7_i_15_n_0
);
W_29_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_13_3,
   I1 => x111_out_3,
   I2 => M_reg_14_21,
   I3 => M_reg_14_10,
   I4 => M_reg_14_6,
   O => W_29_7_i_16_n_0
);
W_29_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x111_out_2,
   I1 => M_reg_14_5,
   I2 => M_reg_14_9,
   I3 => M_reg_14_20,
   I4 => M_reg_13_2,
   O => W_29_7_i_17_n_0
);
W_29_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x102_out_16,
   I1 => x102_out_23,
   I2 => x102_out_25,
   I3 => W_29_7_i_10_n_0,
   I4 => W_29_7_i_11_n_0,
   O => W_29_7_i_2_n_0
);
W_29_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x102_out_15,
   I1 => x102_out_22,
   I2 => x102_out_24,
   I3 => W_29_7_i_12_n_0,
   I4 => W_29_7_i_13_n_0,
   O => W_29_7_i_3_n_0
);
W_29_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x102_out_14,
   I1 => x102_out_21,
   I2 => x102_out_23,
   I3 => W_29_7_i_14_n_0,
   I4 => W_29_7_i_15_n_0,
   O => W_29_7_i_4_n_0
);
W_29_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x102_out_13,
   I1 => x102_out_20,
   I2 => x102_out_22,
   I3 => W_29_7_i_16_n_0,
   I4 => W_29_7_i_17_n_0,
   O => W_29_7_i_5_n_0
);
W_29_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_29_7_i_2_n_0,
   I1 => W_29_11_i_16_n_0,
   I2 => x102_out_17,
   I3 => x102_out_24,
   I4 => x102_out_26,
   I5 => W_29_11_i_17_n_0,
   O => W_29_7_i_6_n_0
);
W_29_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_29_7_i_3_n_0,
   I1 => W_29_7_i_10_n_0,
   I2 => x102_out_16,
   I3 => x102_out_23,
   I4 => x102_out_25,
   I5 => W_29_7_i_11_n_0,
   O => W_29_7_i_7_n_0
);
W_29_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_29_7_i_4_n_0,
   I1 => W_29_7_i_12_n_0,
   I2 => x102_out_15,
   I3 => x102_out_22,
   I4 => x102_out_24,
   I5 => W_29_7_i_13_n_0,
   O => W_29_7_i_8_n_0
);
W_29_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_29_7_i_5_n_0,
   I1 => W_29_7_i_14_n_0,
   I2 => x102_out_14,
   I3 => x102_out_21,
   I4 => x102_out_23,
   I5 => W_29_7_i_15_n_0,
   O => W_29_7_i_9_n_0
);
W_30_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_14_10,
   I1 => x110_out_10,
   I2 => M_reg_15_28,
   I3 => M_reg_15_17,
   I4 => M_reg_15_13,
   O => W_30_11_i_10_n_0
);
W_30_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x110_out_9,
   I1 => M_reg_15_12,
   I2 => M_reg_15_16,
   I3 => M_reg_15_27,
   I4 => M_reg_14_9,
   O => W_30_11_i_11_n_0
);
W_30_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_14_9,
   I1 => x110_out_9,
   I2 => M_reg_15_27,
   I3 => M_reg_15_16,
   I4 => M_reg_15_12,
   O => W_30_11_i_12_n_0
);
W_30_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x110_out_8,
   I1 => M_reg_15_11,
   I2 => M_reg_15_15,
   I3 => M_reg_15_26,
   I4 => M_reg_14_8,
   O => W_30_11_i_13_n_0
);
W_30_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_14_8,
   I1 => x110_out_8,
   I2 => M_reg_15_26,
   I3 => M_reg_15_15,
   I4 => M_reg_15_11,
   O => W_30_11_i_14_n_0
);
W_30_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x110_out_7,
   I1 => M_reg_15_10,
   I2 => M_reg_15_14,
   I3 => M_reg_15_25,
   I4 => M_reg_14_7,
   O => W_30_11_i_15_n_0
);
W_30_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_14_7,
   I1 => x110_out_7,
   I2 => M_reg_15_25,
   I3 => M_reg_15_14,
   I4 => M_reg_15_10,
   O => W_30_11_i_16_n_0
);
W_30_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x110_out_6,
   I1 => M_reg_15_9,
   I2 => M_reg_15_13,
   I3 => M_reg_15_24,
   I4 => M_reg_14_6,
   O => W_30_11_i_17_n_0
);
W_30_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x100_out_20,
   I1 => x100_out_27,
   I2 => x100_out_29,
   I3 => W_30_11_i_10_n_0,
   I4 => W_30_11_i_11_n_0,
   O => W_30_11_i_2_n_0
);
W_30_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x100_out_19,
   I1 => x100_out_26,
   I2 => x100_out_28,
   I3 => W_30_11_i_12_n_0,
   I4 => W_30_11_i_13_n_0,
   O => W_30_11_i_3_n_0
);
W_30_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x100_out_18,
   I1 => x100_out_25,
   I2 => x100_out_27,
   I3 => W_30_11_i_14_n_0,
   I4 => W_30_11_i_15_n_0,
   O => W_30_11_i_4_n_0
);
W_30_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x100_out_17,
   I1 => x100_out_24,
   I2 => x100_out_26,
   I3 => W_30_11_i_16_n_0,
   I4 => W_30_11_i_17_n_0,
   O => W_30_11_i_5_n_0
);
W_30_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_30_11_i_2_n_0,
   I1 => W_30_15_i_16_n_0,
   I2 => x100_out_21,
   I3 => x100_out_28,
   I4 => x100_out_30,
   I5 => W_30_15_i_17_n_0,
   O => W_30_11_i_6_n_0
);
W_30_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_30_11_i_3_n_0,
   I1 => W_30_11_i_10_n_0,
   I2 => x100_out_20,
   I3 => x100_out_27,
   I4 => x100_out_29,
   I5 => W_30_11_i_11_n_0,
   O => W_30_11_i_7_n_0
);
W_30_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_30_11_i_4_n_0,
   I1 => W_30_11_i_12_n_0,
   I2 => x100_out_19,
   I3 => x100_out_26,
   I4 => x100_out_28,
   I5 => W_30_11_i_13_n_0,
   O => W_30_11_i_8_n_0
);
W_30_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_30_11_i_5_n_0,
   I1 => W_30_11_i_14_n_0,
   I2 => x100_out_18,
   I3 => x100_out_25,
   I4 => x100_out_27,
   I5 => W_30_11_i_15_n_0,
   O => W_30_11_i_9_n_0
);
W_30_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_14_14,
   I1 => x110_out_14,
   I2 => M_reg_15_0,
   I3 => M_reg_15_21,
   I4 => M_reg_15_17,
   O => W_30_15_i_10_n_0
);
W_30_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x110_out_13,
   I1 => M_reg_15_16,
   I2 => M_reg_15_20,
   I3 => M_reg_15_31,
   I4 => M_reg_14_13,
   O => W_30_15_i_11_n_0
);
W_30_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_14_13,
   I1 => x110_out_13,
   I2 => M_reg_15_31,
   I3 => M_reg_15_20,
   I4 => M_reg_15_16,
   O => W_30_15_i_12_n_0
);
W_30_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x110_out_12,
   I1 => M_reg_15_15,
   I2 => M_reg_15_19,
   I3 => M_reg_15_30,
   I4 => M_reg_14_12,
   O => W_30_15_i_13_n_0
);
W_30_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_14_12,
   I1 => x110_out_12,
   I2 => M_reg_15_30,
   I3 => M_reg_15_19,
   I4 => M_reg_15_15,
   O => W_30_15_i_14_n_0
);
W_30_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x110_out_11,
   I1 => M_reg_15_14,
   I2 => M_reg_15_18,
   I3 => M_reg_15_29,
   I4 => M_reg_14_11,
   O => W_30_15_i_15_n_0
);
W_30_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_14_11,
   I1 => x110_out_11,
   I2 => M_reg_15_29,
   I3 => M_reg_15_18,
   I4 => M_reg_15_14,
   O => W_30_15_i_16_n_0
);
W_30_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x110_out_10,
   I1 => M_reg_15_13,
   I2 => M_reg_15_17,
   I3 => M_reg_15_28,
   I4 => M_reg_14_10,
   O => W_30_15_i_17_n_0
);
W_30_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x100_out_24,
   I1 => x100_out_31,
   I2 => x100_out_1,
   I3 => W_30_15_i_10_n_0,
   I4 => W_30_15_i_11_n_0,
   O => W_30_15_i_2_n_0
);
W_30_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x100_out_23,
   I1 => x100_out_30,
   I2 => x100_out_0,
   I3 => W_30_15_i_12_n_0,
   I4 => W_30_15_i_13_n_0,
   O => W_30_15_i_3_n_0
);
W_30_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x100_out_22,
   I1 => x100_out_29,
   I2 => x100_out_31,
   I3 => W_30_15_i_14_n_0,
   I4 => W_30_15_i_15_n_0,
   O => W_30_15_i_4_n_0
);
W_30_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x100_out_21,
   I1 => x100_out_28,
   I2 => x100_out_30,
   I3 => W_30_15_i_16_n_0,
   I4 => W_30_15_i_17_n_0,
   O => W_30_15_i_5_n_0
);
W_30_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_30_15_i_2_n_0,
   I1 => W_30_19_i_16_n_0,
   I2 => x100_out_25,
   I3 => x100_out_0,
   I4 => x100_out_2,
   I5 => W_30_19_i_17_n_0,
   O => W_30_15_i_6_n_0
);
W_30_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_30_15_i_3_n_0,
   I1 => W_30_15_i_10_n_0,
   I2 => x100_out_24,
   I3 => x100_out_31,
   I4 => x100_out_1,
   I5 => W_30_15_i_11_n_0,
   O => W_30_15_i_7_n_0
);
W_30_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_30_15_i_4_n_0,
   I1 => W_30_15_i_12_n_0,
   I2 => x100_out_23,
   I3 => x100_out_30,
   I4 => x100_out_0,
   I5 => W_30_15_i_13_n_0,
   O => W_30_15_i_8_n_0
);
W_30_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_30_15_i_5_n_0,
   I1 => W_30_15_i_14_n_0,
   I2 => x100_out_22,
   I3 => x100_out_29,
   I4 => x100_out_31,
   I5 => W_30_15_i_15_n_0,
   O => W_30_15_i_9_n_0
);
W_30_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_14_18,
   I1 => x110_out_18,
   I2 => M_reg_15_4,
   I3 => M_reg_15_25,
   I4 => M_reg_15_21,
   O => W_30_19_i_10_n_0
);
W_30_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x110_out_17,
   I1 => M_reg_15_20,
   I2 => M_reg_15_24,
   I3 => M_reg_15_3,
   I4 => M_reg_14_17,
   O => W_30_19_i_11_n_0
);
W_30_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_14_17,
   I1 => x110_out_17,
   I2 => M_reg_15_3,
   I3 => M_reg_15_24,
   I4 => M_reg_15_20,
   O => W_30_19_i_12_n_0
);
W_30_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x110_out_16,
   I1 => M_reg_15_19,
   I2 => M_reg_15_23,
   I3 => M_reg_15_2,
   I4 => M_reg_14_16,
   O => W_30_19_i_13_n_0
);
W_30_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_14_16,
   I1 => x110_out_16,
   I2 => M_reg_15_2,
   I3 => M_reg_15_23,
   I4 => M_reg_15_19,
   O => W_30_19_i_14_n_0
);
W_30_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x110_out_15,
   I1 => M_reg_15_18,
   I2 => M_reg_15_22,
   I3 => M_reg_15_1,
   I4 => M_reg_14_15,
   O => W_30_19_i_15_n_0
);
W_30_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_14_15,
   I1 => x110_out_15,
   I2 => M_reg_15_1,
   I3 => M_reg_15_22,
   I4 => M_reg_15_18,
   O => W_30_19_i_16_n_0
);
W_30_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x110_out_14,
   I1 => M_reg_15_17,
   I2 => M_reg_15_21,
   I3 => M_reg_15_0,
   I4 => M_reg_14_14,
   O => W_30_19_i_17_n_0
);
W_30_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x100_out_28,
   I1 => x100_out_3,
   I2 => x100_out_5,
   I3 => W_30_19_i_10_n_0,
   I4 => W_30_19_i_11_n_0,
   O => W_30_19_i_2_n_0
);
W_30_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x100_out_27,
   I1 => x100_out_2,
   I2 => x100_out_4,
   I3 => W_30_19_i_12_n_0,
   I4 => W_30_19_i_13_n_0,
   O => W_30_19_i_3_n_0
);
W_30_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x100_out_26,
   I1 => x100_out_1,
   I2 => x100_out_3,
   I3 => W_30_19_i_14_n_0,
   I4 => W_30_19_i_15_n_0,
   O => W_30_19_i_4_n_0
);
W_30_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x100_out_25,
   I1 => x100_out_0,
   I2 => x100_out_2,
   I3 => W_30_19_i_16_n_0,
   I4 => W_30_19_i_17_n_0,
   O => W_30_19_i_5_n_0
);
W_30_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_30_19_i_2_n_0,
   I1 => W_30_23_i_16_n_0,
   I2 => x100_out_29,
   I3 => x100_out_4,
   I4 => x100_out_6,
   I5 => W_30_23_i_17_n_0,
   O => W_30_19_i_6_n_0
);
W_30_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_30_19_i_3_n_0,
   I1 => W_30_19_i_10_n_0,
   I2 => x100_out_28,
   I3 => x100_out_3,
   I4 => x100_out_5,
   I5 => W_30_19_i_11_n_0,
   O => W_30_19_i_7_n_0
);
W_30_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_30_19_i_4_n_0,
   I1 => W_30_19_i_12_n_0,
   I2 => x100_out_27,
   I3 => x100_out_2,
   I4 => x100_out_4,
   I5 => W_30_19_i_13_n_0,
   O => W_30_19_i_8_n_0
);
W_30_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_30_19_i_5_n_0,
   I1 => W_30_19_i_14_n_0,
   I2 => x100_out_26,
   I3 => x100_out_1,
   I4 => x100_out_3,
   I5 => W_30_19_i_15_n_0,
   O => W_30_19_i_9_n_0
);
W_30_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_14_22,
   I1 => x110_out_22,
   I2 => M_reg_15_8,
   I3 => M_reg_15_29,
   I4 => M_reg_15_25,
   O => W_30_23_i_10_n_0
);
W_30_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x110_out_21,
   I1 => M_reg_15_24,
   I2 => M_reg_15_28,
   I3 => M_reg_15_7,
   I4 => M_reg_14_21,
   O => W_30_23_i_11_n_0
);
W_30_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_14_21,
   I1 => x110_out_21,
   I2 => M_reg_15_7,
   I3 => M_reg_15_28,
   I4 => M_reg_15_24,
   O => W_30_23_i_12_n_0
);
W_30_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x110_out_20,
   I1 => M_reg_15_23,
   I2 => M_reg_15_27,
   I3 => M_reg_15_6,
   I4 => M_reg_14_20,
   O => W_30_23_i_13_n_0
);
W_30_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_14_20,
   I1 => x110_out_20,
   I2 => M_reg_15_6,
   I3 => M_reg_15_27,
   I4 => M_reg_15_23,
   O => W_30_23_i_14_n_0
);
W_30_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x110_out_19,
   I1 => M_reg_15_22,
   I2 => M_reg_15_26,
   I3 => M_reg_15_5,
   I4 => M_reg_14_19,
   O => W_30_23_i_15_n_0
);
W_30_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_14_19,
   I1 => x110_out_19,
   I2 => M_reg_15_5,
   I3 => M_reg_15_26,
   I4 => M_reg_15_22,
   O => W_30_23_i_16_n_0
);
W_30_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x110_out_18,
   I1 => M_reg_15_21,
   I2 => M_reg_15_25,
   I3 => M_reg_15_4,
   I4 => M_reg_14_18,
   O => W_30_23_i_17_n_0
);
W_30_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x100_out_7,
   I1 => x100_out_9,
   I2 => W_30_23_i_10_n_0,
   I3 => W_30_23_i_11_n_0,
   O => W_30_23_i_2_n_0
);
W_30_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x100_out_31,
   I1 => x100_out_6,
   I2 => x100_out_8,
   I3 => W_30_23_i_12_n_0,
   I4 => W_30_23_i_13_n_0,
   O => W_30_23_i_3_n_0
);
W_30_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x100_out_30,
   I1 => x100_out_5,
   I2 => x100_out_7,
   I3 => W_30_23_i_14_n_0,
   I4 => W_30_23_i_15_n_0,
   O => W_30_23_i_4_n_0
);
W_30_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x100_out_29,
   I1 => x100_out_4,
   I2 => x100_out_6,
   I3 => W_30_23_i_16_n_0,
   I4 => W_30_23_i_17_n_0,
   O => W_30_23_i_5_n_0
);
W_30_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x100_out_8,
   I1 => x100_out_10,
   I2 => W_30_27_i_16_n_0,
   I3 => W_30_27_i_17_n_0,
   I4 => W_30_23_i_2_n_0,
   O => W_30_23_i_6_n_0
);
W_30_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x100_out_7,
   I1 => x100_out_9,
   I2 => W_30_23_i_10_n_0,
   I3 => W_30_23_i_11_n_0,
   I4 => W_30_23_i_3_n_0,
   O => W_30_23_i_7_n_0
);
W_30_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_30_23_i_4_n_0,
   I1 => W_30_23_i_12_n_0,
   I2 => x100_out_31,
   I3 => x100_out_6,
   I4 => x100_out_8,
   I5 => W_30_23_i_13_n_0,
   O => W_30_23_i_8_n_0
);
W_30_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_30_23_i_5_n_0,
   I1 => W_30_23_i_14_n_0,
   I2 => x100_out_30,
   I3 => x100_out_5,
   I4 => x100_out_7,
   I5 => W_30_23_i_15_n_0,
   O => W_30_23_i_9_n_0
);
W_30_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_14_26,
   I1 => x110_out_26,
   I2 => M_reg_15_12,
   I3 => M_reg_15_1,
   I4 => M_reg_15_29,
   O => W_30_27_i_10_n_0
);
W_30_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x110_out_25,
   I1 => M_reg_15_28,
   I2 => M_reg_15_0,
   I3 => M_reg_15_11,
   I4 => M_reg_14_25,
   O => W_30_27_i_11_n_0
);
W_30_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_14_25,
   I1 => x110_out_25,
   I2 => M_reg_15_11,
   I3 => M_reg_15_0,
   I4 => M_reg_15_28,
   O => W_30_27_i_12_n_0
);
W_30_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x110_out_24,
   I1 => M_reg_15_27,
   I2 => M_reg_15_31,
   I3 => M_reg_15_10,
   I4 => M_reg_14_24,
   O => W_30_27_i_13_n_0
);
W_30_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_14_24,
   I1 => x110_out_24,
   I2 => M_reg_15_10,
   I3 => M_reg_15_31,
   I4 => M_reg_15_27,
   O => W_30_27_i_14_n_0
);
W_30_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x110_out_23,
   I1 => M_reg_15_26,
   I2 => M_reg_15_30,
   I3 => M_reg_15_9,
   I4 => M_reg_14_23,
   O => W_30_27_i_15_n_0
);
W_30_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_14_23,
   I1 => x110_out_23,
   I2 => M_reg_15_9,
   I3 => M_reg_15_30,
   I4 => M_reg_15_26,
   O => W_30_27_i_16_n_0
);
W_30_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x110_out_22,
   I1 => M_reg_15_25,
   I2 => M_reg_15_29,
   I3 => M_reg_15_8,
   I4 => M_reg_14_22,
   O => W_30_27_i_17_n_0
);
W_30_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x100_out_11,
   I1 => x100_out_13,
   I2 => W_30_27_i_10_n_0,
   I3 => W_30_27_i_11_n_0,
   O => W_30_27_i_2_n_0
);
W_30_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x100_out_10,
   I1 => x100_out_12,
   I2 => W_30_27_i_12_n_0,
   I3 => W_30_27_i_13_n_0,
   O => W_30_27_i_3_n_0
);
W_30_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x100_out_9,
   I1 => x100_out_11,
   I2 => W_30_27_i_14_n_0,
   I3 => W_30_27_i_15_n_0,
   O => W_30_27_i_4_n_0
);
W_30_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x100_out_8,
   I1 => x100_out_10,
   I2 => W_30_27_i_16_n_0,
   I3 => W_30_27_i_17_n_0,
   O => W_30_27_i_5_n_0
);
W_30_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x100_out_12,
   I1 => x100_out_14,
   I2 => W_30_31_i_13_n_0,
   I3 => W_30_31_i_14_n_0,
   I4 => W_30_27_i_2_n_0,
   O => W_30_27_i_6_n_0
);
W_30_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x100_out_11,
   I1 => x100_out_13,
   I2 => W_30_27_i_10_n_0,
   I3 => W_30_27_i_11_n_0,
   I4 => W_30_27_i_3_n_0,
   O => W_30_27_i_7_n_0
);
W_30_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x100_out_10,
   I1 => x100_out_12,
   I2 => W_30_27_i_12_n_0,
   I3 => W_30_27_i_13_n_0,
   I4 => W_30_27_i_4_n_0,
   O => W_30_27_i_8_n_0
);
W_30_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x100_out_9,
   I1 => x100_out_11,
   I2 => W_30_27_i_14_n_0,
   I3 => W_30_27_i_15_n_0,
   I4 => W_30_27_i_5_n_0,
   O => W_30_27_i_9_n_0
);
W_30_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x110_out_28,
   I1 => M_reg_15_31,
   I2 => M_reg_15_3,
   I3 => M_reg_15_14,
   I4 => M_reg_14_28,
   O => W_30_31_i_10_n_0
);
W_30_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_14_28,
   I1 => x110_out_28,
   I2 => M_reg_15_14,
   I3 => M_reg_15_3,
   I4 => M_reg_15_31,
   O => W_30_31_i_11_n_0
);
W_30_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x110_out_27,
   I1 => M_reg_15_30,
   I2 => M_reg_15_2,
   I3 => M_reg_15_13,
   I4 => M_reg_14_27,
   O => W_30_31_i_12_n_0
);
W_30_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_14_27,
   I1 => x110_out_27,
   I2 => M_reg_15_13,
   I3 => M_reg_15_2,
   I4 => M_reg_15_30,
   O => W_30_31_i_13_n_0
);
W_30_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x110_out_26,
   I1 => M_reg_15_29,
   I2 => M_reg_15_1,
   I3 => M_reg_15_12,
   I4 => M_reg_14_26,
   O => W_30_31_i_14_n_0
);
W_30_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x110_out_29,
   I1 => M_reg_15_4,
   I2 => M_reg_15_15,
   I3 => M_reg_14_29,
   O => W_30_31_i_15_n_0
);
W_30_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x100_out_17,
   I1 => x100_out_15,
   O => SIGMA_LCASE_1275_out_0_30
);
W_30_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => M_reg_15_6,
   I1 => M_reg_15_17,
   I2 => x110_out_31,
   I3 => M_reg_14_31,
   I4 => x100_out_16,
   I5 => x100_out_18,
   O => W_30_31_i_17_n_0
);
W_30_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => M_reg_15_16,
   I1 => M_reg_15_5,
   O => SIGMA_LCASE_0271_out_30
);
W_30_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => M_reg_14_30,
   I1 => x110_out_30,
   I2 => M_reg_15_16,
   I3 => M_reg_15_5,
   O => W_30_31_i_19_n_0
);
W_30_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x100_out_14,
   I1 => x100_out_16,
   I2 => W_30_31_i_9_n_0,
   I3 => W_30_31_i_10_n_0,
   O => W_30_31_i_2_n_0
);
W_30_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x100_out_13,
   I1 => x100_out_15,
   I2 => W_30_31_i_11_n_0,
   I3 => W_30_31_i_12_n_0,
   O => W_30_31_i_3_n_0
);
W_30_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x100_out_12,
   I1 => x100_out_14,
   I2 => W_30_31_i_13_n_0,
   I3 => W_30_31_i_14_n_0,
   O => W_30_31_i_4_n_0
);
W_30_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_30_31_i_15_n_0,
   I1 => SIGMA_LCASE_1275_out_0_30,
   I2 => W_30_31_i_17_n_0,
   I3 => x110_out_30,
   I4 => SIGMA_LCASE_0271_out_30,
   I5 => M_reg_14_30,
   O => W_30_31_i_5_n_0
);
W_30_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_30_31_i_2_n_0,
   I1 => W_30_31_i_19_n_0,
   I2 => x100_out_15,
   I3 => x100_out_17,
   I4 => W_30_31_i_15_n_0,
   O => W_30_31_i_6_n_0
);
W_30_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x100_out_14,
   I1 => x100_out_16,
   I2 => W_30_31_i_9_n_0,
   I3 => W_30_31_i_10_n_0,
   I4 => W_30_31_i_3_n_0,
   O => W_30_31_i_7_n_0
);
W_30_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x100_out_13,
   I1 => x100_out_15,
   I2 => W_30_31_i_11_n_0,
   I3 => W_30_31_i_12_n_0,
   I4 => W_30_31_i_4_n_0,
   O => W_30_31_i_8_n_0
);
W_30_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => M_reg_14_29,
   I1 => x110_out_29,
   I2 => M_reg_15_15,
   I3 => M_reg_15_4,
   O => W_30_31_i_9_n_0
);
W_30_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_14_2,
   I1 => x110_out_2,
   I2 => M_reg_15_20,
   I3 => M_reg_15_9,
   I4 => M_reg_15_5,
   O => W_30_3_i_10_n_0
);
W_30_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x110_out_1,
   I1 => M_reg_15_4,
   I2 => M_reg_15_8,
   I3 => M_reg_15_19,
   I4 => M_reg_14_1,
   O => W_30_3_i_11_n_0
);
W_30_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => M_reg_15_19,
   I1 => M_reg_15_8,
   I2 => M_reg_15_4,
   O => SIGMA_LCASE_0271_out_1
);
W_30_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x100_out_21,
   I1 => x100_out_19,
   I2 => x100_out_12,
   O => SIGMA_LCASE_1275_out_0_2
);
W_30_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x100_out_20,
   I1 => x100_out_18,
   I2 => x100_out_11,
   O => SIGMA_LCASE_1275_out_1
);
W_30_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x100_out_12,
   I1 => x100_out_19,
   I2 => x100_out_21,
   I3 => W_30_3_i_10_n_0,
   I4 => W_30_3_i_11_n_0,
   O => W_30_3_i_2_n_0
);
W_30_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_30_3_i_11_n_0,
   I1 => x100_out_21,
   I2 => x100_out_19,
   I3 => x100_out_12,
   I4 => W_30_3_i_10_n_0,
   O => W_30_3_i_3_n_0
);
W_30_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_0271_out_1,
   I1 => x110_out_1,
   I2 => M_reg_14_1,
   I3 => x100_out_11,
   I4 => x100_out_18,
   I5 => x100_out_20,
   O => W_30_3_i_4_n_0
);
W_30_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_14_0,
   I1 => x110_out_0,
   I2 => M_reg_15_18,
   I3 => M_reg_15_7,
   I4 => M_reg_15_3,
   O => W_30_3_i_5_n_0
);
W_30_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_30_3_i_2_n_0,
   I1 => W_30_7_i_16_n_0,
   I2 => x100_out_13,
   I3 => x100_out_20,
   I4 => x100_out_22,
   I5 => W_30_7_i_17_n_0,
   O => W_30_3_i_6_n_0
);
W_30_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_30_3_i_10_n_0,
   I1 => SIGMA_LCASE_1275_out_0_2,
   I2 => M_reg_14_1,
   I3 => x110_out_1,
   I4 => SIGMA_LCASE_0271_out_1,
   I5 => SIGMA_LCASE_1275_out_1,
   O => W_30_3_i_7_n_0
);
W_30_3_i_8 : LUT6
  generic map(
   INIT => X"566565566aa6a66a"
  )
 port map (
   I0 => W_30_3_i_4_n_0,
   I1 => M_reg_14_0,
   I2 => M_reg_15_18,
   I3 => M_reg_15_7,
   I4 => M_reg_15_3,
   I5 => x110_out_0,
   O => W_30_3_i_8_n_0
);
W_30_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_30_3_i_5_n_0,
   I1 => x100_out_10,
   I2 => x100_out_17,
   I3 => x100_out_19,
   O => W_30_3_i_9_n_0
);
W_30_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_14_6,
   I1 => x110_out_6,
   I2 => M_reg_15_24,
   I3 => M_reg_15_13,
   I4 => M_reg_15_9,
   O => W_30_7_i_10_n_0
);
W_30_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x110_out_5,
   I1 => M_reg_15_8,
   I2 => M_reg_15_12,
   I3 => M_reg_15_23,
   I4 => M_reg_14_5,
   O => W_30_7_i_11_n_0
);
W_30_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_14_5,
   I1 => x110_out_5,
   I2 => M_reg_15_23,
   I3 => M_reg_15_12,
   I4 => M_reg_15_8,
   O => W_30_7_i_12_n_0
);
W_30_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x110_out_4,
   I1 => M_reg_15_7,
   I2 => M_reg_15_11,
   I3 => M_reg_15_22,
   I4 => M_reg_14_4,
   O => W_30_7_i_13_n_0
);
W_30_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_14_4,
   I1 => x110_out_4,
   I2 => M_reg_15_22,
   I3 => M_reg_15_11,
   I4 => M_reg_15_7,
   O => W_30_7_i_14_n_0
);
W_30_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x110_out_3,
   I1 => M_reg_15_6,
   I2 => M_reg_15_10,
   I3 => M_reg_15_21,
   I4 => M_reg_14_3,
   O => W_30_7_i_15_n_0
);
W_30_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_14_3,
   I1 => x110_out_3,
   I2 => M_reg_15_21,
   I3 => M_reg_15_10,
   I4 => M_reg_15_6,
   O => W_30_7_i_16_n_0
);
W_30_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x110_out_2,
   I1 => M_reg_15_5,
   I2 => M_reg_15_9,
   I3 => M_reg_15_20,
   I4 => M_reg_14_2,
   O => W_30_7_i_17_n_0
);
W_30_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x100_out_16,
   I1 => x100_out_23,
   I2 => x100_out_25,
   I3 => W_30_7_i_10_n_0,
   I4 => W_30_7_i_11_n_0,
   O => W_30_7_i_2_n_0
);
W_30_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x100_out_15,
   I1 => x100_out_22,
   I2 => x100_out_24,
   I3 => W_30_7_i_12_n_0,
   I4 => W_30_7_i_13_n_0,
   O => W_30_7_i_3_n_0
);
W_30_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x100_out_14,
   I1 => x100_out_21,
   I2 => x100_out_23,
   I3 => W_30_7_i_14_n_0,
   I4 => W_30_7_i_15_n_0,
   O => W_30_7_i_4_n_0
);
W_30_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x100_out_13,
   I1 => x100_out_20,
   I2 => x100_out_22,
   I3 => W_30_7_i_16_n_0,
   I4 => W_30_7_i_17_n_0,
   O => W_30_7_i_5_n_0
);
W_30_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_30_7_i_2_n_0,
   I1 => W_30_11_i_16_n_0,
   I2 => x100_out_17,
   I3 => x100_out_24,
   I4 => x100_out_26,
   I5 => W_30_11_i_17_n_0,
   O => W_30_7_i_6_n_0
);
W_30_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_30_7_i_3_n_0,
   I1 => W_30_7_i_10_n_0,
   I2 => x100_out_16,
   I3 => x100_out_23,
   I4 => x100_out_25,
   I5 => W_30_7_i_11_n_0,
   O => W_30_7_i_7_n_0
);
W_30_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_30_7_i_4_n_0,
   I1 => W_30_7_i_12_n_0,
   I2 => x100_out_15,
   I3 => x100_out_22,
   I4 => x100_out_24,
   I5 => W_30_7_i_13_n_0,
   O => W_30_7_i_8_n_0
);
W_30_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_30_7_i_5_n_0,
   I1 => W_30_7_i_14_n_0,
   I2 => x100_out_14,
   I3 => x100_out_21,
   I4 => x100_out_23,
   I5 => W_30_7_i_15_n_0,
   O => W_30_7_i_9_n_0
);
W_31_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_15_10,
   I1 => x108_out_10,
   I2 => x117_out_28,
   I3 => x117_out_17,
   I4 => x117_out_13,
   O => W_31_11_i_10_n_0
);
W_31_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x108_out_9,
   I1 => x117_out_12,
   I2 => x117_out_16,
   I3 => x117_out_27,
   I4 => M_reg_15_9,
   O => W_31_11_i_11_n_0
);
W_31_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_15_9,
   I1 => x108_out_9,
   I2 => x117_out_27,
   I3 => x117_out_16,
   I4 => x117_out_12,
   O => W_31_11_i_12_n_0
);
W_31_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x108_out_8,
   I1 => x117_out_11,
   I2 => x117_out_15,
   I3 => x117_out_26,
   I4 => M_reg_15_8,
   O => W_31_11_i_13_n_0
);
W_31_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_15_8,
   I1 => x108_out_8,
   I2 => x117_out_26,
   I3 => x117_out_15,
   I4 => x117_out_11,
   O => W_31_11_i_14_n_0
);
W_31_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x108_out_7,
   I1 => x117_out_10,
   I2 => x117_out_14,
   I3 => x117_out_25,
   I4 => M_reg_15_7,
   O => W_31_11_i_15_n_0
);
W_31_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_15_7,
   I1 => x108_out_7,
   I2 => x117_out_25,
   I3 => x117_out_14,
   I4 => x117_out_10,
   O => W_31_11_i_16_n_0
);
W_31_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x108_out_6,
   I1 => x117_out_9,
   I2 => x117_out_13,
   I3 => x117_out_24,
   I4 => M_reg_15_6,
   O => W_31_11_i_17_n_0
);
W_31_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x98_out_20,
   I1 => x98_out_27,
   I2 => x98_out_29,
   I3 => W_31_11_i_10_n_0,
   I4 => W_31_11_i_11_n_0,
   O => W_31_11_i_2_n_0
);
W_31_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x98_out_19,
   I1 => x98_out_26,
   I2 => x98_out_28,
   I3 => W_31_11_i_12_n_0,
   I4 => W_31_11_i_13_n_0,
   O => W_31_11_i_3_n_0
);
W_31_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x98_out_18,
   I1 => x98_out_25,
   I2 => x98_out_27,
   I3 => W_31_11_i_14_n_0,
   I4 => W_31_11_i_15_n_0,
   O => W_31_11_i_4_n_0
);
W_31_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x98_out_17,
   I1 => x98_out_24,
   I2 => x98_out_26,
   I3 => W_31_11_i_16_n_0,
   I4 => W_31_11_i_17_n_0,
   O => W_31_11_i_5_n_0
);
W_31_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_31_11_i_2_n_0,
   I1 => W_31_15_i_16_n_0,
   I2 => x98_out_21,
   I3 => x98_out_28,
   I4 => x98_out_30,
   I5 => W_31_15_i_17_n_0,
   O => W_31_11_i_6_n_0
);
W_31_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_31_11_i_3_n_0,
   I1 => W_31_11_i_10_n_0,
   I2 => x98_out_20,
   I3 => x98_out_27,
   I4 => x98_out_29,
   I5 => W_31_11_i_11_n_0,
   O => W_31_11_i_7_n_0
);
W_31_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_31_11_i_4_n_0,
   I1 => W_31_11_i_12_n_0,
   I2 => x98_out_19,
   I3 => x98_out_26,
   I4 => x98_out_28,
   I5 => W_31_11_i_13_n_0,
   O => W_31_11_i_8_n_0
);
W_31_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_31_11_i_5_n_0,
   I1 => W_31_11_i_14_n_0,
   I2 => x98_out_18,
   I3 => x98_out_25,
   I4 => x98_out_27,
   I5 => W_31_11_i_15_n_0,
   O => W_31_11_i_9_n_0
);
W_31_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_15_14,
   I1 => x108_out_14,
   I2 => x117_out_0,
   I3 => x117_out_21,
   I4 => x117_out_17,
   O => W_31_15_i_10_n_0
);
W_31_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x108_out_13,
   I1 => x117_out_16,
   I2 => x117_out_20,
   I3 => x117_out_31,
   I4 => M_reg_15_13,
   O => W_31_15_i_11_n_0
);
W_31_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_15_13,
   I1 => x108_out_13,
   I2 => x117_out_31,
   I3 => x117_out_20,
   I4 => x117_out_16,
   O => W_31_15_i_12_n_0
);
W_31_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x108_out_12,
   I1 => x117_out_15,
   I2 => x117_out_19,
   I3 => x117_out_30,
   I4 => M_reg_15_12,
   O => W_31_15_i_13_n_0
);
W_31_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_15_12,
   I1 => x108_out_12,
   I2 => x117_out_30,
   I3 => x117_out_19,
   I4 => x117_out_15,
   O => W_31_15_i_14_n_0
);
W_31_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x108_out_11,
   I1 => x117_out_14,
   I2 => x117_out_18,
   I3 => x117_out_29,
   I4 => M_reg_15_11,
   O => W_31_15_i_15_n_0
);
W_31_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_15_11,
   I1 => x108_out_11,
   I2 => x117_out_29,
   I3 => x117_out_18,
   I4 => x117_out_14,
   O => W_31_15_i_16_n_0
);
W_31_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x108_out_10,
   I1 => x117_out_13,
   I2 => x117_out_17,
   I3 => x117_out_28,
   I4 => M_reg_15_10,
   O => W_31_15_i_17_n_0
);
W_31_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x98_out_24,
   I1 => x98_out_31,
   I2 => x98_out_1,
   I3 => W_31_15_i_10_n_0,
   I4 => W_31_15_i_11_n_0,
   O => W_31_15_i_2_n_0
);
W_31_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x98_out_23,
   I1 => x98_out_30,
   I2 => x98_out_0,
   I3 => W_31_15_i_12_n_0,
   I4 => W_31_15_i_13_n_0,
   O => W_31_15_i_3_n_0
);
W_31_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x98_out_22,
   I1 => x98_out_29,
   I2 => x98_out_31,
   I3 => W_31_15_i_14_n_0,
   I4 => W_31_15_i_15_n_0,
   O => W_31_15_i_4_n_0
);
W_31_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x98_out_21,
   I1 => x98_out_28,
   I2 => x98_out_30,
   I3 => W_31_15_i_16_n_0,
   I4 => W_31_15_i_17_n_0,
   O => W_31_15_i_5_n_0
);
W_31_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_31_15_i_2_n_0,
   I1 => W_31_19_i_16_n_0,
   I2 => x98_out_25,
   I3 => x98_out_0,
   I4 => x98_out_2,
   I5 => W_31_19_i_17_n_0,
   O => W_31_15_i_6_n_0
);
W_31_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_31_15_i_3_n_0,
   I1 => W_31_15_i_10_n_0,
   I2 => x98_out_24,
   I3 => x98_out_31,
   I4 => x98_out_1,
   I5 => W_31_15_i_11_n_0,
   O => W_31_15_i_7_n_0
);
W_31_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_31_15_i_4_n_0,
   I1 => W_31_15_i_12_n_0,
   I2 => x98_out_23,
   I3 => x98_out_30,
   I4 => x98_out_0,
   I5 => W_31_15_i_13_n_0,
   O => W_31_15_i_8_n_0
);
W_31_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_31_15_i_5_n_0,
   I1 => W_31_15_i_14_n_0,
   I2 => x98_out_22,
   I3 => x98_out_29,
   I4 => x98_out_31,
   I5 => W_31_15_i_15_n_0,
   O => W_31_15_i_9_n_0
);
W_31_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_15_18,
   I1 => x108_out_18,
   I2 => x117_out_4,
   I3 => x117_out_25,
   I4 => x117_out_21,
   O => W_31_19_i_10_n_0
);
W_31_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x108_out_17,
   I1 => x117_out_20,
   I2 => x117_out_24,
   I3 => x117_out_3,
   I4 => M_reg_15_17,
   O => W_31_19_i_11_n_0
);
W_31_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_15_17,
   I1 => x108_out_17,
   I2 => x117_out_3,
   I3 => x117_out_24,
   I4 => x117_out_20,
   O => W_31_19_i_12_n_0
);
W_31_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x108_out_16,
   I1 => x117_out_19,
   I2 => x117_out_23,
   I3 => x117_out_2,
   I4 => M_reg_15_16,
   O => W_31_19_i_13_n_0
);
W_31_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_15_16,
   I1 => x108_out_16,
   I2 => x117_out_2,
   I3 => x117_out_23,
   I4 => x117_out_19,
   O => W_31_19_i_14_n_0
);
W_31_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x108_out_15,
   I1 => x117_out_18,
   I2 => x117_out_22,
   I3 => x117_out_1,
   I4 => M_reg_15_15,
   O => W_31_19_i_15_n_0
);
W_31_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_15_15,
   I1 => x108_out_15,
   I2 => x117_out_1,
   I3 => x117_out_22,
   I4 => x117_out_18,
   O => W_31_19_i_16_n_0
);
W_31_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x108_out_14,
   I1 => x117_out_17,
   I2 => x117_out_21,
   I3 => x117_out_0,
   I4 => M_reg_15_14,
   O => W_31_19_i_17_n_0
);
W_31_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x98_out_28,
   I1 => x98_out_3,
   I2 => x98_out_5,
   I3 => W_31_19_i_10_n_0,
   I4 => W_31_19_i_11_n_0,
   O => W_31_19_i_2_n_0
);
W_31_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x98_out_27,
   I1 => x98_out_2,
   I2 => x98_out_4,
   I3 => W_31_19_i_12_n_0,
   I4 => W_31_19_i_13_n_0,
   O => W_31_19_i_3_n_0
);
W_31_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x98_out_26,
   I1 => x98_out_1,
   I2 => x98_out_3,
   I3 => W_31_19_i_14_n_0,
   I4 => W_31_19_i_15_n_0,
   O => W_31_19_i_4_n_0
);
W_31_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x98_out_25,
   I1 => x98_out_0,
   I2 => x98_out_2,
   I3 => W_31_19_i_16_n_0,
   I4 => W_31_19_i_17_n_0,
   O => W_31_19_i_5_n_0
);
W_31_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_31_19_i_2_n_0,
   I1 => W_31_23_i_16_n_0,
   I2 => x98_out_29,
   I3 => x98_out_4,
   I4 => x98_out_6,
   I5 => W_31_23_i_17_n_0,
   O => W_31_19_i_6_n_0
);
W_31_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_31_19_i_3_n_0,
   I1 => W_31_19_i_10_n_0,
   I2 => x98_out_28,
   I3 => x98_out_3,
   I4 => x98_out_5,
   I5 => W_31_19_i_11_n_0,
   O => W_31_19_i_7_n_0
);
W_31_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_31_19_i_4_n_0,
   I1 => W_31_19_i_12_n_0,
   I2 => x98_out_27,
   I3 => x98_out_2,
   I4 => x98_out_4,
   I5 => W_31_19_i_13_n_0,
   O => W_31_19_i_8_n_0
);
W_31_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_31_19_i_5_n_0,
   I1 => W_31_19_i_14_n_0,
   I2 => x98_out_26,
   I3 => x98_out_1,
   I4 => x98_out_3,
   I5 => W_31_19_i_15_n_0,
   O => W_31_19_i_9_n_0
);
W_31_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_15_22,
   I1 => x108_out_22,
   I2 => x117_out_8,
   I3 => x117_out_29,
   I4 => x117_out_25,
   O => W_31_23_i_10_n_0
);
W_31_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x108_out_21,
   I1 => x117_out_24,
   I2 => x117_out_28,
   I3 => x117_out_7,
   I4 => M_reg_15_21,
   O => W_31_23_i_11_n_0
);
W_31_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_15_21,
   I1 => x108_out_21,
   I2 => x117_out_7,
   I3 => x117_out_28,
   I4 => x117_out_24,
   O => W_31_23_i_12_n_0
);
W_31_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x108_out_20,
   I1 => x117_out_23,
   I2 => x117_out_27,
   I3 => x117_out_6,
   I4 => M_reg_15_20,
   O => W_31_23_i_13_n_0
);
W_31_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_15_20,
   I1 => x108_out_20,
   I2 => x117_out_6,
   I3 => x117_out_27,
   I4 => x117_out_23,
   O => W_31_23_i_14_n_0
);
W_31_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x108_out_19,
   I1 => x117_out_22,
   I2 => x117_out_26,
   I3 => x117_out_5,
   I4 => M_reg_15_19,
   O => W_31_23_i_15_n_0
);
W_31_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_15_19,
   I1 => x108_out_19,
   I2 => x117_out_5,
   I3 => x117_out_26,
   I4 => x117_out_22,
   O => W_31_23_i_16_n_0
);
W_31_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x108_out_18,
   I1 => x117_out_21,
   I2 => x117_out_25,
   I3 => x117_out_4,
   I4 => M_reg_15_18,
   O => W_31_23_i_17_n_0
);
W_31_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x98_out_7,
   I1 => x98_out_9,
   I2 => W_31_23_i_10_n_0,
   I3 => W_31_23_i_11_n_0,
   O => W_31_23_i_2_n_0
);
W_31_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x98_out_31,
   I1 => x98_out_6,
   I2 => x98_out_8,
   I3 => W_31_23_i_12_n_0,
   I4 => W_31_23_i_13_n_0,
   O => W_31_23_i_3_n_0
);
W_31_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x98_out_30,
   I1 => x98_out_5,
   I2 => x98_out_7,
   I3 => W_31_23_i_14_n_0,
   I4 => W_31_23_i_15_n_0,
   O => W_31_23_i_4_n_0
);
W_31_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x98_out_29,
   I1 => x98_out_4,
   I2 => x98_out_6,
   I3 => W_31_23_i_16_n_0,
   I4 => W_31_23_i_17_n_0,
   O => W_31_23_i_5_n_0
);
W_31_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x98_out_8,
   I1 => x98_out_10,
   I2 => W_31_27_i_16_n_0,
   I3 => W_31_27_i_17_n_0,
   I4 => W_31_23_i_2_n_0,
   O => W_31_23_i_6_n_0
);
W_31_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x98_out_7,
   I1 => x98_out_9,
   I2 => W_31_23_i_10_n_0,
   I3 => W_31_23_i_11_n_0,
   I4 => W_31_23_i_3_n_0,
   O => W_31_23_i_7_n_0
);
W_31_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_31_23_i_4_n_0,
   I1 => W_31_23_i_12_n_0,
   I2 => x98_out_31,
   I3 => x98_out_6,
   I4 => x98_out_8,
   I5 => W_31_23_i_13_n_0,
   O => W_31_23_i_8_n_0
);
W_31_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_31_23_i_5_n_0,
   I1 => W_31_23_i_14_n_0,
   I2 => x98_out_30,
   I3 => x98_out_5,
   I4 => x98_out_7,
   I5 => W_31_23_i_15_n_0,
   O => W_31_23_i_9_n_0
);
W_31_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_15_26,
   I1 => x108_out_26,
   I2 => x117_out_12,
   I3 => x117_out_1,
   I4 => x117_out_29,
   O => W_31_27_i_10_n_0
);
W_31_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x108_out_25,
   I1 => x117_out_28,
   I2 => x117_out_0,
   I3 => x117_out_11,
   I4 => M_reg_15_25,
   O => W_31_27_i_11_n_0
);
W_31_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_15_25,
   I1 => x108_out_25,
   I2 => x117_out_11,
   I3 => x117_out_0,
   I4 => x117_out_28,
   O => W_31_27_i_12_n_0
);
W_31_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x108_out_24,
   I1 => x117_out_27,
   I2 => x117_out_31,
   I3 => x117_out_10,
   I4 => M_reg_15_24,
   O => W_31_27_i_13_n_0
);
W_31_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_15_24,
   I1 => x108_out_24,
   I2 => x117_out_10,
   I3 => x117_out_31,
   I4 => x117_out_27,
   O => W_31_27_i_14_n_0
);
W_31_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x108_out_23,
   I1 => x117_out_26,
   I2 => x117_out_30,
   I3 => x117_out_9,
   I4 => M_reg_15_23,
   O => W_31_27_i_15_n_0
);
W_31_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_15_23,
   I1 => x108_out_23,
   I2 => x117_out_9,
   I3 => x117_out_30,
   I4 => x117_out_26,
   O => W_31_27_i_16_n_0
);
W_31_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x108_out_22,
   I1 => x117_out_25,
   I2 => x117_out_29,
   I3 => x117_out_8,
   I4 => M_reg_15_22,
   O => W_31_27_i_17_n_0
);
W_31_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x98_out_11,
   I1 => x98_out_13,
   I2 => W_31_27_i_10_n_0,
   I3 => W_31_27_i_11_n_0,
   O => W_31_27_i_2_n_0
);
W_31_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x98_out_10,
   I1 => x98_out_12,
   I2 => W_31_27_i_12_n_0,
   I3 => W_31_27_i_13_n_0,
   O => W_31_27_i_3_n_0
);
W_31_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x98_out_9,
   I1 => x98_out_11,
   I2 => W_31_27_i_14_n_0,
   I3 => W_31_27_i_15_n_0,
   O => W_31_27_i_4_n_0
);
W_31_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x98_out_8,
   I1 => x98_out_10,
   I2 => W_31_27_i_16_n_0,
   I3 => W_31_27_i_17_n_0,
   O => W_31_27_i_5_n_0
);
W_31_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x98_out_12,
   I1 => x98_out_14,
   I2 => W_31_31_i_13_n_0,
   I3 => W_31_31_i_14_n_0,
   I4 => W_31_27_i_2_n_0,
   O => W_31_27_i_6_n_0
);
W_31_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x98_out_11,
   I1 => x98_out_13,
   I2 => W_31_27_i_10_n_0,
   I3 => W_31_27_i_11_n_0,
   I4 => W_31_27_i_3_n_0,
   O => W_31_27_i_7_n_0
);
W_31_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x98_out_10,
   I1 => x98_out_12,
   I2 => W_31_27_i_12_n_0,
   I3 => W_31_27_i_13_n_0,
   I4 => W_31_27_i_4_n_0,
   O => W_31_27_i_8_n_0
);
W_31_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x98_out_9,
   I1 => x98_out_11,
   I2 => W_31_27_i_14_n_0,
   I3 => W_31_27_i_15_n_0,
   I4 => W_31_27_i_5_n_0,
   O => W_31_27_i_9_n_0
);
W_31_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x108_out_28,
   I1 => x117_out_31,
   I2 => x117_out_3,
   I3 => x117_out_14,
   I4 => M_reg_15_28,
   O => W_31_31_i_10_n_0
);
W_31_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_15_28,
   I1 => x108_out_28,
   I2 => x117_out_14,
   I3 => x117_out_3,
   I4 => x117_out_31,
   O => W_31_31_i_11_n_0
);
W_31_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x108_out_27,
   I1 => x117_out_30,
   I2 => x117_out_2,
   I3 => x117_out_13,
   I4 => M_reg_15_27,
   O => W_31_31_i_12_n_0
);
W_31_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_15_27,
   I1 => x108_out_27,
   I2 => x117_out_13,
   I3 => x117_out_2,
   I4 => x117_out_30,
   O => W_31_31_i_13_n_0
);
W_31_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x108_out_26,
   I1 => x117_out_29,
   I2 => x117_out_1,
   I3 => x117_out_12,
   I4 => M_reg_15_26,
   O => W_31_31_i_14_n_0
);
W_31_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x108_out_29,
   I1 => x117_out_4,
   I2 => x117_out_15,
   I3 => M_reg_15_29,
   O => W_31_31_i_15_n_0
);
W_31_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x98_out_17,
   I1 => x98_out_15,
   O => SIGMA_LCASE_1267_out_0_30
);
W_31_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => x117_out_6,
   I1 => x117_out_17,
   I2 => x108_out_31,
   I3 => M_reg_15_31,
   I4 => x98_out_16,
   I5 => x98_out_18,
   O => W_31_31_i_17_n_0
);
W_31_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x117_out_16,
   I1 => x117_out_5,
   O => SIGMA_LCASE_0263_out_30
);
W_31_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => M_reg_15_30,
   I1 => x108_out_30,
   I2 => x117_out_16,
   I3 => x117_out_5,
   O => W_31_31_i_19_n_0
);
W_31_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x98_out_14,
   I1 => x98_out_16,
   I2 => W_31_31_i_9_n_0,
   I3 => W_31_31_i_10_n_0,
   O => W_31_31_i_2_n_0
);
W_31_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x98_out_13,
   I1 => x98_out_15,
   I2 => W_31_31_i_11_n_0,
   I3 => W_31_31_i_12_n_0,
   O => W_31_31_i_3_n_0
);
W_31_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x98_out_12,
   I1 => x98_out_14,
   I2 => W_31_31_i_13_n_0,
   I3 => W_31_31_i_14_n_0,
   O => W_31_31_i_4_n_0
);
W_31_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_31_31_i_15_n_0,
   I1 => SIGMA_LCASE_1267_out_0_30,
   I2 => W_31_31_i_17_n_0,
   I3 => x108_out_30,
   I4 => SIGMA_LCASE_0263_out_30,
   I5 => M_reg_15_30,
   O => W_31_31_i_5_n_0
);
W_31_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_31_31_i_2_n_0,
   I1 => W_31_31_i_19_n_0,
   I2 => x98_out_15,
   I3 => x98_out_17,
   I4 => W_31_31_i_15_n_0,
   O => W_31_31_i_6_n_0
);
W_31_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x98_out_14,
   I1 => x98_out_16,
   I2 => W_31_31_i_9_n_0,
   I3 => W_31_31_i_10_n_0,
   I4 => W_31_31_i_3_n_0,
   O => W_31_31_i_7_n_0
);
W_31_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x98_out_13,
   I1 => x98_out_15,
   I2 => W_31_31_i_11_n_0,
   I3 => W_31_31_i_12_n_0,
   I4 => W_31_31_i_4_n_0,
   O => W_31_31_i_8_n_0
);
W_31_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => M_reg_15_29,
   I1 => x108_out_29,
   I2 => x117_out_15,
   I3 => x117_out_4,
   O => W_31_31_i_9_n_0
);
W_31_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_15_2,
   I1 => x108_out_2,
   I2 => x117_out_20,
   I3 => x117_out_9,
   I4 => x117_out_5,
   O => W_31_3_i_10_n_0
);
W_31_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x108_out_1,
   I1 => x117_out_4,
   I2 => x117_out_8,
   I3 => x117_out_19,
   I4 => M_reg_15_1,
   O => W_31_3_i_11_n_0
);
W_31_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x117_out_19,
   I1 => x117_out_8,
   I2 => x117_out_4,
   O => SIGMA_LCASE_0263_out_1
);
W_31_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x98_out_21,
   I1 => x98_out_19,
   I2 => x98_out_12,
   O => SIGMA_LCASE_1267_out_0_2
);
W_31_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x98_out_20,
   I1 => x98_out_18,
   I2 => x98_out_11,
   O => SIGMA_LCASE_1267_out_1
);
W_31_3_i_15 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_15_1,
   I1 => x108_out_1,
   I2 => x117_out_19,
   I3 => x117_out_8,
   I4 => x117_out_4,
   O => W_31_3_i_15_n_0
);
W_31_3_i_16 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x117_out_18,
   I1 => x117_out_7,
   I2 => x117_out_3,
   O => SIGMA_LCASE_0263_out_0
);
W_31_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x98_out_12,
   I1 => x98_out_19,
   I2 => x98_out_21,
   I3 => W_31_3_i_10_n_0,
   I4 => W_31_3_i_11_n_0,
   O => W_31_3_i_2_n_0
);
W_31_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_31_3_i_11_n_0,
   I1 => x98_out_21,
   I2 => x98_out_19,
   I3 => x98_out_12,
   I4 => W_31_3_i_10_n_0,
   O => W_31_3_i_3_n_0
);
W_31_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_0263_out_1,
   I1 => x108_out_1,
   I2 => M_reg_15_1,
   I3 => x98_out_11,
   I4 => x98_out_18,
   I5 => x98_out_20,
   O => W_31_3_i_4_n_0
);
W_31_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_15_0,
   I1 => x108_out_0,
   I2 => x117_out_18,
   I3 => x117_out_7,
   I4 => x117_out_3,
   O => W_31_3_i_5_n_0
);
W_31_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_31_3_i_2_n_0,
   I1 => W_31_7_i_16_n_0,
   I2 => x98_out_13,
   I3 => x98_out_20,
   I4 => x98_out_22,
   I5 => W_31_7_i_17_n_0,
   O => W_31_3_i_6_n_0
);
W_31_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_31_3_i_10_n_0,
   I1 => SIGMA_LCASE_1267_out_0_2,
   I2 => M_reg_15_1,
   I3 => x108_out_1,
   I4 => SIGMA_LCASE_0263_out_1,
   I5 => SIGMA_LCASE_1267_out_1,
   O => W_31_3_i_7_n_0
);
W_31_3_i_8 : LUT5
  generic map(
   INIT => X"99969666"
  )
 port map (
   I0 => SIGMA_LCASE_1267_out_1,
   I1 => W_31_3_i_15_n_0,
   I2 => M_reg_15_0,
   I3 => SIGMA_LCASE_0263_out_0,
   I4 => x108_out_0,
   O => W_31_3_i_8_n_0
);
W_31_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_31_3_i_5_n_0,
   I1 => x98_out_10,
   I2 => x98_out_17,
   I3 => x98_out_19,
   O => W_31_3_i_9_n_0
);
W_31_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_15_6,
   I1 => x108_out_6,
   I2 => x117_out_24,
   I3 => x117_out_13,
   I4 => x117_out_9,
   O => W_31_7_i_10_n_0
);
W_31_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x108_out_5,
   I1 => x117_out_8,
   I2 => x117_out_12,
   I3 => x117_out_23,
   I4 => M_reg_15_5,
   O => W_31_7_i_11_n_0
);
W_31_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_15_5,
   I1 => x108_out_5,
   I2 => x117_out_23,
   I3 => x117_out_12,
   I4 => x117_out_8,
   O => W_31_7_i_12_n_0
);
W_31_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x108_out_4,
   I1 => x117_out_7,
   I2 => x117_out_11,
   I3 => x117_out_22,
   I4 => M_reg_15_4,
   O => W_31_7_i_13_n_0
);
W_31_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_15_4,
   I1 => x108_out_4,
   I2 => x117_out_22,
   I3 => x117_out_11,
   I4 => x117_out_7,
   O => W_31_7_i_14_n_0
);
W_31_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x108_out_3,
   I1 => x117_out_6,
   I2 => x117_out_10,
   I3 => x117_out_21,
   I4 => M_reg_15_3,
   O => W_31_7_i_15_n_0
);
W_31_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => M_reg_15_3,
   I1 => x108_out_3,
   I2 => x117_out_21,
   I3 => x117_out_10,
   I4 => x117_out_6,
   O => W_31_7_i_16_n_0
);
W_31_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x108_out_2,
   I1 => x117_out_5,
   I2 => x117_out_9,
   I3 => x117_out_20,
   I4 => M_reg_15_2,
   O => W_31_7_i_17_n_0
);
W_31_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x98_out_16,
   I1 => x98_out_23,
   I2 => x98_out_25,
   I3 => W_31_7_i_10_n_0,
   I4 => W_31_7_i_11_n_0,
   O => W_31_7_i_2_n_0
);
W_31_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x98_out_15,
   I1 => x98_out_22,
   I2 => x98_out_24,
   I3 => W_31_7_i_12_n_0,
   I4 => W_31_7_i_13_n_0,
   O => W_31_7_i_3_n_0
);
W_31_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x98_out_14,
   I1 => x98_out_21,
   I2 => x98_out_23,
   I3 => W_31_7_i_14_n_0,
   I4 => W_31_7_i_15_n_0,
   O => W_31_7_i_4_n_0
);
W_31_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x98_out_13,
   I1 => x98_out_20,
   I2 => x98_out_22,
   I3 => W_31_7_i_16_n_0,
   I4 => W_31_7_i_17_n_0,
   O => W_31_7_i_5_n_0
);
W_31_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_31_7_i_2_n_0,
   I1 => W_31_11_i_16_n_0,
   I2 => x98_out_17,
   I3 => x98_out_24,
   I4 => x98_out_26,
   I5 => W_31_11_i_17_n_0,
   O => W_31_7_i_6_n_0
);
W_31_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_31_7_i_3_n_0,
   I1 => W_31_7_i_10_n_0,
   I2 => x98_out_16,
   I3 => x98_out_23,
   I4 => x98_out_25,
   I5 => W_31_7_i_11_n_0,
   O => W_31_7_i_7_n_0
);
W_31_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_31_7_i_4_n_0,
   I1 => W_31_7_i_12_n_0,
   I2 => x98_out_15,
   I3 => x98_out_22,
   I4 => x98_out_24,
   I5 => W_31_7_i_13_n_0,
   O => W_31_7_i_8_n_0
);
W_31_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_31_7_i_5_n_0,
   I1 => W_31_7_i_14_n_0,
   I2 => x98_out_14,
   I3 => x98_out_21,
   I4 => x98_out_23,
   I5 => W_31_7_i_15_n_0,
   O => W_31_7_i_9_n_0
);
W_32_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x117_out_10,
   I1 => x106_out_10,
   I2 => x116_out_28,
   I3 => x116_out_17,
   I4 => x116_out_13,
   O => W_32_11_i_10_n_0
);
W_32_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x106_out_9,
   I1 => x116_out_12,
   I2 => x116_out_16,
   I3 => x116_out_27,
   I4 => x117_out_9,
   O => W_32_11_i_11_n_0
);
W_32_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x117_out_9,
   I1 => x106_out_9,
   I2 => x116_out_27,
   I3 => x116_out_16,
   I4 => x116_out_12,
   O => W_32_11_i_12_n_0
);
W_32_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x106_out_8,
   I1 => x116_out_11,
   I2 => x116_out_15,
   I3 => x116_out_26,
   I4 => x117_out_8,
   O => W_32_11_i_13_n_0
);
W_32_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x117_out_8,
   I1 => x106_out_8,
   I2 => x116_out_26,
   I3 => x116_out_15,
   I4 => x116_out_11,
   O => W_32_11_i_14_n_0
);
W_32_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x106_out_7,
   I1 => x116_out_10,
   I2 => x116_out_14,
   I3 => x116_out_25,
   I4 => x117_out_7,
   O => W_32_11_i_15_n_0
);
W_32_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x117_out_7,
   I1 => x106_out_7,
   I2 => x116_out_25,
   I3 => x116_out_14,
   I4 => x116_out_10,
   O => W_32_11_i_16_n_0
);
W_32_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x106_out_6,
   I1 => x116_out_9,
   I2 => x116_out_13,
   I3 => x116_out_24,
   I4 => x117_out_6,
   O => W_32_11_i_17_n_0
);
W_32_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x96_out_20,
   I1 => x96_out_27,
   I2 => x96_out_29,
   I3 => W_32_11_i_10_n_0,
   I4 => W_32_11_i_11_n_0,
   O => W_32_11_i_2_n_0
);
W_32_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x96_out_19,
   I1 => x96_out_26,
   I2 => x96_out_28,
   I3 => W_32_11_i_12_n_0,
   I4 => W_32_11_i_13_n_0,
   O => W_32_11_i_3_n_0
);
W_32_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x96_out_18,
   I1 => x96_out_25,
   I2 => x96_out_27,
   I3 => W_32_11_i_14_n_0,
   I4 => W_32_11_i_15_n_0,
   O => W_32_11_i_4_n_0
);
W_32_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x96_out_17,
   I1 => x96_out_24,
   I2 => x96_out_26,
   I3 => W_32_11_i_16_n_0,
   I4 => W_32_11_i_17_n_0,
   O => W_32_11_i_5_n_0
);
W_32_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_32_11_i_2_n_0,
   I1 => W_32_15_i_16_n_0,
   I2 => x96_out_21,
   I3 => x96_out_28,
   I4 => x96_out_30,
   I5 => W_32_15_i_17_n_0,
   O => W_32_11_i_6_n_0
);
W_32_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_32_11_i_3_n_0,
   I1 => W_32_11_i_10_n_0,
   I2 => x96_out_20,
   I3 => x96_out_27,
   I4 => x96_out_29,
   I5 => W_32_11_i_11_n_0,
   O => W_32_11_i_7_n_0
);
W_32_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_32_11_i_4_n_0,
   I1 => W_32_11_i_12_n_0,
   I2 => x96_out_19,
   I3 => x96_out_26,
   I4 => x96_out_28,
   I5 => W_32_11_i_13_n_0,
   O => W_32_11_i_8_n_0
);
W_32_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_32_11_i_5_n_0,
   I1 => W_32_11_i_14_n_0,
   I2 => x96_out_18,
   I3 => x96_out_25,
   I4 => x96_out_27,
   I5 => W_32_11_i_15_n_0,
   O => W_32_11_i_9_n_0
);
W_32_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x117_out_14,
   I1 => x106_out_14,
   I2 => x116_out_0,
   I3 => x116_out_21,
   I4 => x116_out_17,
   O => W_32_15_i_10_n_0
);
W_32_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x106_out_13,
   I1 => x116_out_16,
   I2 => x116_out_20,
   I3 => x116_out_31,
   I4 => x117_out_13,
   O => W_32_15_i_11_n_0
);
W_32_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x117_out_13,
   I1 => x106_out_13,
   I2 => x116_out_31,
   I3 => x116_out_20,
   I4 => x116_out_16,
   O => W_32_15_i_12_n_0
);
W_32_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x106_out_12,
   I1 => x116_out_15,
   I2 => x116_out_19,
   I3 => x116_out_30,
   I4 => x117_out_12,
   O => W_32_15_i_13_n_0
);
W_32_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x117_out_12,
   I1 => x106_out_12,
   I2 => x116_out_30,
   I3 => x116_out_19,
   I4 => x116_out_15,
   O => W_32_15_i_14_n_0
);
W_32_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x106_out_11,
   I1 => x116_out_14,
   I2 => x116_out_18,
   I3 => x116_out_29,
   I4 => x117_out_11,
   O => W_32_15_i_15_n_0
);
W_32_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x117_out_11,
   I1 => x106_out_11,
   I2 => x116_out_29,
   I3 => x116_out_18,
   I4 => x116_out_14,
   O => W_32_15_i_16_n_0
);
W_32_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x106_out_10,
   I1 => x116_out_13,
   I2 => x116_out_17,
   I3 => x116_out_28,
   I4 => x117_out_10,
   O => W_32_15_i_17_n_0
);
W_32_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x96_out_24,
   I1 => x96_out_31,
   I2 => x96_out_1,
   I3 => W_32_15_i_10_n_0,
   I4 => W_32_15_i_11_n_0,
   O => W_32_15_i_2_n_0
);
W_32_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x96_out_23,
   I1 => x96_out_30,
   I2 => x96_out_0,
   I3 => W_32_15_i_12_n_0,
   I4 => W_32_15_i_13_n_0,
   O => W_32_15_i_3_n_0
);
W_32_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x96_out_22,
   I1 => x96_out_29,
   I2 => x96_out_31,
   I3 => W_32_15_i_14_n_0,
   I4 => W_32_15_i_15_n_0,
   O => W_32_15_i_4_n_0
);
W_32_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x96_out_21,
   I1 => x96_out_28,
   I2 => x96_out_30,
   I3 => W_32_15_i_16_n_0,
   I4 => W_32_15_i_17_n_0,
   O => W_32_15_i_5_n_0
);
W_32_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_32_15_i_2_n_0,
   I1 => W_32_19_i_16_n_0,
   I2 => x96_out_25,
   I3 => x96_out_0,
   I4 => x96_out_2,
   I5 => W_32_19_i_17_n_0,
   O => W_32_15_i_6_n_0
);
W_32_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_32_15_i_3_n_0,
   I1 => W_32_15_i_10_n_0,
   I2 => x96_out_24,
   I3 => x96_out_31,
   I4 => x96_out_1,
   I5 => W_32_15_i_11_n_0,
   O => W_32_15_i_7_n_0
);
W_32_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_32_15_i_4_n_0,
   I1 => W_32_15_i_12_n_0,
   I2 => x96_out_23,
   I3 => x96_out_30,
   I4 => x96_out_0,
   I5 => W_32_15_i_13_n_0,
   O => W_32_15_i_8_n_0
);
W_32_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_32_15_i_5_n_0,
   I1 => W_32_15_i_14_n_0,
   I2 => x96_out_22,
   I3 => x96_out_29,
   I4 => x96_out_31,
   I5 => W_32_15_i_15_n_0,
   O => W_32_15_i_9_n_0
);
W_32_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x117_out_18,
   I1 => x106_out_18,
   I2 => x116_out_4,
   I3 => x116_out_25,
   I4 => x116_out_21,
   O => W_32_19_i_10_n_0
);
W_32_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x106_out_17,
   I1 => x116_out_20,
   I2 => x116_out_24,
   I3 => x116_out_3,
   I4 => x117_out_17,
   O => W_32_19_i_11_n_0
);
W_32_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x117_out_17,
   I1 => x106_out_17,
   I2 => x116_out_3,
   I3 => x116_out_24,
   I4 => x116_out_20,
   O => W_32_19_i_12_n_0
);
W_32_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x106_out_16,
   I1 => x116_out_19,
   I2 => x116_out_23,
   I3 => x116_out_2,
   I4 => x117_out_16,
   O => W_32_19_i_13_n_0
);
W_32_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x117_out_16,
   I1 => x106_out_16,
   I2 => x116_out_2,
   I3 => x116_out_23,
   I4 => x116_out_19,
   O => W_32_19_i_14_n_0
);
W_32_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x106_out_15,
   I1 => x116_out_18,
   I2 => x116_out_22,
   I3 => x116_out_1,
   I4 => x117_out_15,
   O => W_32_19_i_15_n_0
);
W_32_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x117_out_15,
   I1 => x106_out_15,
   I2 => x116_out_1,
   I3 => x116_out_22,
   I4 => x116_out_18,
   O => W_32_19_i_16_n_0
);
W_32_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x106_out_14,
   I1 => x116_out_17,
   I2 => x116_out_21,
   I3 => x116_out_0,
   I4 => x117_out_14,
   O => W_32_19_i_17_n_0
);
W_32_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x96_out_28,
   I1 => x96_out_3,
   I2 => x96_out_5,
   I3 => W_32_19_i_10_n_0,
   I4 => W_32_19_i_11_n_0,
   O => W_32_19_i_2_n_0
);
W_32_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x96_out_27,
   I1 => x96_out_2,
   I2 => x96_out_4,
   I3 => W_32_19_i_12_n_0,
   I4 => W_32_19_i_13_n_0,
   O => W_32_19_i_3_n_0
);
W_32_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x96_out_26,
   I1 => x96_out_1,
   I2 => x96_out_3,
   I3 => W_32_19_i_14_n_0,
   I4 => W_32_19_i_15_n_0,
   O => W_32_19_i_4_n_0
);
W_32_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x96_out_25,
   I1 => x96_out_0,
   I2 => x96_out_2,
   I3 => W_32_19_i_16_n_0,
   I4 => W_32_19_i_17_n_0,
   O => W_32_19_i_5_n_0
);
W_32_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_32_19_i_2_n_0,
   I1 => W_32_23_i_16_n_0,
   I2 => x96_out_29,
   I3 => x96_out_4,
   I4 => x96_out_6,
   I5 => W_32_23_i_17_n_0,
   O => W_32_19_i_6_n_0
);
W_32_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_32_19_i_3_n_0,
   I1 => W_32_19_i_10_n_0,
   I2 => x96_out_28,
   I3 => x96_out_3,
   I4 => x96_out_5,
   I5 => W_32_19_i_11_n_0,
   O => W_32_19_i_7_n_0
);
W_32_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_32_19_i_4_n_0,
   I1 => W_32_19_i_12_n_0,
   I2 => x96_out_27,
   I3 => x96_out_2,
   I4 => x96_out_4,
   I5 => W_32_19_i_13_n_0,
   O => W_32_19_i_8_n_0
);
W_32_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_32_19_i_5_n_0,
   I1 => W_32_19_i_14_n_0,
   I2 => x96_out_26,
   I3 => x96_out_1,
   I4 => x96_out_3,
   I5 => W_32_19_i_15_n_0,
   O => W_32_19_i_9_n_0
);
W_32_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x117_out_22,
   I1 => x106_out_22,
   I2 => x116_out_8,
   I3 => x116_out_29,
   I4 => x116_out_25,
   O => W_32_23_i_10_n_0
);
W_32_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x106_out_21,
   I1 => x116_out_24,
   I2 => x116_out_28,
   I3 => x116_out_7,
   I4 => x117_out_21,
   O => W_32_23_i_11_n_0
);
W_32_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x117_out_21,
   I1 => x106_out_21,
   I2 => x116_out_7,
   I3 => x116_out_28,
   I4 => x116_out_24,
   O => W_32_23_i_12_n_0
);
W_32_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x106_out_20,
   I1 => x116_out_23,
   I2 => x116_out_27,
   I3 => x116_out_6,
   I4 => x117_out_20,
   O => W_32_23_i_13_n_0
);
W_32_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x117_out_20,
   I1 => x106_out_20,
   I2 => x116_out_6,
   I3 => x116_out_27,
   I4 => x116_out_23,
   O => W_32_23_i_14_n_0
);
W_32_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x106_out_19,
   I1 => x116_out_22,
   I2 => x116_out_26,
   I3 => x116_out_5,
   I4 => x117_out_19,
   O => W_32_23_i_15_n_0
);
W_32_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x117_out_19,
   I1 => x106_out_19,
   I2 => x116_out_5,
   I3 => x116_out_26,
   I4 => x116_out_22,
   O => W_32_23_i_16_n_0
);
W_32_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x106_out_18,
   I1 => x116_out_21,
   I2 => x116_out_25,
   I3 => x116_out_4,
   I4 => x117_out_18,
   O => W_32_23_i_17_n_0
);
W_32_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x96_out_7,
   I1 => x96_out_9,
   I2 => W_32_23_i_10_n_0,
   I3 => W_32_23_i_11_n_0,
   O => W_32_23_i_2_n_0
);
W_32_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x96_out_31,
   I1 => x96_out_6,
   I2 => x96_out_8,
   I3 => W_32_23_i_12_n_0,
   I4 => W_32_23_i_13_n_0,
   O => W_32_23_i_3_n_0
);
W_32_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x96_out_30,
   I1 => x96_out_5,
   I2 => x96_out_7,
   I3 => W_32_23_i_14_n_0,
   I4 => W_32_23_i_15_n_0,
   O => W_32_23_i_4_n_0
);
W_32_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x96_out_29,
   I1 => x96_out_4,
   I2 => x96_out_6,
   I3 => W_32_23_i_16_n_0,
   I4 => W_32_23_i_17_n_0,
   O => W_32_23_i_5_n_0
);
W_32_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x96_out_8,
   I1 => x96_out_10,
   I2 => W_32_27_i_16_n_0,
   I3 => W_32_27_i_17_n_0,
   I4 => W_32_23_i_2_n_0,
   O => W_32_23_i_6_n_0
);
W_32_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x96_out_7,
   I1 => x96_out_9,
   I2 => W_32_23_i_10_n_0,
   I3 => W_32_23_i_11_n_0,
   I4 => W_32_23_i_3_n_0,
   O => W_32_23_i_7_n_0
);
W_32_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_32_23_i_4_n_0,
   I1 => W_32_23_i_12_n_0,
   I2 => x96_out_31,
   I3 => x96_out_6,
   I4 => x96_out_8,
   I5 => W_32_23_i_13_n_0,
   O => W_32_23_i_8_n_0
);
W_32_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_32_23_i_5_n_0,
   I1 => W_32_23_i_14_n_0,
   I2 => x96_out_30,
   I3 => x96_out_5,
   I4 => x96_out_7,
   I5 => W_32_23_i_15_n_0,
   O => W_32_23_i_9_n_0
);
W_32_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x117_out_26,
   I1 => x106_out_26,
   I2 => x116_out_12,
   I3 => x116_out_1,
   I4 => x116_out_29,
   O => W_32_27_i_10_n_0
);
W_32_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x106_out_25,
   I1 => x116_out_28,
   I2 => x116_out_0,
   I3 => x116_out_11,
   I4 => x117_out_25,
   O => W_32_27_i_11_n_0
);
W_32_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x117_out_25,
   I1 => x106_out_25,
   I2 => x116_out_11,
   I3 => x116_out_0,
   I4 => x116_out_28,
   O => W_32_27_i_12_n_0
);
W_32_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x106_out_24,
   I1 => x116_out_27,
   I2 => x116_out_31,
   I3 => x116_out_10,
   I4 => x117_out_24,
   O => W_32_27_i_13_n_0
);
W_32_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x117_out_24,
   I1 => x106_out_24,
   I2 => x116_out_10,
   I3 => x116_out_31,
   I4 => x116_out_27,
   O => W_32_27_i_14_n_0
);
W_32_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x106_out_23,
   I1 => x116_out_26,
   I2 => x116_out_30,
   I3 => x116_out_9,
   I4 => x117_out_23,
   O => W_32_27_i_15_n_0
);
W_32_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x117_out_23,
   I1 => x106_out_23,
   I2 => x116_out_9,
   I3 => x116_out_30,
   I4 => x116_out_26,
   O => W_32_27_i_16_n_0
);
W_32_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x106_out_22,
   I1 => x116_out_25,
   I2 => x116_out_29,
   I3 => x116_out_8,
   I4 => x117_out_22,
   O => W_32_27_i_17_n_0
);
W_32_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x96_out_11,
   I1 => x96_out_13,
   I2 => W_32_27_i_10_n_0,
   I3 => W_32_27_i_11_n_0,
   O => W_32_27_i_2_n_0
);
W_32_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x96_out_10,
   I1 => x96_out_12,
   I2 => W_32_27_i_12_n_0,
   I3 => W_32_27_i_13_n_0,
   O => W_32_27_i_3_n_0
);
W_32_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x96_out_9,
   I1 => x96_out_11,
   I2 => W_32_27_i_14_n_0,
   I3 => W_32_27_i_15_n_0,
   O => W_32_27_i_4_n_0
);
W_32_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x96_out_8,
   I1 => x96_out_10,
   I2 => W_32_27_i_16_n_0,
   I3 => W_32_27_i_17_n_0,
   O => W_32_27_i_5_n_0
);
W_32_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x96_out_12,
   I1 => x96_out_14,
   I2 => W_32_31_i_14_n_0,
   I3 => W_32_31_i_15_n_0,
   I4 => W_32_27_i_2_n_0,
   O => W_32_27_i_6_n_0
);
W_32_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x96_out_11,
   I1 => x96_out_13,
   I2 => W_32_27_i_10_n_0,
   I3 => W_32_27_i_11_n_0,
   I4 => W_32_27_i_3_n_0,
   O => W_32_27_i_7_n_0
);
W_32_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x96_out_10,
   I1 => x96_out_12,
   I2 => W_32_27_i_12_n_0,
   I3 => W_32_27_i_13_n_0,
   I4 => W_32_27_i_4_n_0,
   O => W_32_27_i_8_n_0
);
W_32_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x96_out_9,
   I1 => x96_out_11,
   I2 => W_32_27_i_14_n_0,
   I3 => W_32_27_i_15_n_0,
   I4 => W_32_27_i_5_n_0,
   O => W_32_27_i_9_n_0
);
W_32_31_i_1 : LUT2
  generic map(
   INIT => X"2"
  )
 port map (
   I0 => W_32,
   I1 => rst_IBUF,
   O => W_reg_32_0
);
W_32_31_i_10 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x117_out_29,
   I1 => x106_out_29,
   I2 => x116_out_15,
   I3 => x116_out_4,
   O => W_32_31_i_10_n_0
);
W_32_31_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x106_out_28,
   I1 => x116_out_31,
   I2 => x116_out_3,
   I3 => x116_out_14,
   I4 => x117_out_28,
   O => W_32_31_i_11_n_0
);
W_32_31_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x117_out_28,
   I1 => x106_out_28,
   I2 => x116_out_14,
   I3 => x116_out_3,
   I4 => x116_out_31,
   O => W_32_31_i_12_n_0
);
W_32_31_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x106_out_27,
   I1 => x116_out_30,
   I2 => x116_out_2,
   I3 => x116_out_13,
   I4 => x117_out_27,
   O => W_32_31_i_13_n_0
);
W_32_31_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x117_out_27,
   I1 => x106_out_27,
   I2 => x116_out_13,
   I3 => x116_out_2,
   I4 => x116_out_30,
   O => W_32_31_i_14_n_0
);
W_32_31_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x106_out_26,
   I1 => x116_out_29,
   I2 => x116_out_1,
   I3 => x116_out_12,
   I4 => x117_out_26,
   O => W_32_31_i_15_n_0
);
W_32_31_i_16 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x106_out_29,
   I1 => x116_out_4,
   I2 => x116_out_15,
   I3 => x117_out_29,
   O => W_32_31_i_16_n_0
);
W_32_31_i_17 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x96_out_17,
   I1 => x96_out_15,
   O => SIGMA_LCASE_1259_out_0_30
);
W_32_31_i_18 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => x116_out_6,
   I1 => x116_out_17,
   I2 => x106_out_31,
   I3 => x117_out_31,
   I4 => x96_out_16,
   I5 => x96_out_18,
   O => W_32_31_i_18_n_0
);
W_32_31_i_19 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x116_out_16,
   I1 => x116_out_5,
   O => SIGMA_LCASE_0255_out_30
);
W_32_31_i_20 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x117_out_30,
   I1 => x106_out_30,
   I2 => x116_out_16,
   I3 => x116_out_5,
   O => W_32_31_i_20_n_0
);
W_32_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x96_out_14,
   I1 => x96_out_16,
   I2 => W_32_31_i_10_n_0,
   I3 => W_32_31_i_11_n_0,
   O => W_32_31_i_3_n_0
);
W_32_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x96_out_13,
   I1 => x96_out_15,
   I2 => W_32_31_i_12_n_0,
   I3 => W_32_31_i_13_n_0,
   O => W_32_31_i_4_n_0
);
W_32_31_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x96_out_12,
   I1 => x96_out_14,
   I2 => W_32_31_i_14_n_0,
   I3 => W_32_31_i_15_n_0,
   O => W_32_31_i_5_n_0
);
W_32_31_i_6 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_32_31_i_16_n_0,
   I1 => SIGMA_LCASE_1259_out_0_30,
   I2 => W_32_31_i_18_n_0,
   I3 => x106_out_30,
   I4 => SIGMA_LCASE_0255_out_30,
   I5 => x117_out_30,
   O => W_32_31_i_6_n_0
);
W_32_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_32_31_i_3_n_0,
   I1 => W_32_31_i_20_n_0,
   I2 => x96_out_15,
   I3 => x96_out_17,
   I4 => W_32_31_i_16_n_0,
   O => W_32_31_i_7_n_0
);
W_32_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x96_out_14,
   I1 => x96_out_16,
   I2 => W_32_31_i_10_n_0,
   I3 => W_32_31_i_11_n_0,
   I4 => W_32_31_i_4_n_0,
   O => W_32_31_i_8_n_0
);
W_32_31_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x96_out_13,
   I1 => x96_out_15,
   I2 => W_32_31_i_12_n_0,
   I3 => W_32_31_i_13_n_0,
   I4 => W_32_31_i_5_n_0,
   O => W_32_31_i_9_n_0
);
W_32_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x117_out_2,
   I1 => x106_out_2,
   I2 => x116_out_20,
   I3 => x116_out_9,
   I4 => x116_out_5,
   O => W_32_3_i_10_n_0
);
W_32_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x106_out_1,
   I1 => x116_out_4,
   I2 => x116_out_8,
   I3 => x116_out_19,
   I4 => x117_out_1,
   O => W_32_3_i_11_n_0
);
W_32_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x116_out_19,
   I1 => x116_out_8,
   I2 => x116_out_4,
   O => SIGMA_LCASE_0255_out_1
);
W_32_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x96_out_21,
   I1 => x96_out_19,
   I2 => x96_out_12,
   O => SIGMA_LCASE_1259_out_0_2
);
W_32_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x96_out_20,
   I1 => x96_out_18,
   I2 => x96_out_11,
   O => SIGMA_LCASE_1259_out_1
);
W_32_3_i_15 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x117_out_1,
   I1 => x106_out_1,
   I2 => x116_out_19,
   I3 => x116_out_8,
   I4 => x116_out_4,
   O => W_32_3_i_15_n_0
);
W_32_3_i_16 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x116_out_18,
   I1 => x116_out_7,
   I2 => x116_out_3,
   O => SIGMA_LCASE_0255_out_0
);
W_32_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x96_out_12,
   I1 => x96_out_19,
   I2 => x96_out_21,
   I3 => W_32_3_i_10_n_0,
   I4 => W_32_3_i_11_n_0,
   O => W_32_3_i_2_n_0
);
W_32_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_32_3_i_11_n_0,
   I1 => x96_out_21,
   I2 => x96_out_19,
   I3 => x96_out_12,
   I4 => W_32_3_i_10_n_0,
   O => W_32_3_i_3_n_0
);
W_32_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_0255_out_1,
   I1 => x106_out_1,
   I2 => x117_out_1,
   I3 => x96_out_11,
   I4 => x96_out_18,
   I5 => x96_out_20,
   O => W_32_3_i_4_n_0
);
W_32_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x117_out_0,
   I1 => x106_out_0,
   I2 => x116_out_18,
   I3 => x116_out_7,
   I4 => x116_out_3,
   O => W_32_3_i_5_n_0
);
W_32_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_32_3_i_2_n_0,
   I1 => W_32_7_i_16_n_0,
   I2 => x96_out_13,
   I3 => x96_out_20,
   I4 => x96_out_22,
   I5 => W_32_7_i_17_n_0,
   O => W_32_3_i_6_n_0
);
W_32_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_32_3_i_10_n_0,
   I1 => SIGMA_LCASE_1259_out_0_2,
   I2 => x117_out_1,
   I3 => x106_out_1,
   I4 => SIGMA_LCASE_0255_out_1,
   I5 => SIGMA_LCASE_1259_out_1,
   O => W_32_3_i_7_n_0
);
W_32_3_i_8 : LUT5
  generic map(
   INIT => X"99969666"
  )
 port map (
   I0 => SIGMA_LCASE_1259_out_1,
   I1 => W_32_3_i_15_n_0,
   I2 => x117_out_0,
   I3 => SIGMA_LCASE_0255_out_0,
   I4 => x106_out_0,
   O => W_32_3_i_8_n_0
);
W_32_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_32_3_i_5_n_0,
   I1 => x96_out_10,
   I2 => x96_out_17,
   I3 => x96_out_19,
   O => W_32_3_i_9_n_0
);
W_32_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x117_out_6,
   I1 => x106_out_6,
   I2 => x116_out_24,
   I3 => x116_out_13,
   I4 => x116_out_9,
   O => W_32_7_i_10_n_0
);
W_32_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x106_out_5,
   I1 => x116_out_8,
   I2 => x116_out_12,
   I3 => x116_out_23,
   I4 => x117_out_5,
   O => W_32_7_i_11_n_0
);
W_32_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x117_out_5,
   I1 => x106_out_5,
   I2 => x116_out_23,
   I3 => x116_out_12,
   I4 => x116_out_8,
   O => W_32_7_i_12_n_0
);
W_32_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x106_out_4,
   I1 => x116_out_7,
   I2 => x116_out_11,
   I3 => x116_out_22,
   I4 => x117_out_4,
   O => W_32_7_i_13_n_0
);
W_32_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x117_out_4,
   I1 => x106_out_4,
   I2 => x116_out_22,
   I3 => x116_out_11,
   I4 => x116_out_7,
   O => W_32_7_i_14_n_0
);
W_32_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x106_out_3,
   I1 => x116_out_6,
   I2 => x116_out_10,
   I3 => x116_out_21,
   I4 => x117_out_3,
   O => W_32_7_i_15_n_0
);
W_32_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x117_out_3,
   I1 => x106_out_3,
   I2 => x116_out_21,
   I3 => x116_out_10,
   I4 => x116_out_6,
   O => W_32_7_i_16_n_0
);
W_32_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x106_out_2,
   I1 => x116_out_5,
   I2 => x116_out_9,
   I3 => x116_out_20,
   I4 => x117_out_2,
   O => W_32_7_i_17_n_0
);
W_32_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x96_out_16,
   I1 => x96_out_23,
   I2 => x96_out_25,
   I3 => W_32_7_i_10_n_0,
   I4 => W_32_7_i_11_n_0,
   O => W_32_7_i_2_n_0
);
W_32_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x96_out_15,
   I1 => x96_out_22,
   I2 => x96_out_24,
   I3 => W_32_7_i_12_n_0,
   I4 => W_32_7_i_13_n_0,
   O => W_32_7_i_3_n_0
);
W_32_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x96_out_14,
   I1 => x96_out_21,
   I2 => x96_out_23,
   I3 => W_32_7_i_14_n_0,
   I4 => W_32_7_i_15_n_0,
   O => W_32_7_i_4_n_0
);
W_32_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x96_out_13,
   I1 => x96_out_20,
   I2 => x96_out_22,
   I3 => W_32_7_i_16_n_0,
   I4 => W_32_7_i_17_n_0,
   O => W_32_7_i_5_n_0
);
W_32_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_32_7_i_2_n_0,
   I1 => W_32_11_i_16_n_0,
   I2 => x96_out_17,
   I3 => x96_out_24,
   I4 => x96_out_26,
   I5 => W_32_11_i_17_n_0,
   O => W_32_7_i_6_n_0
);
W_32_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_32_7_i_3_n_0,
   I1 => W_32_7_i_10_n_0,
   I2 => x96_out_16,
   I3 => x96_out_23,
   I4 => x96_out_25,
   I5 => W_32_7_i_11_n_0,
   O => W_32_7_i_7_n_0
);
W_32_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_32_7_i_4_n_0,
   I1 => W_32_7_i_12_n_0,
   I2 => x96_out_15,
   I3 => x96_out_22,
   I4 => x96_out_24,
   I5 => W_32_7_i_13_n_0,
   O => W_32_7_i_8_n_0
);
W_32_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_32_7_i_5_n_0,
   I1 => W_32_7_i_14_n_0,
   I2 => x96_out_14,
   I3 => x96_out_21,
   I4 => x96_out_23,
   I5 => W_32_7_i_15_n_0,
   O => W_32_7_i_9_n_0
);
W_33_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x116_out_10,
   I1 => x104_out_10,
   I2 => x115_out_28,
   I3 => x115_out_17,
   I4 => x115_out_13,
   O => W_33_11_i_10_n_0
);
W_33_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x104_out_9,
   I1 => x115_out_12,
   I2 => x115_out_16,
   I3 => x115_out_27,
   I4 => x116_out_9,
   O => W_33_11_i_11_n_0
);
W_33_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x116_out_9,
   I1 => x104_out_9,
   I2 => x115_out_27,
   I3 => x115_out_16,
   I4 => x115_out_12,
   O => W_33_11_i_12_n_0
);
W_33_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x104_out_8,
   I1 => x115_out_11,
   I2 => x115_out_15,
   I3 => x115_out_26,
   I4 => x116_out_8,
   O => W_33_11_i_13_n_0
);
W_33_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x116_out_8,
   I1 => x104_out_8,
   I2 => x115_out_26,
   I3 => x115_out_15,
   I4 => x115_out_11,
   O => W_33_11_i_14_n_0
);
W_33_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x104_out_7,
   I1 => x115_out_10,
   I2 => x115_out_14,
   I3 => x115_out_25,
   I4 => x116_out_7,
   O => W_33_11_i_15_n_0
);
W_33_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x116_out_7,
   I1 => x104_out_7,
   I2 => x115_out_25,
   I3 => x115_out_14,
   I4 => x115_out_10,
   O => W_33_11_i_16_n_0
);
W_33_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x104_out_6,
   I1 => x115_out_9,
   I2 => x115_out_13,
   I3 => x115_out_24,
   I4 => x116_out_6,
   O => W_33_11_i_17_n_0
);
W_33_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x94_out_20,
   I1 => x94_out_27,
   I2 => x94_out_29,
   I3 => W_33_11_i_10_n_0,
   I4 => W_33_11_i_11_n_0,
   O => W_33_11_i_2_n_0
);
W_33_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x94_out_19,
   I1 => x94_out_26,
   I2 => x94_out_28,
   I3 => W_33_11_i_12_n_0,
   I4 => W_33_11_i_13_n_0,
   O => W_33_11_i_3_n_0
);
W_33_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x94_out_18,
   I1 => x94_out_25,
   I2 => x94_out_27,
   I3 => W_33_11_i_14_n_0,
   I4 => W_33_11_i_15_n_0,
   O => W_33_11_i_4_n_0
);
W_33_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x94_out_17,
   I1 => x94_out_24,
   I2 => x94_out_26,
   I3 => W_33_11_i_16_n_0,
   I4 => W_33_11_i_17_n_0,
   O => W_33_11_i_5_n_0
);
W_33_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_33_11_i_2_n_0,
   I1 => W_33_15_i_16_n_0,
   I2 => x94_out_21,
   I3 => x94_out_28,
   I4 => x94_out_30,
   I5 => W_33_15_i_17_n_0,
   O => W_33_11_i_6_n_0
);
W_33_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_33_11_i_3_n_0,
   I1 => W_33_11_i_10_n_0,
   I2 => x94_out_20,
   I3 => x94_out_27,
   I4 => x94_out_29,
   I5 => W_33_11_i_11_n_0,
   O => W_33_11_i_7_n_0
);
W_33_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_33_11_i_4_n_0,
   I1 => W_33_11_i_12_n_0,
   I2 => x94_out_19,
   I3 => x94_out_26,
   I4 => x94_out_28,
   I5 => W_33_11_i_13_n_0,
   O => W_33_11_i_8_n_0
);
W_33_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_33_11_i_5_n_0,
   I1 => W_33_11_i_14_n_0,
   I2 => x94_out_18,
   I3 => x94_out_25,
   I4 => x94_out_27,
   I5 => W_33_11_i_15_n_0,
   O => W_33_11_i_9_n_0
);
W_33_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x116_out_14,
   I1 => x104_out_14,
   I2 => x115_out_0,
   I3 => x115_out_21,
   I4 => x115_out_17,
   O => W_33_15_i_10_n_0
);
W_33_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x104_out_13,
   I1 => x115_out_16,
   I2 => x115_out_20,
   I3 => x115_out_31,
   I4 => x116_out_13,
   O => W_33_15_i_11_n_0
);
W_33_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x116_out_13,
   I1 => x104_out_13,
   I2 => x115_out_31,
   I3 => x115_out_20,
   I4 => x115_out_16,
   O => W_33_15_i_12_n_0
);
W_33_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x104_out_12,
   I1 => x115_out_15,
   I2 => x115_out_19,
   I3 => x115_out_30,
   I4 => x116_out_12,
   O => W_33_15_i_13_n_0
);
W_33_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x116_out_12,
   I1 => x104_out_12,
   I2 => x115_out_30,
   I3 => x115_out_19,
   I4 => x115_out_15,
   O => W_33_15_i_14_n_0
);
W_33_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x104_out_11,
   I1 => x115_out_14,
   I2 => x115_out_18,
   I3 => x115_out_29,
   I4 => x116_out_11,
   O => W_33_15_i_15_n_0
);
W_33_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x116_out_11,
   I1 => x104_out_11,
   I2 => x115_out_29,
   I3 => x115_out_18,
   I4 => x115_out_14,
   O => W_33_15_i_16_n_0
);
W_33_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x104_out_10,
   I1 => x115_out_13,
   I2 => x115_out_17,
   I3 => x115_out_28,
   I4 => x116_out_10,
   O => W_33_15_i_17_n_0
);
W_33_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x94_out_24,
   I1 => x94_out_31,
   I2 => x94_out_1,
   I3 => W_33_15_i_10_n_0,
   I4 => W_33_15_i_11_n_0,
   O => W_33_15_i_2_n_0
);
W_33_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x94_out_23,
   I1 => x94_out_30,
   I2 => x94_out_0,
   I3 => W_33_15_i_12_n_0,
   I4 => W_33_15_i_13_n_0,
   O => W_33_15_i_3_n_0
);
W_33_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x94_out_22,
   I1 => x94_out_29,
   I2 => x94_out_31,
   I3 => W_33_15_i_14_n_0,
   I4 => W_33_15_i_15_n_0,
   O => W_33_15_i_4_n_0
);
W_33_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x94_out_21,
   I1 => x94_out_28,
   I2 => x94_out_30,
   I3 => W_33_15_i_16_n_0,
   I4 => W_33_15_i_17_n_0,
   O => W_33_15_i_5_n_0
);
W_33_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_33_15_i_2_n_0,
   I1 => W_33_19_i_16_n_0,
   I2 => x94_out_25,
   I3 => x94_out_0,
   I4 => x94_out_2,
   I5 => W_33_19_i_17_n_0,
   O => W_33_15_i_6_n_0
);
W_33_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_33_15_i_3_n_0,
   I1 => W_33_15_i_10_n_0,
   I2 => x94_out_24,
   I3 => x94_out_31,
   I4 => x94_out_1,
   I5 => W_33_15_i_11_n_0,
   O => W_33_15_i_7_n_0
);
W_33_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_33_15_i_4_n_0,
   I1 => W_33_15_i_12_n_0,
   I2 => x94_out_23,
   I3 => x94_out_30,
   I4 => x94_out_0,
   I5 => W_33_15_i_13_n_0,
   O => W_33_15_i_8_n_0
);
W_33_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_33_15_i_5_n_0,
   I1 => W_33_15_i_14_n_0,
   I2 => x94_out_22,
   I3 => x94_out_29,
   I4 => x94_out_31,
   I5 => W_33_15_i_15_n_0,
   O => W_33_15_i_9_n_0
);
W_33_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x116_out_18,
   I1 => x104_out_18,
   I2 => x115_out_4,
   I3 => x115_out_25,
   I4 => x115_out_21,
   O => W_33_19_i_10_n_0
);
W_33_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x104_out_17,
   I1 => x115_out_20,
   I2 => x115_out_24,
   I3 => x115_out_3,
   I4 => x116_out_17,
   O => W_33_19_i_11_n_0
);
W_33_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x116_out_17,
   I1 => x104_out_17,
   I2 => x115_out_3,
   I3 => x115_out_24,
   I4 => x115_out_20,
   O => W_33_19_i_12_n_0
);
W_33_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x104_out_16,
   I1 => x115_out_19,
   I2 => x115_out_23,
   I3 => x115_out_2,
   I4 => x116_out_16,
   O => W_33_19_i_13_n_0
);
W_33_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x116_out_16,
   I1 => x104_out_16,
   I2 => x115_out_2,
   I3 => x115_out_23,
   I4 => x115_out_19,
   O => W_33_19_i_14_n_0
);
W_33_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x104_out_15,
   I1 => x115_out_18,
   I2 => x115_out_22,
   I3 => x115_out_1,
   I4 => x116_out_15,
   O => W_33_19_i_15_n_0
);
W_33_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x116_out_15,
   I1 => x104_out_15,
   I2 => x115_out_1,
   I3 => x115_out_22,
   I4 => x115_out_18,
   O => W_33_19_i_16_n_0
);
W_33_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x104_out_14,
   I1 => x115_out_17,
   I2 => x115_out_21,
   I3 => x115_out_0,
   I4 => x116_out_14,
   O => W_33_19_i_17_n_0
);
W_33_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x94_out_28,
   I1 => x94_out_3,
   I2 => x94_out_5,
   I3 => W_33_19_i_10_n_0,
   I4 => W_33_19_i_11_n_0,
   O => W_33_19_i_2_n_0
);
W_33_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x94_out_27,
   I1 => x94_out_2,
   I2 => x94_out_4,
   I3 => W_33_19_i_12_n_0,
   I4 => W_33_19_i_13_n_0,
   O => W_33_19_i_3_n_0
);
W_33_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x94_out_26,
   I1 => x94_out_1,
   I2 => x94_out_3,
   I3 => W_33_19_i_14_n_0,
   I4 => W_33_19_i_15_n_0,
   O => W_33_19_i_4_n_0
);
W_33_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x94_out_25,
   I1 => x94_out_0,
   I2 => x94_out_2,
   I3 => W_33_19_i_16_n_0,
   I4 => W_33_19_i_17_n_0,
   O => W_33_19_i_5_n_0
);
W_33_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_33_19_i_2_n_0,
   I1 => W_33_23_i_16_n_0,
   I2 => x94_out_29,
   I3 => x94_out_4,
   I4 => x94_out_6,
   I5 => W_33_23_i_17_n_0,
   O => W_33_19_i_6_n_0
);
W_33_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_33_19_i_3_n_0,
   I1 => W_33_19_i_10_n_0,
   I2 => x94_out_28,
   I3 => x94_out_3,
   I4 => x94_out_5,
   I5 => W_33_19_i_11_n_0,
   O => W_33_19_i_7_n_0
);
W_33_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_33_19_i_4_n_0,
   I1 => W_33_19_i_12_n_0,
   I2 => x94_out_27,
   I3 => x94_out_2,
   I4 => x94_out_4,
   I5 => W_33_19_i_13_n_0,
   O => W_33_19_i_8_n_0
);
W_33_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_33_19_i_5_n_0,
   I1 => W_33_19_i_14_n_0,
   I2 => x94_out_26,
   I3 => x94_out_1,
   I4 => x94_out_3,
   I5 => W_33_19_i_15_n_0,
   O => W_33_19_i_9_n_0
);
W_33_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x116_out_22,
   I1 => x104_out_22,
   I2 => x115_out_8,
   I3 => x115_out_29,
   I4 => x115_out_25,
   O => W_33_23_i_10_n_0
);
W_33_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x104_out_21,
   I1 => x115_out_24,
   I2 => x115_out_28,
   I3 => x115_out_7,
   I4 => x116_out_21,
   O => W_33_23_i_11_n_0
);
W_33_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x116_out_21,
   I1 => x104_out_21,
   I2 => x115_out_7,
   I3 => x115_out_28,
   I4 => x115_out_24,
   O => W_33_23_i_12_n_0
);
W_33_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x104_out_20,
   I1 => x115_out_23,
   I2 => x115_out_27,
   I3 => x115_out_6,
   I4 => x116_out_20,
   O => W_33_23_i_13_n_0
);
W_33_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x116_out_20,
   I1 => x104_out_20,
   I2 => x115_out_6,
   I3 => x115_out_27,
   I4 => x115_out_23,
   O => W_33_23_i_14_n_0
);
W_33_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x104_out_19,
   I1 => x115_out_22,
   I2 => x115_out_26,
   I3 => x115_out_5,
   I4 => x116_out_19,
   O => W_33_23_i_15_n_0
);
W_33_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x116_out_19,
   I1 => x104_out_19,
   I2 => x115_out_5,
   I3 => x115_out_26,
   I4 => x115_out_22,
   O => W_33_23_i_16_n_0
);
W_33_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x104_out_18,
   I1 => x115_out_21,
   I2 => x115_out_25,
   I3 => x115_out_4,
   I4 => x116_out_18,
   O => W_33_23_i_17_n_0
);
W_33_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x94_out_7,
   I1 => x94_out_9,
   I2 => W_33_23_i_10_n_0,
   I3 => W_33_23_i_11_n_0,
   O => W_33_23_i_2_n_0
);
W_33_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x94_out_31,
   I1 => x94_out_6,
   I2 => x94_out_8,
   I3 => W_33_23_i_12_n_0,
   I4 => W_33_23_i_13_n_0,
   O => W_33_23_i_3_n_0
);
W_33_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x94_out_30,
   I1 => x94_out_5,
   I2 => x94_out_7,
   I3 => W_33_23_i_14_n_0,
   I4 => W_33_23_i_15_n_0,
   O => W_33_23_i_4_n_0
);
W_33_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x94_out_29,
   I1 => x94_out_4,
   I2 => x94_out_6,
   I3 => W_33_23_i_16_n_0,
   I4 => W_33_23_i_17_n_0,
   O => W_33_23_i_5_n_0
);
W_33_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x94_out_8,
   I1 => x94_out_10,
   I2 => W_33_27_i_16_n_0,
   I3 => W_33_27_i_17_n_0,
   I4 => W_33_23_i_2_n_0,
   O => W_33_23_i_6_n_0
);
W_33_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x94_out_7,
   I1 => x94_out_9,
   I2 => W_33_23_i_10_n_0,
   I3 => W_33_23_i_11_n_0,
   I4 => W_33_23_i_3_n_0,
   O => W_33_23_i_7_n_0
);
W_33_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_33_23_i_4_n_0,
   I1 => W_33_23_i_12_n_0,
   I2 => x94_out_31,
   I3 => x94_out_6,
   I4 => x94_out_8,
   I5 => W_33_23_i_13_n_0,
   O => W_33_23_i_8_n_0
);
W_33_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_33_23_i_5_n_0,
   I1 => W_33_23_i_14_n_0,
   I2 => x94_out_30,
   I3 => x94_out_5,
   I4 => x94_out_7,
   I5 => W_33_23_i_15_n_0,
   O => W_33_23_i_9_n_0
);
W_33_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x116_out_26,
   I1 => x104_out_26,
   I2 => x115_out_12,
   I3 => x115_out_1,
   I4 => x115_out_29,
   O => W_33_27_i_10_n_0
);
W_33_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x104_out_25,
   I1 => x115_out_28,
   I2 => x115_out_0,
   I3 => x115_out_11,
   I4 => x116_out_25,
   O => W_33_27_i_11_n_0
);
W_33_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x116_out_25,
   I1 => x104_out_25,
   I2 => x115_out_11,
   I3 => x115_out_0,
   I4 => x115_out_28,
   O => W_33_27_i_12_n_0
);
W_33_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x104_out_24,
   I1 => x115_out_27,
   I2 => x115_out_31,
   I3 => x115_out_10,
   I4 => x116_out_24,
   O => W_33_27_i_13_n_0
);
W_33_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x116_out_24,
   I1 => x104_out_24,
   I2 => x115_out_10,
   I3 => x115_out_31,
   I4 => x115_out_27,
   O => W_33_27_i_14_n_0
);
W_33_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x104_out_23,
   I1 => x115_out_26,
   I2 => x115_out_30,
   I3 => x115_out_9,
   I4 => x116_out_23,
   O => W_33_27_i_15_n_0
);
W_33_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x116_out_23,
   I1 => x104_out_23,
   I2 => x115_out_9,
   I3 => x115_out_30,
   I4 => x115_out_26,
   O => W_33_27_i_16_n_0
);
W_33_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x104_out_22,
   I1 => x115_out_25,
   I2 => x115_out_29,
   I3 => x115_out_8,
   I4 => x116_out_22,
   O => W_33_27_i_17_n_0
);
W_33_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x94_out_11,
   I1 => x94_out_13,
   I2 => W_33_27_i_10_n_0,
   I3 => W_33_27_i_11_n_0,
   O => W_33_27_i_2_n_0
);
W_33_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x94_out_10,
   I1 => x94_out_12,
   I2 => W_33_27_i_12_n_0,
   I3 => W_33_27_i_13_n_0,
   O => W_33_27_i_3_n_0
);
W_33_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x94_out_9,
   I1 => x94_out_11,
   I2 => W_33_27_i_14_n_0,
   I3 => W_33_27_i_15_n_0,
   O => W_33_27_i_4_n_0
);
W_33_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x94_out_8,
   I1 => x94_out_10,
   I2 => W_33_27_i_16_n_0,
   I3 => W_33_27_i_17_n_0,
   O => W_33_27_i_5_n_0
);
W_33_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x94_out_12,
   I1 => x94_out_14,
   I2 => W_33_31_i_13_n_0,
   I3 => W_33_31_i_14_n_0,
   I4 => W_33_27_i_2_n_0,
   O => W_33_27_i_6_n_0
);
W_33_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x94_out_11,
   I1 => x94_out_13,
   I2 => W_33_27_i_10_n_0,
   I3 => W_33_27_i_11_n_0,
   I4 => W_33_27_i_3_n_0,
   O => W_33_27_i_7_n_0
);
W_33_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x94_out_10,
   I1 => x94_out_12,
   I2 => W_33_27_i_12_n_0,
   I3 => W_33_27_i_13_n_0,
   I4 => W_33_27_i_4_n_0,
   O => W_33_27_i_8_n_0
);
W_33_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x94_out_9,
   I1 => x94_out_11,
   I2 => W_33_27_i_14_n_0,
   I3 => W_33_27_i_15_n_0,
   I4 => W_33_27_i_5_n_0,
   O => W_33_27_i_9_n_0
);
W_33_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x104_out_28,
   I1 => x115_out_31,
   I2 => x115_out_3,
   I3 => x115_out_14,
   I4 => x116_out_28,
   O => W_33_31_i_10_n_0
);
W_33_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x116_out_28,
   I1 => x104_out_28,
   I2 => x115_out_14,
   I3 => x115_out_3,
   I4 => x115_out_31,
   O => W_33_31_i_11_n_0
);
W_33_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x104_out_27,
   I1 => x115_out_30,
   I2 => x115_out_2,
   I3 => x115_out_13,
   I4 => x116_out_27,
   O => W_33_31_i_12_n_0
);
W_33_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x116_out_27,
   I1 => x104_out_27,
   I2 => x115_out_13,
   I3 => x115_out_2,
   I4 => x115_out_30,
   O => W_33_31_i_13_n_0
);
W_33_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x104_out_26,
   I1 => x115_out_29,
   I2 => x115_out_1,
   I3 => x115_out_12,
   I4 => x116_out_26,
   O => W_33_31_i_14_n_0
);
W_33_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x104_out_29,
   I1 => x115_out_4,
   I2 => x115_out_15,
   I3 => x116_out_29,
   O => W_33_31_i_15_n_0
);
W_33_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x94_out_17,
   I1 => x94_out_15,
   O => SIGMA_LCASE_1251_out_0_30
);
W_33_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => x115_out_6,
   I1 => x115_out_17,
   I2 => x104_out_31,
   I3 => x116_out_31,
   I4 => x94_out_16,
   I5 => x94_out_18,
   O => W_33_31_i_17_n_0
);
W_33_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x115_out_16,
   I1 => x115_out_5,
   O => SIGMA_LCASE_0247_out_30
);
W_33_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x116_out_30,
   I1 => x104_out_30,
   I2 => x115_out_16,
   I3 => x115_out_5,
   O => W_33_31_i_19_n_0
);
W_33_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x94_out_14,
   I1 => x94_out_16,
   I2 => W_33_31_i_9_n_0,
   I3 => W_33_31_i_10_n_0,
   O => W_33_31_i_2_n_0
);
W_33_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x94_out_13,
   I1 => x94_out_15,
   I2 => W_33_31_i_11_n_0,
   I3 => W_33_31_i_12_n_0,
   O => W_33_31_i_3_n_0
);
W_33_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x94_out_12,
   I1 => x94_out_14,
   I2 => W_33_31_i_13_n_0,
   I3 => W_33_31_i_14_n_0,
   O => W_33_31_i_4_n_0
);
W_33_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_33_31_i_15_n_0,
   I1 => SIGMA_LCASE_1251_out_0_30,
   I2 => W_33_31_i_17_n_0,
   I3 => x104_out_30,
   I4 => SIGMA_LCASE_0247_out_30,
   I5 => x116_out_30,
   O => W_33_31_i_5_n_0
);
W_33_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_33_31_i_2_n_0,
   I1 => W_33_31_i_19_n_0,
   I2 => x94_out_15,
   I3 => x94_out_17,
   I4 => W_33_31_i_15_n_0,
   O => W_33_31_i_6_n_0
);
W_33_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x94_out_14,
   I1 => x94_out_16,
   I2 => W_33_31_i_9_n_0,
   I3 => W_33_31_i_10_n_0,
   I4 => W_33_31_i_3_n_0,
   O => W_33_31_i_7_n_0
);
W_33_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x94_out_13,
   I1 => x94_out_15,
   I2 => W_33_31_i_11_n_0,
   I3 => W_33_31_i_12_n_0,
   I4 => W_33_31_i_4_n_0,
   O => W_33_31_i_8_n_0
);
W_33_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x116_out_29,
   I1 => x104_out_29,
   I2 => x115_out_15,
   I3 => x115_out_4,
   O => W_33_31_i_9_n_0
);
W_33_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x116_out_2,
   I1 => x104_out_2,
   I2 => x115_out_20,
   I3 => x115_out_9,
   I4 => x115_out_5,
   O => W_33_3_i_10_n_0
);
W_33_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x104_out_1,
   I1 => x115_out_4,
   I2 => x115_out_8,
   I3 => x115_out_19,
   I4 => x116_out_1,
   O => W_33_3_i_11_n_0
);
W_33_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x115_out_19,
   I1 => x115_out_8,
   I2 => x115_out_4,
   O => SIGMA_LCASE_0247_out_1
);
W_33_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x94_out_21,
   I1 => x94_out_19,
   I2 => x94_out_12,
   O => SIGMA_LCASE_1251_out_0_2
);
W_33_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x94_out_20,
   I1 => x94_out_18,
   I2 => x94_out_11,
   O => SIGMA_LCASE_1251_out_1
);
W_33_3_i_15 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x116_out_1,
   I1 => x104_out_1,
   I2 => x115_out_19,
   I3 => x115_out_8,
   I4 => x115_out_4,
   O => W_33_3_i_15_n_0
);
W_33_3_i_16 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x115_out_18,
   I1 => x115_out_7,
   I2 => x115_out_3,
   O => SIGMA_LCASE_0247_out_0
);
W_33_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x94_out_12,
   I1 => x94_out_19,
   I2 => x94_out_21,
   I3 => W_33_3_i_10_n_0,
   I4 => W_33_3_i_11_n_0,
   O => W_33_3_i_2_n_0
);
W_33_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_33_3_i_11_n_0,
   I1 => x94_out_21,
   I2 => x94_out_19,
   I3 => x94_out_12,
   I4 => W_33_3_i_10_n_0,
   O => W_33_3_i_3_n_0
);
W_33_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_0247_out_1,
   I1 => x104_out_1,
   I2 => x116_out_1,
   I3 => x94_out_11,
   I4 => x94_out_18,
   I5 => x94_out_20,
   O => W_33_3_i_4_n_0
);
W_33_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x116_out_0,
   I1 => x104_out_0,
   I2 => x115_out_18,
   I3 => x115_out_7,
   I4 => x115_out_3,
   O => W_33_3_i_5_n_0
);
W_33_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_33_3_i_2_n_0,
   I1 => W_33_7_i_16_n_0,
   I2 => x94_out_13,
   I3 => x94_out_20,
   I4 => x94_out_22,
   I5 => W_33_7_i_17_n_0,
   O => W_33_3_i_6_n_0
);
W_33_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_33_3_i_10_n_0,
   I1 => SIGMA_LCASE_1251_out_0_2,
   I2 => x116_out_1,
   I3 => x104_out_1,
   I4 => SIGMA_LCASE_0247_out_1,
   I5 => SIGMA_LCASE_1251_out_1,
   O => W_33_3_i_7_n_0
);
W_33_3_i_8 : LUT5
  generic map(
   INIT => X"99969666"
  )
 port map (
   I0 => SIGMA_LCASE_1251_out_1,
   I1 => W_33_3_i_15_n_0,
   I2 => x116_out_0,
   I3 => SIGMA_LCASE_0247_out_0,
   I4 => x104_out_0,
   O => W_33_3_i_8_n_0
);
W_33_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_33_3_i_5_n_0,
   I1 => x94_out_10,
   I2 => x94_out_17,
   I3 => x94_out_19,
   O => W_33_3_i_9_n_0
);
W_33_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x116_out_6,
   I1 => x104_out_6,
   I2 => x115_out_24,
   I3 => x115_out_13,
   I4 => x115_out_9,
   O => W_33_7_i_10_n_0
);
W_33_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x104_out_5,
   I1 => x115_out_8,
   I2 => x115_out_12,
   I3 => x115_out_23,
   I4 => x116_out_5,
   O => W_33_7_i_11_n_0
);
W_33_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x116_out_5,
   I1 => x104_out_5,
   I2 => x115_out_23,
   I3 => x115_out_12,
   I4 => x115_out_8,
   O => W_33_7_i_12_n_0
);
W_33_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x104_out_4,
   I1 => x115_out_7,
   I2 => x115_out_11,
   I3 => x115_out_22,
   I4 => x116_out_4,
   O => W_33_7_i_13_n_0
);
W_33_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x116_out_4,
   I1 => x104_out_4,
   I2 => x115_out_22,
   I3 => x115_out_11,
   I4 => x115_out_7,
   O => W_33_7_i_14_n_0
);
W_33_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x104_out_3,
   I1 => x115_out_6,
   I2 => x115_out_10,
   I3 => x115_out_21,
   I4 => x116_out_3,
   O => W_33_7_i_15_n_0
);
W_33_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x116_out_3,
   I1 => x104_out_3,
   I2 => x115_out_21,
   I3 => x115_out_10,
   I4 => x115_out_6,
   O => W_33_7_i_16_n_0
);
W_33_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x104_out_2,
   I1 => x115_out_5,
   I2 => x115_out_9,
   I3 => x115_out_20,
   I4 => x116_out_2,
   O => W_33_7_i_17_n_0
);
W_33_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x94_out_16,
   I1 => x94_out_23,
   I2 => x94_out_25,
   I3 => W_33_7_i_10_n_0,
   I4 => W_33_7_i_11_n_0,
   O => W_33_7_i_2_n_0
);
W_33_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x94_out_15,
   I1 => x94_out_22,
   I2 => x94_out_24,
   I3 => W_33_7_i_12_n_0,
   I4 => W_33_7_i_13_n_0,
   O => W_33_7_i_3_n_0
);
W_33_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x94_out_14,
   I1 => x94_out_21,
   I2 => x94_out_23,
   I3 => W_33_7_i_14_n_0,
   I4 => W_33_7_i_15_n_0,
   O => W_33_7_i_4_n_0
);
W_33_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x94_out_13,
   I1 => x94_out_20,
   I2 => x94_out_22,
   I3 => W_33_7_i_16_n_0,
   I4 => W_33_7_i_17_n_0,
   O => W_33_7_i_5_n_0
);
W_33_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_33_7_i_2_n_0,
   I1 => W_33_11_i_16_n_0,
   I2 => x94_out_17,
   I3 => x94_out_24,
   I4 => x94_out_26,
   I5 => W_33_11_i_17_n_0,
   O => W_33_7_i_6_n_0
);
W_33_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_33_7_i_3_n_0,
   I1 => W_33_7_i_10_n_0,
   I2 => x94_out_16,
   I3 => x94_out_23,
   I4 => x94_out_25,
   I5 => W_33_7_i_11_n_0,
   O => W_33_7_i_7_n_0
);
W_33_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_33_7_i_4_n_0,
   I1 => W_33_7_i_12_n_0,
   I2 => x94_out_15,
   I3 => x94_out_22,
   I4 => x94_out_24,
   I5 => W_33_7_i_13_n_0,
   O => W_33_7_i_8_n_0
);
W_33_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_33_7_i_5_n_0,
   I1 => W_33_7_i_14_n_0,
   I2 => x94_out_14,
   I3 => x94_out_21,
   I4 => x94_out_23,
   I5 => W_33_7_i_15_n_0,
   O => W_33_7_i_9_n_0
);
W_34_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x115_out_10,
   I1 => x102_out_10,
   I2 => x114_out_28,
   I3 => x114_out_17,
   I4 => x114_out_13,
   O => W_34_11_i_10_n_0
);
W_34_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x102_out_9,
   I1 => x114_out_12,
   I2 => x114_out_16,
   I3 => x114_out_27,
   I4 => x115_out_9,
   O => W_34_11_i_11_n_0
);
W_34_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x115_out_9,
   I1 => x102_out_9,
   I2 => x114_out_27,
   I3 => x114_out_16,
   I4 => x114_out_12,
   O => W_34_11_i_12_n_0
);
W_34_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x102_out_8,
   I1 => x114_out_11,
   I2 => x114_out_15,
   I3 => x114_out_26,
   I4 => x115_out_8,
   O => W_34_11_i_13_n_0
);
W_34_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x115_out_8,
   I1 => x102_out_8,
   I2 => x114_out_26,
   I3 => x114_out_15,
   I4 => x114_out_11,
   O => W_34_11_i_14_n_0
);
W_34_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x102_out_7,
   I1 => x114_out_10,
   I2 => x114_out_14,
   I3 => x114_out_25,
   I4 => x115_out_7,
   O => W_34_11_i_15_n_0
);
W_34_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x115_out_7,
   I1 => x102_out_7,
   I2 => x114_out_25,
   I3 => x114_out_14,
   I4 => x114_out_10,
   O => W_34_11_i_16_n_0
);
W_34_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x102_out_6,
   I1 => x114_out_9,
   I2 => x114_out_13,
   I3 => x114_out_24,
   I4 => x115_out_6,
   O => W_34_11_i_17_n_0
);
W_34_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x92_out_20,
   I1 => x92_out_27,
   I2 => x92_out_29,
   I3 => W_34_11_i_10_n_0,
   I4 => W_34_11_i_11_n_0,
   O => W_34_11_i_2_n_0
);
W_34_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x92_out_19,
   I1 => x92_out_26,
   I2 => x92_out_28,
   I3 => W_34_11_i_12_n_0,
   I4 => W_34_11_i_13_n_0,
   O => W_34_11_i_3_n_0
);
W_34_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x92_out_18,
   I1 => x92_out_25,
   I2 => x92_out_27,
   I3 => W_34_11_i_14_n_0,
   I4 => W_34_11_i_15_n_0,
   O => W_34_11_i_4_n_0
);
W_34_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x92_out_17,
   I1 => x92_out_24,
   I2 => x92_out_26,
   I3 => W_34_11_i_16_n_0,
   I4 => W_34_11_i_17_n_0,
   O => W_34_11_i_5_n_0
);
W_34_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_34_11_i_2_n_0,
   I1 => W_34_15_i_16_n_0,
   I2 => x92_out_21,
   I3 => x92_out_28,
   I4 => x92_out_30,
   I5 => W_34_15_i_17_n_0,
   O => W_34_11_i_6_n_0
);
W_34_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_34_11_i_3_n_0,
   I1 => W_34_11_i_10_n_0,
   I2 => x92_out_20,
   I3 => x92_out_27,
   I4 => x92_out_29,
   I5 => W_34_11_i_11_n_0,
   O => W_34_11_i_7_n_0
);
W_34_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_34_11_i_4_n_0,
   I1 => W_34_11_i_12_n_0,
   I2 => x92_out_19,
   I3 => x92_out_26,
   I4 => x92_out_28,
   I5 => W_34_11_i_13_n_0,
   O => W_34_11_i_8_n_0
);
W_34_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_34_11_i_5_n_0,
   I1 => W_34_11_i_14_n_0,
   I2 => x92_out_18,
   I3 => x92_out_25,
   I4 => x92_out_27,
   I5 => W_34_11_i_15_n_0,
   O => W_34_11_i_9_n_0
);
W_34_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x115_out_14,
   I1 => x102_out_14,
   I2 => x114_out_0,
   I3 => x114_out_21,
   I4 => x114_out_17,
   O => W_34_15_i_10_n_0
);
W_34_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x102_out_13,
   I1 => x114_out_16,
   I2 => x114_out_20,
   I3 => x114_out_31,
   I4 => x115_out_13,
   O => W_34_15_i_11_n_0
);
W_34_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x115_out_13,
   I1 => x102_out_13,
   I2 => x114_out_31,
   I3 => x114_out_20,
   I4 => x114_out_16,
   O => W_34_15_i_12_n_0
);
W_34_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x102_out_12,
   I1 => x114_out_15,
   I2 => x114_out_19,
   I3 => x114_out_30,
   I4 => x115_out_12,
   O => W_34_15_i_13_n_0
);
W_34_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x115_out_12,
   I1 => x102_out_12,
   I2 => x114_out_30,
   I3 => x114_out_19,
   I4 => x114_out_15,
   O => W_34_15_i_14_n_0
);
W_34_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x102_out_11,
   I1 => x114_out_14,
   I2 => x114_out_18,
   I3 => x114_out_29,
   I4 => x115_out_11,
   O => W_34_15_i_15_n_0
);
W_34_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x115_out_11,
   I1 => x102_out_11,
   I2 => x114_out_29,
   I3 => x114_out_18,
   I4 => x114_out_14,
   O => W_34_15_i_16_n_0
);
W_34_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x102_out_10,
   I1 => x114_out_13,
   I2 => x114_out_17,
   I3 => x114_out_28,
   I4 => x115_out_10,
   O => W_34_15_i_17_n_0
);
W_34_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x92_out_24,
   I1 => x92_out_31,
   I2 => x92_out_1,
   I3 => W_34_15_i_10_n_0,
   I4 => W_34_15_i_11_n_0,
   O => W_34_15_i_2_n_0
);
W_34_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x92_out_23,
   I1 => x92_out_30,
   I2 => x92_out_0,
   I3 => W_34_15_i_12_n_0,
   I4 => W_34_15_i_13_n_0,
   O => W_34_15_i_3_n_0
);
W_34_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x92_out_22,
   I1 => x92_out_29,
   I2 => x92_out_31,
   I3 => W_34_15_i_14_n_0,
   I4 => W_34_15_i_15_n_0,
   O => W_34_15_i_4_n_0
);
W_34_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x92_out_21,
   I1 => x92_out_28,
   I2 => x92_out_30,
   I3 => W_34_15_i_16_n_0,
   I4 => W_34_15_i_17_n_0,
   O => W_34_15_i_5_n_0
);
W_34_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_34_15_i_2_n_0,
   I1 => W_34_19_i_16_n_0,
   I2 => x92_out_25,
   I3 => x92_out_0,
   I4 => x92_out_2,
   I5 => W_34_19_i_17_n_0,
   O => W_34_15_i_6_n_0
);
W_34_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_34_15_i_3_n_0,
   I1 => W_34_15_i_10_n_0,
   I2 => x92_out_24,
   I3 => x92_out_31,
   I4 => x92_out_1,
   I5 => W_34_15_i_11_n_0,
   O => W_34_15_i_7_n_0
);
W_34_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_34_15_i_4_n_0,
   I1 => W_34_15_i_12_n_0,
   I2 => x92_out_23,
   I3 => x92_out_30,
   I4 => x92_out_0,
   I5 => W_34_15_i_13_n_0,
   O => W_34_15_i_8_n_0
);
W_34_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_34_15_i_5_n_0,
   I1 => W_34_15_i_14_n_0,
   I2 => x92_out_22,
   I3 => x92_out_29,
   I4 => x92_out_31,
   I5 => W_34_15_i_15_n_0,
   O => W_34_15_i_9_n_0
);
W_34_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x115_out_18,
   I1 => x102_out_18,
   I2 => x114_out_4,
   I3 => x114_out_25,
   I4 => x114_out_21,
   O => W_34_19_i_10_n_0
);
W_34_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x102_out_17,
   I1 => x114_out_20,
   I2 => x114_out_24,
   I3 => x114_out_3,
   I4 => x115_out_17,
   O => W_34_19_i_11_n_0
);
W_34_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x115_out_17,
   I1 => x102_out_17,
   I2 => x114_out_3,
   I3 => x114_out_24,
   I4 => x114_out_20,
   O => W_34_19_i_12_n_0
);
W_34_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x102_out_16,
   I1 => x114_out_19,
   I2 => x114_out_23,
   I3 => x114_out_2,
   I4 => x115_out_16,
   O => W_34_19_i_13_n_0
);
W_34_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x115_out_16,
   I1 => x102_out_16,
   I2 => x114_out_2,
   I3 => x114_out_23,
   I4 => x114_out_19,
   O => W_34_19_i_14_n_0
);
W_34_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x102_out_15,
   I1 => x114_out_18,
   I2 => x114_out_22,
   I3 => x114_out_1,
   I4 => x115_out_15,
   O => W_34_19_i_15_n_0
);
W_34_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x115_out_15,
   I1 => x102_out_15,
   I2 => x114_out_1,
   I3 => x114_out_22,
   I4 => x114_out_18,
   O => W_34_19_i_16_n_0
);
W_34_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x102_out_14,
   I1 => x114_out_17,
   I2 => x114_out_21,
   I3 => x114_out_0,
   I4 => x115_out_14,
   O => W_34_19_i_17_n_0
);
W_34_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x92_out_28,
   I1 => x92_out_3,
   I2 => x92_out_5,
   I3 => W_34_19_i_10_n_0,
   I4 => W_34_19_i_11_n_0,
   O => W_34_19_i_2_n_0
);
W_34_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x92_out_27,
   I1 => x92_out_2,
   I2 => x92_out_4,
   I3 => W_34_19_i_12_n_0,
   I4 => W_34_19_i_13_n_0,
   O => W_34_19_i_3_n_0
);
W_34_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x92_out_26,
   I1 => x92_out_1,
   I2 => x92_out_3,
   I3 => W_34_19_i_14_n_0,
   I4 => W_34_19_i_15_n_0,
   O => W_34_19_i_4_n_0
);
W_34_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x92_out_25,
   I1 => x92_out_0,
   I2 => x92_out_2,
   I3 => W_34_19_i_16_n_0,
   I4 => W_34_19_i_17_n_0,
   O => W_34_19_i_5_n_0
);
W_34_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_34_19_i_2_n_0,
   I1 => W_34_23_i_16_n_0,
   I2 => x92_out_29,
   I3 => x92_out_4,
   I4 => x92_out_6,
   I5 => W_34_23_i_17_n_0,
   O => W_34_19_i_6_n_0
);
W_34_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_34_19_i_3_n_0,
   I1 => W_34_19_i_10_n_0,
   I2 => x92_out_28,
   I3 => x92_out_3,
   I4 => x92_out_5,
   I5 => W_34_19_i_11_n_0,
   O => W_34_19_i_7_n_0
);
W_34_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_34_19_i_4_n_0,
   I1 => W_34_19_i_12_n_0,
   I2 => x92_out_27,
   I3 => x92_out_2,
   I4 => x92_out_4,
   I5 => W_34_19_i_13_n_0,
   O => W_34_19_i_8_n_0
);
W_34_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_34_19_i_5_n_0,
   I1 => W_34_19_i_14_n_0,
   I2 => x92_out_26,
   I3 => x92_out_1,
   I4 => x92_out_3,
   I5 => W_34_19_i_15_n_0,
   O => W_34_19_i_9_n_0
);
W_34_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x115_out_22,
   I1 => x102_out_22,
   I2 => x114_out_8,
   I3 => x114_out_29,
   I4 => x114_out_25,
   O => W_34_23_i_10_n_0
);
W_34_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x102_out_21,
   I1 => x114_out_24,
   I2 => x114_out_28,
   I3 => x114_out_7,
   I4 => x115_out_21,
   O => W_34_23_i_11_n_0
);
W_34_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x115_out_21,
   I1 => x102_out_21,
   I2 => x114_out_7,
   I3 => x114_out_28,
   I4 => x114_out_24,
   O => W_34_23_i_12_n_0
);
W_34_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x102_out_20,
   I1 => x114_out_23,
   I2 => x114_out_27,
   I3 => x114_out_6,
   I4 => x115_out_20,
   O => W_34_23_i_13_n_0
);
W_34_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x115_out_20,
   I1 => x102_out_20,
   I2 => x114_out_6,
   I3 => x114_out_27,
   I4 => x114_out_23,
   O => W_34_23_i_14_n_0
);
W_34_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x102_out_19,
   I1 => x114_out_22,
   I2 => x114_out_26,
   I3 => x114_out_5,
   I4 => x115_out_19,
   O => W_34_23_i_15_n_0
);
W_34_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x115_out_19,
   I1 => x102_out_19,
   I2 => x114_out_5,
   I3 => x114_out_26,
   I4 => x114_out_22,
   O => W_34_23_i_16_n_0
);
W_34_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x102_out_18,
   I1 => x114_out_21,
   I2 => x114_out_25,
   I3 => x114_out_4,
   I4 => x115_out_18,
   O => W_34_23_i_17_n_0
);
W_34_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x92_out_7,
   I1 => x92_out_9,
   I2 => W_34_23_i_10_n_0,
   I3 => W_34_23_i_11_n_0,
   O => W_34_23_i_2_n_0
);
W_34_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x92_out_31,
   I1 => x92_out_6,
   I2 => x92_out_8,
   I3 => W_34_23_i_12_n_0,
   I4 => W_34_23_i_13_n_0,
   O => W_34_23_i_3_n_0
);
W_34_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x92_out_30,
   I1 => x92_out_5,
   I2 => x92_out_7,
   I3 => W_34_23_i_14_n_0,
   I4 => W_34_23_i_15_n_0,
   O => W_34_23_i_4_n_0
);
W_34_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x92_out_29,
   I1 => x92_out_4,
   I2 => x92_out_6,
   I3 => W_34_23_i_16_n_0,
   I4 => W_34_23_i_17_n_0,
   O => W_34_23_i_5_n_0
);
W_34_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x92_out_8,
   I1 => x92_out_10,
   I2 => W_34_27_i_16_n_0,
   I3 => W_34_27_i_17_n_0,
   I4 => W_34_23_i_2_n_0,
   O => W_34_23_i_6_n_0
);
W_34_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x92_out_7,
   I1 => x92_out_9,
   I2 => W_34_23_i_10_n_0,
   I3 => W_34_23_i_11_n_0,
   I4 => W_34_23_i_3_n_0,
   O => W_34_23_i_7_n_0
);
W_34_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_34_23_i_4_n_0,
   I1 => W_34_23_i_12_n_0,
   I2 => x92_out_31,
   I3 => x92_out_6,
   I4 => x92_out_8,
   I5 => W_34_23_i_13_n_0,
   O => W_34_23_i_8_n_0
);
W_34_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_34_23_i_5_n_0,
   I1 => W_34_23_i_14_n_0,
   I2 => x92_out_30,
   I3 => x92_out_5,
   I4 => x92_out_7,
   I5 => W_34_23_i_15_n_0,
   O => W_34_23_i_9_n_0
);
W_34_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x115_out_26,
   I1 => x102_out_26,
   I2 => x114_out_12,
   I3 => x114_out_1,
   I4 => x114_out_29,
   O => W_34_27_i_10_n_0
);
W_34_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x102_out_25,
   I1 => x114_out_28,
   I2 => x114_out_0,
   I3 => x114_out_11,
   I4 => x115_out_25,
   O => W_34_27_i_11_n_0
);
W_34_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x115_out_25,
   I1 => x102_out_25,
   I2 => x114_out_11,
   I3 => x114_out_0,
   I4 => x114_out_28,
   O => W_34_27_i_12_n_0
);
W_34_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x102_out_24,
   I1 => x114_out_27,
   I2 => x114_out_31,
   I3 => x114_out_10,
   I4 => x115_out_24,
   O => W_34_27_i_13_n_0
);
W_34_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x115_out_24,
   I1 => x102_out_24,
   I2 => x114_out_10,
   I3 => x114_out_31,
   I4 => x114_out_27,
   O => W_34_27_i_14_n_0
);
W_34_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x102_out_23,
   I1 => x114_out_26,
   I2 => x114_out_30,
   I3 => x114_out_9,
   I4 => x115_out_23,
   O => W_34_27_i_15_n_0
);
W_34_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x115_out_23,
   I1 => x102_out_23,
   I2 => x114_out_9,
   I3 => x114_out_30,
   I4 => x114_out_26,
   O => W_34_27_i_16_n_0
);
W_34_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x102_out_22,
   I1 => x114_out_25,
   I2 => x114_out_29,
   I3 => x114_out_8,
   I4 => x115_out_22,
   O => W_34_27_i_17_n_0
);
W_34_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x92_out_11,
   I1 => x92_out_13,
   I2 => W_34_27_i_10_n_0,
   I3 => W_34_27_i_11_n_0,
   O => W_34_27_i_2_n_0
);
W_34_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x92_out_10,
   I1 => x92_out_12,
   I2 => W_34_27_i_12_n_0,
   I3 => W_34_27_i_13_n_0,
   O => W_34_27_i_3_n_0
);
W_34_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x92_out_9,
   I1 => x92_out_11,
   I2 => W_34_27_i_14_n_0,
   I3 => W_34_27_i_15_n_0,
   O => W_34_27_i_4_n_0
);
W_34_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x92_out_8,
   I1 => x92_out_10,
   I2 => W_34_27_i_16_n_0,
   I3 => W_34_27_i_17_n_0,
   O => W_34_27_i_5_n_0
);
W_34_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x92_out_12,
   I1 => x92_out_14,
   I2 => W_34_31_i_13_n_0,
   I3 => W_34_31_i_14_n_0,
   I4 => W_34_27_i_2_n_0,
   O => W_34_27_i_6_n_0
);
W_34_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x92_out_11,
   I1 => x92_out_13,
   I2 => W_34_27_i_10_n_0,
   I3 => W_34_27_i_11_n_0,
   I4 => W_34_27_i_3_n_0,
   O => W_34_27_i_7_n_0
);
W_34_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x92_out_10,
   I1 => x92_out_12,
   I2 => W_34_27_i_12_n_0,
   I3 => W_34_27_i_13_n_0,
   I4 => W_34_27_i_4_n_0,
   O => W_34_27_i_8_n_0
);
W_34_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x92_out_9,
   I1 => x92_out_11,
   I2 => W_34_27_i_14_n_0,
   I3 => W_34_27_i_15_n_0,
   I4 => W_34_27_i_5_n_0,
   O => W_34_27_i_9_n_0
);
W_34_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x102_out_28,
   I1 => x114_out_31,
   I2 => x114_out_3,
   I3 => x114_out_14,
   I4 => x115_out_28,
   O => W_34_31_i_10_n_0
);
W_34_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x115_out_28,
   I1 => x102_out_28,
   I2 => x114_out_14,
   I3 => x114_out_3,
   I4 => x114_out_31,
   O => W_34_31_i_11_n_0
);
W_34_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x102_out_27,
   I1 => x114_out_30,
   I2 => x114_out_2,
   I3 => x114_out_13,
   I4 => x115_out_27,
   O => W_34_31_i_12_n_0
);
W_34_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x115_out_27,
   I1 => x102_out_27,
   I2 => x114_out_13,
   I3 => x114_out_2,
   I4 => x114_out_30,
   O => W_34_31_i_13_n_0
);
W_34_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x102_out_26,
   I1 => x114_out_29,
   I2 => x114_out_1,
   I3 => x114_out_12,
   I4 => x115_out_26,
   O => W_34_31_i_14_n_0
);
W_34_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x102_out_29,
   I1 => x114_out_4,
   I2 => x114_out_15,
   I3 => x115_out_29,
   O => W_34_31_i_15_n_0
);
W_34_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x92_out_17,
   I1 => x92_out_15,
   O => SIGMA_LCASE_1243_out_0_30
);
W_34_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => x114_out_6,
   I1 => x114_out_17,
   I2 => x102_out_31,
   I3 => x115_out_31,
   I4 => x92_out_16,
   I5 => x92_out_18,
   O => W_34_31_i_17_n_0
);
W_34_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x114_out_16,
   I1 => x114_out_5,
   O => SIGMA_LCASE_0239_out_30
);
W_34_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x115_out_30,
   I1 => x102_out_30,
   I2 => x114_out_16,
   I3 => x114_out_5,
   O => W_34_31_i_19_n_0
);
W_34_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x92_out_14,
   I1 => x92_out_16,
   I2 => W_34_31_i_9_n_0,
   I3 => W_34_31_i_10_n_0,
   O => W_34_31_i_2_n_0
);
W_34_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x92_out_13,
   I1 => x92_out_15,
   I2 => W_34_31_i_11_n_0,
   I3 => W_34_31_i_12_n_0,
   O => W_34_31_i_3_n_0
);
W_34_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x92_out_12,
   I1 => x92_out_14,
   I2 => W_34_31_i_13_n_0,
   I3 => W_34_31_i_14_n_0,
   O => W_34_31_i_4_n_0
);
W_34_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_34_31_i_15_n_0,
   I1 => SIGMA_LCASE_1243_out_0_30,
   I2 => W_34_31_i_17_n_0,
   I3 => x102_out_30,
   I4 => SIGMA_LCASE_0239_out_30,
   I5 => x115_out_30,
   O => W_34_31_i_5_n_0
);
W_34_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_34_31_i_2_n_0,
   I1 => W_34_31_i_19_n_0,
   I2 => x92_out_15,
   I3 => x92_out_17,
   I4 => W_34_31_i_15_n_0,
   O => W_34_31_i_6_n_0
);
W_34_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x92_out_14,
   I1 => x92_out_16,
   I2 => W_34_31_i_9_n_0,
   I3 => W_34_31_i_10_n_0,
   I4 => W_34_31_i_3_n_0,
   O => W_34_31_i_7_n_0
);
W_34_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x92_out_13,
   I1 => x92_out_15,
   I2 => W_34_31_i_11_n_0,
   I3 => W_34_31_i_12_n_0,
   I4 => W_34_31_i_4_n_0,
   O => W_34_31_i_8_n_0
);
W_34_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x115_out_29,
   I1 => x102_out_29,
   I2 => x114_out_15,
   I3 => x114_out_4,
   O => W_34_31_i_9_n_0
);
W_34_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x115_out_2,
   I1 => x102_out_2,
   I2 => x114_out_20,
   I3 => x114_out_9,
   I4 => x114_out_5,
   O => W_34_3_i_10_n_0
);
W_34_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x102_out_1,
   I1 => x114_out_4,
   I2 => x114_out_8,
   I3 => x114_out_19,
   I4 => x115_out_1,
   O => W_34_3_i_11_n_0
);
W_34_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x114_out_19,
   I1 => x114_out_8,
   I2 => x114_out_4,
   O => SIGMA_LCASE_0239_out_1
);
W_34_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x92_out_21,
   I1 => x92_out_19,
   I2 => x92_out_12,
   O => SIGMA_LCASE_1243_out_0_2
);
W_34_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x92_out_20,
   I1 => x92_out_18,
   I2 => x92_out_11,
   O => SIGMA_LCASE_1243_out_1
);
W_34_3_i_15 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x115_out_1,
   I1 => x102_out_1,
   I2 => x114_out_19,
   I3 => x114_out_8,
   I4 => x114_out_4,
   O => W_34_3_i_15_n_0
);
W_34_3_i_16 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x114_out_18,
   I1 => x114_out_7,
   I2 => x114_out_3,
   O => SIGMA_LCASE_0239_out_0
);
W_34_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x92_out_12,
   I1 => x92_out_19,
   I2 => x92_out_21,
   I3 => W_34_3_i_10_n_0,
   I4 => W_34_3_i_11_n_0,
   O => W_34_3_i_2_n_0
);
W_34_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_34_3_i_11_n_0,
   I1 => x92_out_21,
   I2 => x92_out_19,
   I3 => x92_out_12,
   I4 => W_34_3_i_10_n_0,
   O => W_34_3_i_3_n_0
);
W_34_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_0239_out_1,
   I1 => x102_out_1,
   I2 => x115_out_1,
   I3 => x92_out_11,
   I4 => x92_out_18,
   I5 => x92_out_20,
   O => W_34_3_i_4_n_0
);
W_34_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x115_out_0,
   I1 => x102_out_0,
   I2 => x114_out_18,
   I3 => x114_out_7,
   I4 => x114_out_3,
   O => W_34_3_i_5_n_0
);
W_34_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_34_3_i_2_n_0,
   I1 => W_34_7_i_16_n_0,
   I2 => x92_out_13,
   I3 => x92_out_20,
   I4 => x92_out_22,
   I5 => W_34_7_i_17_n_0,
   O => W_34_3_i_6_n_0
);
W_34_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_34_3_i_10_n_0,
   I1 => SIGMA_LCASE_1243_out_0_2,
   I2 => x115_out_1,
   I3 => x102_out_1,
   I4 => SIGMA_LCASE_0239_out_1,
   I5 => SIGMA_LCASE_1243_out_1,
   O => W_34_3_i_7_n_0
);
W_34_3_i_8 : LUT5
  generic map(
   INIT => X"99969666"
  )
 port map (
   I0 => SIGMA_LCASE_1243_out_1,
   I1 => W_34_3_i_15_n_0,
   I2 => x115_out_0,
   I3 => SIGMA_LCASE_0239_out_0,
   I4 => x102_out_0,
   O => W_34_3_i_8_n_0
);
W_34_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_34_3_i_5_n_0,
   I1 => x92_out_10,
   I2 => x92_out_17,
   I3 => x92_out_19,
   O => W_34_3_i_9_n_0
);
W_34_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x115_out_6,
   I1 => x102_out_6,
   I2 => x114_out_24,
   I3 => x114_out_13,
   I4 => x114_out_9,
   O => W_34_7_i_10_n_0
);
W_34_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x102_out_5,
   I1 => x114_out_8,
   I2 => x114_out_12,
   I3 => x114_out_23,
   I4 => x115_out_5,
   O => W_34_7_i_11_n_0
);
W_34_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x115_out_5,
   I1 => x102_out_5,
   I2 => x114_out_23,
   I3 => x114_out_12,
   I4 => x114_out_8,
   O => W_34_7_i_12_n_0
);
W_34_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x102_out_4,
   I1 => x114_out_7,
   I2 => x114_out_11,
   I3 => x114_out_22,
   I4 => x115_out_4,
   O => W_34_7_i_13_n_0
);
W_34_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x115_out_4,
   I1 => x102_out_4,
   I2 => x114_out_22,
   I3 => x114_out_11,
   I4 => x114_out_7,
   O => W_34_7_i_14_n_0
);
W_34_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x102_out_3,
   I1 => x114_out_6,
   I2 => x114_out_10,
   I3 => x114_out_21,
   I4 => x115_out_3,
   O => W_34_7_i_15_n_0
);
W_34_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x115_out_3,
   I1 => x102_out_3,
   I2 => x114_out_21,
   I3 => x114_out_10,
   I4 => x114_out_6,
   O => W_34_7_i_16_n_0
);
W_34_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x102_out_2,
   I1 => x114_out_5,
   I2 => x114_out_9,
   I3 => x114_out_20,
   I4 => x115_out_2,
   O => W_34_7_i_17_n_0
);
W_34_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x92_out_16,
   I1 => x92_out_23,
   I2 => x92_out_25,
   I3 => W_34_7_i_10_n_0,
   I4 => W_34_7_i_11_n_0,
   O => W_34_7_i_2_n_0
);
W_34_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x92_out_15,
   I1 => x92_out_22,
   I2 => x92_out_24,
   I3 => W_34_7_i_12_n_0,
   I4 => W_34_7_i_13_n_0,
   O => W_34_7_i_3_n_0
);
W_34_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x92_out_14,
   I1 => x92_out_21,
   I2 => x92_out_23,
   I3 => W_34_7_i_14_n_0,
   I4 => W_34_7_i_15_n_0,
   O => W_34_7_i_4_n_0
);
W_34_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x92_out_13,
   I1 => x92_out_20,
   I2 => x92_out_22,
   I3 => W_34_7_i_16_n_0,
   I4 => W_34_7_i_17_n_0,
   O => W_34_7_i_5_n_0
);
W_34_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_34_7_i_2_n_0,
   I1 => W_34_11_i_16_n_0,
   I2 => x92_out_17,
   I3 => x92_out_24,
   I4 => x92_out_26,
   I5 => W_34_11_i_17_n_0,
   O => W_34_7_i_6_n_0
);
W_34_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_34_7_i_3_n_0,
   I1 => W_34_7_i_10_n_0,
   I2 => x92_out_16,
   I3 => x92_out_23,
   I4 => x92_out_25,
   I5 => W_34_7_i_11_n_0,
   O => W_34_7_i_7_n_0
);
W_34_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_34_7_i_4_n_0,
   I1 => W_34_7_i_12_n_0,
   I2 => x92_out_15,
   I3 => x92_out_22,
   I4 => x92_out_24,
   I5 => W_34_7_i_13_n_0,
   O => W_34_7_i_8_n_0
);
W_34_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_34_7_i_5_n_0,
   I1 => W_34_7_i_14_n_0,
   I2 => x92_out_14,
   I3 => x92_out_21,
   I4 => x92_out_23,
   I5 => W_34_7_i_15_n_0,
   O => W_34_7_i_9_n_0
);
W_35_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x114_out_10,
   I1 => x100_out_10,
   I2 => x113_out_28,
   I3 => x113_out_17,
   I4 => x113_out_13,
   O => W_35_11_i_10_n_0
);
W_35_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x100_out_9,
   I1 => x113_out_12,
   I2 => x113_out_16,
   I3 => x113_out_27,
   I4 => x114_out_9,
   O => W_35_11_i_11_n_0
);
W_35_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x114_out_9,
   I1 => x100_out_9,
   I2 => x113_out_27,
   I3 => x113_out_16,
   I4 => x113_out_12,
   O => W_35_11_i_12_n_0
);
W_35_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x100_out_8,
   I1 => x113_out_11,
   I2 => x113_out_15,
   I3 => x113_out_26,
   I4 => x114_out_8,
   O => W_35_11_i_13_n_0
);
W_35_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x114_out_8,
   I1 => x100_out_8,
   I2 => x113_out_26,
   I3 => x113_out_15,
   I4 => x113_out_11,
   O => W_35_11_i_14_n_0
);
W_35_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x100_out_7,
   I1 => x113_out_10,
   I2 => x113_out_14,
   I3 => x113_out_25,
   I4 => x114_out_7,
   O => W_35_11_i_15_n_0
);
W_35_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x114_out_7,
   I1 => x100_out_7,
   I2 => x113_out_25,
   I3 => x113_out_14,
   I4 => x113_out_10,
   O => W_35_11_i_16_n_0
);
W_35_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x100_out_6,
   I1 => x113_out_9,
   I2 => x113_out_13,
   I3 => x113_out_24,
   I4 => x114_out_6,
   O => W_35_11_i_17_n_0
);
W_35_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x89_out_20,
   I1 => x89_out_27,
   I2 => x89_out_29,
   I3 => W_35_11_i_10_n_0,
   I4 => W_35_11_i_11_n_0,
   O => W_35_11_i_2_n_0
);
W_35_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x89_out_19,
   I1 => x89_out_26,
   I2 => x89_out_28,
   I3 => W_35_11_i_12_n_0,
   I4 => W_35_11_i_13_n_0,
   O => W_35_11_i_3_n_0
);
W_35_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x89_out_18,
   I1 => x89_out_25,
   I2 => x89_out_27,
   I3 => W_35_11_i_14_n_0,
   I4 => W_35_11_i_15_n_0,
   O => W_35_11_i_4_n_0
);
W_35_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x89_out_17,
   I1 => x89_out_24,
   I2 => x89_out_26,
   I3 => W_35_11_i_16_n_0,
   I4 => W_35_11_i_17_n_0,
   O => W_35_11_i_5_n_0
);
W_35_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_35_11_i_2_n_0,
   I1 => W_35_15_i_16_n_0,
   I2 => x89_out_21,
   I3 => x89_out_28,
   I4 => x89_out_30,
   I5 => W_35_15_i_17_n_0,
   O => W_35_11_i_6_n_0
);
W_35_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_35_11_i_3_n_0,
   I1 => W_35_11_i_10_n_0,
   I2 => x89_out_20,
   I3 => x89_out_27,
   I4 => x89_out_29,
   I5 => W_35_11_i_11_n_0,
   O => W_35_11_i_7_n_0
);
W_35_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_35_11_i_4_n_0,
   I1 => W_35_11_i_12_n_0,
   I2 => x89_out_19,
   I3 => x89_out_26,
   I4 => x89_out_28,
   I5 => W_35_11_i_13_n_0,
   O => W_35_11_i_8_n_0
);
W_35_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_35_11_i_5_n_0,
   I1 => W_35_11_i_14_n_0,
   I2 => x89_out_18,
   I3 => x89_out_25,
   I4 => x89_out_27,
   I5 => W_35_11_i_15_n_0,
   O => W_35_11_i_9_n_0
);
W_35_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x114_out_14,
   I1 => x100_out_14,
   I2 => x113_out_0,
   I3 => x113_out_21,
   I4 => x113_out_17,
   O => W_35_15_i_10_n_0
);
W_35_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x100_out_13,
   I1 => x113_out_16,
   I2 => x113_out_20,
   I3 => x113_out_31,
   I4 => x114_out_13,
   O => W_35_15_i_11_n_0
);
W_35_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x114_out_13,
   I1 => x100_out_13,
   I2 => x113_out_31,
   I3 => x113_out_20,
   I4 => x113_out_16,
   O => W_35_15_i_12_n_0
);
W_35_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x100_out_12,
   I1 => x113_out_15,
   I2 => x113_out_19,
   I3 => x113_out_30,
   I4 => x114_out_12,
   O => W_35_15_i_13_n_0
);
W_35_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x114_out_12,
   I1 => x100_out_12,
   I2 => x113_out_30,
   I3 => x113_out_19,
   I4 => x113_out_15,
   O => W_35_15_i_14_n_0
);
W_35_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x100_out_11,
   I1 => x113_out_14,
   I2 => x113_out_18,
   I3 => x113_out_29,
   I4 => x114_out_11,
   O => W_35_15_i_15_n_0
);
W_35_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x114_out_11,
   I1 => x100_out_11,
   I2 => x113_out_29,
   I3 => x113_out_18,
   I4 => x113_out_14,
   O => W_35_15_i_16_n_0
);
W_35_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x100_out_10,
   I1 => x113_out_13,
   I2 => x113_out_17,
   I3 => x113_out_28,
   I4 => x114_out_10,
   O => W_35_15_i_17_n_0
);
W_35_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x89_out_24,
   I1 => x89_out_31,
   I2 => x89_out_1,
   I3 => W_35_15_i_10_n_0,
   I4 => W_35_15_i_11_n_0,
   O => W_35_15_i_2_n_0
);
W_35_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x89_out_23,
   I1 => x89_out_30,
   I2 => x89_out_0,
   I3 => W_35_15_i_12_n_0,
   I4 => W_35_15_i_13_n_0,
   O => W_35_15_i_3_n_0
);
W_35_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x89_out_22,
   I1 => x89_out_29,
   I2 => x89_out_31,
   I3 => W_35_15_i_14_n_0,
   I4 => W_35_15_i_15_n_0,
   O => W_35_15_i_4_n_0
);
W_35_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x89_out_21,
   I1 => x89_out_28,
   I2 => x89_out_30,
   I3 => W_35_15_i_16_n_0,
   I4 => W_35_15_i_17_n_0,
   O => W_35_15_i_5_n_0
);
W_35_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_35_15_i_2_n_0,
   I1 => W_35_19_i_16_n_0,
   I2 => x89_out_25,
   I3 => x89_out_0,
   I4 => x89_out_2,
   I5 => W_35_19_i_17_n_0,
   O => W_35_15_i_6_n_0
);
W_35_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_35_15_i_3_n_0,
   I1 => W_35_15_i_10_n_0,
   I2 => x89_out_24,
   I3 => x89_out_31,
   I4 => x89_out_1,
   I5 => W_35_15_i_11_n_0,
   O => W_35_15_i_7_n_0
);
W_35_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_35_15_i_4_n_0,
   I1 => W_35_15_i_12_n_0,
   I2 => x89_out_23,
   I3 => x89_out_30,
   I4 => x89_out_0,
   I5 => W_35_15_i_13_n_0,
   O => W_35_15_i_8_n_0
);
W_35_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_35_15_i_5_n_0,
   I1 => W_35_15_i_14_n_0,
   I2 => x89_out_22,
   I3 => x89_out_29,
   I4 => x89_out_31,
   I5 => W_35_15_i_15_n_0,
   O => W_35_15_i_9_n_0
);
W_35_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x114_out_18,
   I1 => x100_out_18,
   I2 => x113_out_4,
   I3 => x113_out_25,
   I4 => x113_out_21,
   O => W_35_19_i_10_n_0
);
W_35_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x100_out_17,
   I1 => x113_out_20,
   I2 => x113_out_24,
   I3 => x113_out_3,
   I4 => x114_out_17,
   O => W_35_19_i_11_n_0
);
W_35_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x114_out_17,
   I1 => x100_out_17,
   I2 => x113_out_3,
   I3 => x113_out_24,
   I4 => x113_out_20,
   O => W_35_19_i_12_n_0
);
W_35_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x100_out_16,
   I1 => x113_out_19,
   I2 => x113_out_23,
   I3 => x113_out_2,
   I4 => x114_out_16,
   O => W_35_19_i_13_n_0
);
W_35_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x114_out_16,
   I1 => x100_out_16,
   I2 => x113_out_2,
   I3 => x113_out_23,
   I4 => x113_out_19,
   O => W_35_19_i_14_n_0
);
W_35_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x100_out_15,
   I1 => x113_out_18,
   I2 => x113_out_22,
   I3 => x113_out_1,
   I4 => x114_out_15,
   O => W_35_19_i_15_n_0
);
W_35_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x114_out_15,
   I1 => x100_out_15,
   I2 => x113_out_1,
   I3 => x113_out_22,
   I4 => x113_out_18,
   O => W_35_19_i_16_n_0
);
W_35_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x100_out_14,
   I1 => x113_out_17,
   I2 => x113_out_21,
   I3 => x113_out_0,
   I4 => x114_out_14,
   O => W_35_19_i_17_n_0
);
W_35_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x89_out_28,
   I1 => x89_out_3,
   I2 => x89_out_5,
   I3 => W_35_19_i_10_n_0,
   I4 => W_35_19_i_11_n_0,
   O => W_35_19_i_2_n_0
);
W_35_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x89_out_27,
   I1 => x89_out_2,
   I2 => x89_out_4,
   I3 => W_35_19_i_12_n_0,
   I4 => W_35_19_i_13_n_0,
   O => W_35_19_i_3_n_0
);
W_35_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x89_out_26,
   I1 => x89_out_1,
   I2 => x89_out_3,
   I3 => W_35_19_i_14_n_0,
   I4 => W_35_19_i_15_n_0,
   O => W_35_19_i_4_n_0
);
W_35_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x89_out_25,
   I1 => x89_out_0,
   I2 => x89_out_2,
   I3 => W_35_19_i_16_n_0,
   I4 => W_35_19_i_17_n_0,
   O => W_35_19_i_5_n_0
);
W_35_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_35_19_i_2_n_0,
   I1 => W_35_23_i_16_n_0,
   I2 => x89_out_29,
   I3 => x89_out_4,
   I4 => x89_out_6,
   I5 => W_35_23_i_17_n_0,
   O => W_35_19_i_6_n_0
);
W_35_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_35_19_i_3_n_0,
   I1 => W_35_19_i_10_n_0,
   I2 => x89_out_28,
   I3 => x89_out_3,
   I4 => x89_out_5,
   I5 => W_35_19_i_11_n_0,
   O => W_35_19_i_7_n_0
);
W_35_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_35_19_i_4_n_0,
   I1 => W_35_19_i_12_n_0,
   I2 => x89_out_27,
   I3 => x89_out_2,
   I4 => x89_out_4,
   I5 => W_35_19_i_13_n_0,
   O => W_35_19_i_8_n_0
);
W_35_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_35_19_i_5_n_0,
   I1 => W_35_19_i_14_n_0,
   I2 => x89_out_26,
   I3 => x89_out_1,
   I4 => x89_out_3,
   I5 => W_35_19_i_15_n_0,
   O => W_35_19_i_9_n_0
);
W_35_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x114_out_22,
   I1 => x100_out_22,
   I2 => x113_out_8,
   I3 => x113_out_29,
   I4 => x113_out_25,
   O => W_35_23_i_10_n_0
);
W_35_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x100_out_21,
   I1 => x113_out_24,
   I2 => x113_out_28,
   I3 => x113_out_7,
   I4 => x114_out_21,
   O => W_35_23_i_11_n_0
);
W_35_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x114_out_21,
   I1 => x100_out_21,
   I2 => x113_out_7,
   I3 => x113_out_28,
   I4 => x113_out_24,
   O => W_35_23_i_12_n_0
);
W_35_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x100_out_20,
   I1 => x113_out_23,
   I2 => x113_out_27,
   I3 => x113_out_6,
   I4 => x114_out_20,
   O => W_35_23_i_13_n_0
);
W_35_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x114_out_20,
   I1 => x100_out_20,
   I2 => x113_out_6,
   I3 => x113_out_27,
   I4 => x113_out_23,
   O => W_35_23_i_14_n_0
);
W_35_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x100_out_19,
   I1 => x113_out_22,
   I2 => x113_out_26,
   I3 => x113_out_5,
   I4 => x114_out_19,
   O => W_35_23_i_15_n_0
);
W_35_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x114_out_19,
   I1 => x100_out_19,
   I2 => x113_out_5,
   I3 => x113_out_26,
   I4 => x113_out_22,
   O => W_35_23_i_16_n_0
);
W_35_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x100_out_18,
   I1 => x113_out_21,
   I2 => x113_out_25,
   I3 => x113_out_4,
   I4 => x114_out_18,
   O => W_35_23_i_17_n_0
);
W_35_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x89_out_7,
   I1 => x89_out_9,
   I2 => W_35_23_i_10_n_0,
   I3 => W_35_23_i_11_n_0,
   O => W_35_23_i_2_n_0
);
W_35_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x89_out_31,
   I1 => x89_out_6,
   I2 => x89_out_8,
   I3 => W_35_23_i_12_n_0,
   I4 => W_35_23_i_13_n_0,
   O => W_35_23_i_3_n_0
);
W_35_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x89_out_30,
   I1 => x89_out_5,
   I2 => x89_out_7,
   I3 => W_35_23_i_14_n_0,
   I4 => W_35_23_i_15_n_0,
   O => W_35_23_i_4_n_0
);
W_35_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x89_out_29,
   I1 => x89_out_4,
   I2 => x89_out_6,
   I3 => W_35_23_i_16_n_0,
   I4 => W_35_23_i_17_n_0,
   O => W_35_23_i_5_n_0
);
W_35_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x89_out_8,
   I1 => x89_out_10,
   I2 => W_35_27_i_16_n_0,
   I3 => W_35_27_i_17_n_0,
   I4 => W_35_23_i_2_n_0,
   O => W_35_23_i_6_n_0
);
W_35_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x89_out_7,
   I1 => x89_out_9,
   I2 => W_35_23_i_10_n_0,
   I3 => W_35_23_i_11_n_0,
   I4 => W_35_23_i_3_n_0,
   O => W_35_23_i_7_n_0
);
W_35_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_35_23_i_4_n_0,
   I1 => W_35_23_i_12_n_0,
   I2 => x89_out_31,
   I3 => x89_out_6,
   I4 => x89_out_8,
   I5 => W_35_23_i_13_n_0,
   O => W_35_23_i_8_n_0
);
W_35_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_35_23_i_5_n_0,
   I1 => W_35_23_i_14_n_0,
   I2 => x89_out_30,
   I3 => x89_out_5,
   I4 => x89_out_7,
   I5 => W_35_23_i_15_n_0,
   O => W_35_23_i_9_n_0
);
W_35_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x114_out_26,
   I1 => x100_out_26,
   I2 => x113_out_12,
   I3 => x113_out_1,
   I4 => x113_out_29,
   O => W_35_27_i_10_n_0
);
W_35_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x100_out_25,
   I1 => x113_out_28,
   I2 => x113_out_0,
   I3 => x113_out_11,
   I4 => x114_out_25,
   O => W_35_27_i_11_n_0
);
W_35_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x114_out_25,
   I1 => x100_out_25,
   I2 => x113_out_11,
   I3 => x113_out_0,
   I4 => x113_out_28,
   O => W_35_27_i_12_n_0
);
W_35_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x100_out_24,
   I1 => x113_out_27,
   I2 => x113_out_31,
   I3 => x113_out_10,
   I4 => x114_out_24,
   O => W_35_27_i_13_n_0
);
W_35_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x114_out_24,
   I1 => x100_out_24,
   I2 => x113_out_10,
   I3 => x113_out_31,
   I4 => x113_out_27,
   O => W_35_27_i_14_n_0
);
W_35_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x100_out_23,
   I1 => x113_out_26,
   I2 => x113_out_30,
   I3 => x113_out_9,
   I4 => x114_out_23,
   O => W_35_27_i_15_n_0
);
W_35_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x114_out_23,
   I1 => x100_out_23,
   I2 => x113_out_9,
   I3 => x113_out_30,
   I4 => x113_out_26,
   O => W_35_27_i_16_n_0
);
W_35_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x100_out_22,
   I1 => x113_out_25,
   I2 => x113_out_29,
   I3 => x113_out_8,
   I4 => x114_out_22,
   O => W_35_27_i_17_n_0
);
W_35_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x89_out_11,
   I1 => x89_out_13,
   I2 => W_35_27_i_10_n_0,
   I3 => W_35_27_i_11_n_0,
   O => W_35_27_i_2_n_0
);
W_35_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x89_out_10,
   I1 => x89_out_12,
   I2 => W_35_27_i_12_n_0,
   I3 => W_35_27_i_13_n_0,
   O => W_35_27_i_3_n_0
);
W_35_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x89_out_9,
   I1 => x89_out_11,
   I2 => W_35_27_i_14_n_0,
   I3 => W_35_27_i_15_n_0,
   O => W_35_27_i_4_n_0
);
W_35_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x89_out_8,
   I1 => x89_out_10,
   I2 => W_35_27_i_16_n_0,
   I3 => W_35_27_i_17_n_0,
   O => W_35_27_i_5_n_0
);
W_35_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x89_out_12,
   I1 => x89_out_14,
   I2 => W_35_31_i_13_n_0,
   I3 => W_35_31_i_14_n_0,
   I4 => W_35_27_i_2_n_0,
   O => W_35_27_i_6_n_0
);
W_35_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x89_out_11,
   I1 => x89_out_13,
   I2 => W_35_27_i_10_n_0,
   I3 => W_35_27_i_11_n_0,
   I4 => W_35_27_i_3_n_0,
   O => W_35_27_i_7_n_0
);
W_35_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x89_out_10,
   I1 => x89_out_12,
   I2 => W_35_27_i_12_n_0,
   I3 => W_35_27_i_13_n_0,
   I4 => W_35_27_i_4_n_0,
   O => W_35_27_i_8_n_0
);
W_35_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x89_out_9,
   I1 => x89_out_11,
   I2 => W_35_27_i_14_n_0,
   I3 => W_35_27_i_15_n_0,
   I4 => W_35_27_i_5_n_0,
   O => W_35_27_i_9_n_0
);
W_35_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x100_out_28,
   I1 => x113_out_31,
   I2 => x113_out_3,
   I3 => x113_out_14,
   I4 => x114_out_28,
   O => W_35_31_i_10_n_0
);
W_35_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x114_out_28,
   I1 => x100_out_28,
   I2 => x113_out_14,
   I3 => x113_out_3,
   I4 => x113_out_31,
   O => W_35_31_i_11_n_0
);
W_35_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x100_out_27,
   I1 => x113_out_30,
   I2 => x113_out_2,
   I3 => x113_out_13,
   I4 => x114_out_27,
   O => W_35_31_i_12_n_0
);
W_35_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x114_out_27,
   I1 => x100_out_27,
   I2 => x113_out_13,
   I3 => x113_out_2,
   I4 => x113_out_30,
   O => W_35_31_i_13_n_0
);
W_35_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x100_out_26,
   I1 => x113_out_29,
   I2 => x113_out_1,
   I3 => x113_out_12,
   I4 => x114_out_26,
   O => W_35_31_i_14_n_0
);
W_35_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x100_out_29,
   I1 => x113_out_4,
   I2 => x113_out_15,
   I3 => x114_out_29,
   O => W_35_31_i_15_n_0
);
W_35_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x89_out_17,
   I1 => x89_out_15,
   O => SIGMA_LCASE_1235_out_0_30
);
W_35_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => x113_out_6,
   I1 => x113_out_17,
   I2 => x100_out_31,
   I3 => x114_out_31,
   I4 => x89_out_16,
   I5 => x89_out_18,
   O => W_35_31_i_17_n_0
);
W_35_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x113_out_16,
   I1 => x113_out_5,
   O => SIGMA_LCASE_0231_out_30
);
W_35_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x114_out_30,
   I1 => x100_out_30,
   I2 => x113_out_16,
   I3 => x113_out_5,
   O => W_35_31_i_19_n_0
);
W_35_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x89_out_14,
   I1 => x89_out_16,
   I2 => W_35_31_i_9_n_0,
   I3 => W_35_31_i_10_n_0,
   O => W_35_31_i_2_n_0
);
W_35_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x89_out_13,
   I1 => x89_out_15,
   I2 => W_35_31_i_11_n_0,
   I3 => W_35_31_i_12_n_0,
   O => W_35_31_i_3_n_0
);
W_35_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x89_out_12,
   I1 => x89_out_14,
   I2 => W_35_31_i_13_n_0,
   I3 => W_35_31_i_14_n_0,
   O => W_35_31_i_4_n_0
);
W_35_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_35_31_i_15_n_0,
   I1 => SIGMA_LCASE_1235_out_0_30,
   I2 => W_35_31_i_17_n_0,
   I3 => x100_out_30,
   I4 => SIGMA_LCASE_0231_out_30,
   I5 => x114_out_30,
   O => W_35_31_i_5_n_0
);
W_35_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_35_31_i_2_n_0,
   I1 => W_35_31_i_19_n_0,
   I2 => x89_out_15,
   I3 => x89_out_17,
   I4 => W_35_31_i_15_n_0,
   O => W_35_31_i_6_n_0
);
W_35_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x89_out_14,
   I1 => x89_out_16,
   I2 => W_35_31_i_9_n_0,
   I3 => W_35_31_i_10_n_0,
   I4 => W_35_31_i_3_n_0,
   O => W_35_31_i_7_n_0
);
W_35_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x89_out_13,
   I1 => x89_out_15,
   I2 => W_35_31_i_11_n_0,
   I3 => W_35_31_i_12_n_0,
   I4 => W_35_31_i_4_n_0,
   O => W_35_31_i_8_n_0
);
W_35_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x114_out_29,
   I1 => x100_out_29,
   I2 => x113_out_15,
   I3 => x113_out_4,
   O => W_35_31_i_9_n_0
);
W_35_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x114_out_2,
   I1 => x100_out_2,
   I2 => x113_out_20,
   I3 => x113_out_9,
   I4 => x113_out_5,
   O => W_35_3_i_10_n_0
);
W_35_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x100_out_1,
   I1 => x113_out_4,
   I2 => x113_out_8,
   I3 => x113_out_19,
   I4 => x114_out_1,
   O => W_35_3_i_11_n_0
);
W_35_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x113_out_19,
   I1 => x113_out_8,
   I2 => x113_out_4,
   O => SIGMA_LCASE_0231_out_1
);
W_35_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x89_out_21,
   I1 => x89_out_19,
   I2 => x89_out_12,
   O => SIGMA_LCASE_1235_out_0_2
);
W_35_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x89_out_20,
   I1 => x89_out_18,
   I2 => x89_out_11,
   O => SIGMA_LCASE_1235_out_1
);
W_35_3_i_15 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x114_out_1,
   I1 => x100_out_1,
   I2 => x113_out_19,
   I3 => x113_out_8,
   I4 => x113_out_4,
   O => W_35_3_i_15_n_0
);
W_35_3_i_16 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x113_out_18,
   I1 => x113_out_7,
   I2 => x113_out_3,
   O => SIGMA_LCASE_0231_out_0
);
W_35_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x89_out_12,
   I1 => x89_out_19,
   I2 => x89_out_21,
   I3 => W_35_3_i_10_n_0,
   I4 => W_35_3_i_11_n_0,
   O => W_35_3_i_2_n_0
);
W_35_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_35_3_i_11_n_0,
   I1 => x89_out_21,
   I2 => x89_out_19,
   I3 => x89_out_12,
   I4 => W_35_3_i_10_n_0,
   O => W_35_3_i_3_n_0
);
W_35_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_0231_out_1,
   I1 => x100_out_1,
   I2 => x114_out_1,
   I3 => x89_out_11,
   I4 => x89_out_18,
   I5 => x89_out_20,
   O => W_35_3_i_4_n_0
);
W_35_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x114_out_0,
   I1 => x100_out_0,
   I2 => x113_out_18,
   I3 => x113_out_7,
   I4 => x113_out_3,
   O => W_35_3_i_5_n_0
);
W_35_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_35_3_i_2_n_0,
   I1 => W_35_7_i_16_n_0,
   I2 => x89_out_13,
   I3 => x89_out_20,
   I4 => x89_out_22,
   I5 => W_35_7_i_17_n_0,
   O => W_35_3_i_6_n_0
);
W_35_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_35_3_i_10_n_0,
   I1 => SIGMA_LCASE_1235_out_0_2,
   I2 => x114_out_1,
   I3 => x100_out_1,
   I4 => SIGMA_LCASE_0231_out_1,
   I5 => SIGMA_LCASE_1235_out_1,
   O => W_35_3_i_7_n_0
);
W_35_3_i_8 : LUT5
  generic map(
   INIT => X"99969666"
  )
 port map (
   I0 => SIGMA_LCASE_1235_out_1,
   I1 => W_35_3_i_15_n_0,
   I2 => x114_out_0,
   I3 => SIGMA_LCASE_0231_out_0,
   I4 => x100_out_0,
   O => W_35_3_i_8_n_0
);
W_35_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_35_3_i_5_n_0,
   I1 => x89_out_10,
   I2 => x89_out_17,
   I3 => x89_out_19,
   O => W_35_3_i_9_n_0
);
W_35_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x114_out_6,
   I1 => x100_out_6,
   I2 => x113_out_24,
   I3 => x113_out_13,
   I4 => x113_out_9,
   O => W_35_7_i_10_n_0
);
W_35_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x100_out_5,
   I1 => x113_out_8,
   I2 => x113_out_12,
   I3 => x113_out_23,
   I4 => x114_out_5,
   O => W_35_7_i_11_n_0
);
W_35_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x114_out_5,
   I1 => x100_out_5,
   I2 => x113_out_23,
   I3 => x113_out_12,
   I4 => x113_out_8,
   O => W_35_7_i_12_n_0
);
W_35_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x100_out_4,
   I1 => x113_out_7,
   I2 => x113_out_11,
   I3 => x113_out_22,
   I4 => x114_out_4,
   O => W_35_7_i_13_n_0
);
W_35_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x114_out_4,
   I1 => x100_out_4,
   I2 => x113_out_22,
   I3 => x113_out_11,
   I4 => x113_out_7,
   O => W_35_7_i_14_n_0
);
W_35_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x100_out_3,
   I1 => x113_out_6,
   I2 => x113_out_10,
   I3 => x113_out_21,
   I4 => x114_out_3,
   O => W_35_7_i_15_n_0
);
W_35_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x114_out_3,
   I1 => x100_out_3,
   I2 => x113_out_21,
   I3 => x113_out_10,
   I4 => x113_out_6,
   O => W_35_7_i_16_n_0
);
W_35_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x100_out_2,
   I1 => x113_out_5,
   I2 => x113_out_9,
   I3 => x113_out_20,
   I4 => x114_out_2,
   O => W_35_7_i_17_n_0
);
W_35_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x89_out_16,
   I1 => x89_out_23,
   I2 => x89_out_25,
   I3 => W_35_7_i_10_n_0,
   I4 => W_35_7_i_11_n_0,
   O => W_35_7_i_2_n_0
);
W_35_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x89_out_15,
   I1 => x89_out_22,
   I2 => x89_out_24,
   I3 => W_35_7_i_12_n_0,
   I4 => W_35_7_i_13_n_0,
   O => W_35_7_i_3_n_0
);
W_35_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x89_out_14,
   I1 => x89_out_21,
   I2 => x89_out_23,
   I3 => W_35_7_i_14_n_0,
   I4 => W_35_7_i_15_n_0,
   O => W_35_7_i_4_n_0
);
W_35_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x89_out_13,
   I1 => x89_out_20,
   I2 => x89_out_22,
   I3 => W_35_7_i_16_n_0,
   I4 => W_35_7_i_17_n_0,
   O => W_35_7_i_5_n_0
);
W_35_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_35_7_i_2_n_0,
   I1 => W_35_11_i_16_n_0,
   I2 => x89_out_17,
   I3 => x89_out_24,
   I4 => x89_out_26,
   I5 => W_35_11_i_17_n_0,
   O => W_35_7_i_6_n_0
);
W_35_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_35_7_i_3_n_0,
   I1 => W_35_7_i_10_n_0,
   I2 => x89_out_16,
   I3 => x89_out_23,
   I4 => x89_out_25,
   I5 => W_35_7_i_11_n_0,
   O => W_35_7_i_7_n_0
);
W_35_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_35_7_i_4_n_0,
   I1 => W_35_7_i_12_n_0,
   I2 => x89_out_15,
   I3 => x89_out_22,
   I4 => x89_out_24,
   I5 => W_35_7_i_13_n_0,
   O => W_35_7_i_8_n_0
);
W_35_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_35_7_i_5_n_0,
   I1 => W_35_7_i_14_n_0,
   I2 => x89_out_14,
   I3 => x89_out_21,
   I4 => x89_out_23,
   I5 => W_35_7_i_15_n_0,
   O => W_35_7_i_9_n_0
);
W_36_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x113_out_10,
   I1 => x98_out_10,
   I2 => x112_out_28,
   I3 => x112_out_17,
   I4 => x112_out_13,
   O => W_36_11_i_10_n_0
);
W_36_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x98_out_9,
   I1 => x112_out_12,
   I2 => x112_out_16,
   I3 => x112_out_27,
   I4 => x113_out_9,
   O => W_36_11_i_11_n_0
);
W_36_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x113_out_9,
   I1 => x98_out_9,
   I2 => x112_out_27,
   I3 => x112_out_16,
   I4 => x112_out_12,
   O => W_36_11_i_12_n_0
);
W_36_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x98_out_8,
   I1 => x112_out_11,
   I2 => x112_out_15,
   I3 => x112_out_26,
   I4 => x113_out_8,
   O => W_36_11_i_13_n_0
);
W_36_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x113_out_8,
   I1 => x98_out_8,
   I2 => x112_out_26,
   I3 => x112_out_15,
   I4 => x112_out_11,
   O => W_36_11_i_14_n_0
);
W_36_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x98_out_7,
   I1 => x112_out_10,
   I2 => x112_out_14,
   I3 => x112_out_25,
   I4 => x113_out_7,
   O => W_36_11_i_15_n_0
);
W_36_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x113_out_7,
   I1 => x98_out_7,
   I2 => x112_out_25,
   I3 => x112_out_14,
   I4 => x112_out_10,
   O => W_36_11_i_16_n_0
);
W_36_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x98_out_6,
   I1 => x112_out_9,
   I2 => x112_out_13,
   I3 => x112_out_24,
   I4 => x113_out_6,
   O => W_36_11_i_17_n_0
);
W_36_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x86_out_20,
   I1 => x86_out_27,
   I2 => x86_out_29,
   I3 => W_36_11_i_10_n_0,
   I4 => W_36_11_i_11_n_0,
   O => W_36_11_i_2_n_0
);
W_36_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x86_out_19,
   I1 => x86_out_26,
   I2 => x86_out_28,
   I3 => W_36_11_i_12_n_0,
   I4 => W_36_11_i_13_n_0,
   O => W_36_11_i_3_n_0
);
W_36_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x86_out_18,
   I1 => x86_out_25,
   I2 => x86_out_27,
   I3 => W_36_11_i_14_n_0,
   I4 => W_36_11_i_15_n_0,
   O => W_36_11_i_4_n_0
);
W_36_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x86_out_17,
   I1 => x86_out_24,
   I2 => x86_out_26,
   I3 => W_36_11_i_16_n_0,
   I4 => W_36_11_i_17_n_0,
   O => W_36_11_i_5_n_0
);
W_36_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_36_11_i_2_n_0,
   I1 => W_36_15_i_16_n_0,
   I2 => x86_out_21,
   I3 => x86_out_28,
   I4 => x86_out_30,
   I5 => W_36_15_i_17_n_0,
   O => W_36_11_i_6_n_0
);
W_36_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_36_11_i_3_n_0,
   I1 => W_36_11_i_10_n_0,
   I2 => x86_out_20,
   I3 => x86_out_27,
   I4 => x86_out_29,
   I5 => W_36_11_i_11_n_0,
   O => W_36_11_i_7_n_0
);
W_36_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_36_11_i_4_n_0,
   I1 => W_36_11_i_12_n_0,
   I2 => x86_out_19,
   I3 => x86_out_26,
   I4 => x86_out_28,
   I5 => W_36_11_i_13_n_0,
   O => W_36_11_i_8_n_0
);
W_36_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_36_11_i_5_n_0,
   I1 => W_36_11_i_14_n_0,
   I2 => x86_out_18,
   I3 => x86_out_25,
   I4 => x86_out_27,
   I5 => W_36_11_i_15_n_0,
   O => W_36_11_i_9_n_0
);
W_36_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x113_out_14,
   I1 => x98_out_14,
   I2 => x112_out_0,
   I3 => x112_out_21,
   I4 => x112_out_17,
   O => W_36_15_i_10_n_0
);
W_36_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x98_out_13,
   I1 => x112_out_16,
   I2 => x112_out_20,
   I3 => x112_out_31,
   I4 => x113_out_13,
   O => W_36_15_i_11_n_0
);
W_36_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x113_out_13,
   I1 => x98_out_13,
   I2 => x112_out_31,
   I3 => x112_out_20,
   I4 => x112_out_16,
   O => W_36_15_i_12_n_0
);
W_36_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x98_out_12,
   I1 => x112_out_15,
   I2 => x112_out_19,
   I3 => x112_out_30,
   I4 => x113_out_12,
   O => W_36_15_i_13_n_0
);
W_36_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x113_out_12,
   I1 => x98_out_12,
   I2 => x112_out_30,
   I3 => x112_out_19,
   I4 => x112_out_15,
   O => W_36_15_i_14_n_0
);
W_36_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x98_out_11,
   I1 => x112_out_14,
   I2 => x112_out_18,
   I3 => x112_out_29,
   I4 => x113_out_11,
   O => W_36_15_i_15_n_0
);
W_36_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x113_out_11,
   I1 => x98_out_11,
   I2 => x112_out_29,
   I3 => x112_out_18,
   I4 => x112_out_14,
   O => W_36_15_i_16_n_0
);
W_36_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x98_out_10,
   I1 => x112_out_13,
   I2 => x112_out_17,
   I3 => x112_out_28,
   I4 => x113_out_10,
   O => W_36_15_i_17_n_0
);
W_36_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x86_out_24,
   I1 => x86_out_31,
   I2 => x86_out_1,
   I3 => W_36_15_i_10_n_0,
   I4 => W_36_15_i_11_n_0,
   O => W_36_15_i_2_n_0
);
W_36_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x86_out_23,
   I1 => x86_out_30,
   I2 => x86_out_0,
   I3 => W_36_15_i_12_n_0,
   I4 => W_36_15_i_13_n_0,
   O => W_36_15_i_3_n_0
);
W_36_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x86_out_22,
   I1 => x86_out_29,
   I2 => x86_out_31,
   I3 => W_36_15_i_14_n_0,
   I4 => W_36_15_i_15_n_0,
   O => W_36_15_i_4_n_0
);
W_36_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x86_out_21,
   I1 => x86_out_28,
   I2 => x86_out_30,
   I3 => W_36_15_i_16_n_0,
   I4 => W_36_15_i_17_n_0,
   O => W_36_15_i_5_n_0
);
W_36_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_36_15_i_2_n_0,
   I1 => W_36_19_i_16_n_0,
   I2 => x86_out_25,
   I3 => x86_out_0,
   I4 => x86_out_2,
   I5 => W_36_19_i_17_n_0,
   O => W_36_15_i_6_n_0
);
W_36_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_36_15_i_3_n_0,
   I1 => W_36_15_i_10_n_0,
   I2 => x86_out_24,
   I3 => x86_out_31,
   I4 => x86_out_1,
   I5 => W_36_15_i_11_n_0,
   O => W_36_15_i_7_n_0
);
W_36_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_36_15_i_4_n_0,
   I1 => W_36_15_i_12_n_0,
   I2 => x86_out_23,
   I3 => x86_out_30,
   I4 => x86_out_0,
   I5 => W_36_15_i_13_n_0,
   O => W_36_15_i_8_n_0
);
W_36_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_36_15_i_5_n_0,
   I1 => W_36_15_i_14_n_0,
   I2 => x86_out_22,
   I3 => x86_out_29,
   I4 => x86_out_31,
   I5 => W_36_15_i_15_n_0,
   O => W_36_15_i_9_n_0
);
W_36_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x113_out_18,
   I1 => x98_out_18,
   I2 => x112_out_4,
   I3 => x112_out_25,
   I4 => x112_out_21,
   O => W_36_19_i_10_n_0
);
W_36_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x98_out_17,
   I1 => x112_out_20,
   I2 => x112_out_24,
   I3 => x112_out_3,
   I4 => x113_out_17,
   O => W_36_19_i_11_n_0
);
W_36_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x113_out_17,
   I1 => x98_out_17,
   I2 => x112_out_3,
   I3 => x112_out_24,
   I4 => x112_out_20,
   O => W_36_19_i_12_n_0
);
W_36_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x98_out_16,
   I1 => x112_out_19,
   I2 => x112_out_23,
   I3 => x112_out_2,
   I4 => x113_out_16,
   O => W_36_19_i_13_n_0
);
W_36_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x113_out_16,
   I1 => x98_out_16,
   I2 => x112_out_2,
   I3 => x112_out_23,
   I4 => x112_out_19,
   O => W_36_19_i_14_n_0
);
W_36_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x98_out_15,
   I1 => x112_out_18,
   I2 => x112_out_22,
   I3 => x112_out_1,
   I4 => x113_out_15,
   O => W_36_19_i_15_n_0
);
W_36_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x113_out_15,
   I1 => x98_out_15,
   I2 => x112_out_1,
   I3 => x112_out_22,
   I4 => x112_out_18,
   O => W_36_19_i_16_n_0
);
W_36_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x98_out_14,
   I1 => x112_out_17,
   I2 => x112_out_21,
   I3 => x112_out_0,
   I4 => x113_out_14,
   O => W_36_19_i_17_n_0
);
W_36_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x86_out_28,
   I1 => x86_out_3,
   I2 => x86_out_5,
   I3 => W_36_19_i_10_n_0,
   I4 => W_36_19_i_11_n_0,
   O => W_36_19_i_2_n_0
);
W_36_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x86_out_27,
   I1 => x86_out_2,
   I2 => x86_out_4,
   I3 => W_36_19_i_12_n_0,
   I4 => W_36_19_i_13_n_0,
   O => W_36_19_i_3_n_0
);
W_36_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x86_out_26,
   I1 => x86_out_1,
   I2 => x86_out_3,
   I3 => W_36_19_i_14_n_0,
   I4 => W_36_19_i_15_n_0,
   O => W_36_19_i_4_n_0
);
W_36_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x86_out_25,
   I1 => x86_out_0,
   I2 => x86_out_2,
   I3 => W_36_19_i_16_n_0,
   I4 => W_36_19_i_17_n_0,
   O => W_36_19_i_5_n_0
);
W_36_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_36_19_i_2_n_0,
   I1 => W_36_23_i_16_n_0,
   I2 => x86_out_29,
   I3 => x86_out_4,
   I4 => x86_out_6,
   I5 => W_36_23_i_17_n_0,
   O => W_36_19_i_6_n_0
);
W_36_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_36_19_i_3_n_0,
   I1 => W_36_19_i_10_n_0,
   I2 => x86_out_28,
   I3 => x86_out_3,
   I4 => x86_out_5,
   I5 => W_36_19_i_11_n_0,
   O => W_36_19_i_7_n_0
);
W_36_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_36_19_i_4_n_0,
   I1 => W_36_19_i_12_n_0,
   I2 => x86_out_27,
   I3 => x86_out_2,
   I4 => x86_out_4,
   I5 => W_36_19_i_13_n_0,
   O => W_36_19_i_8_n_0
);
W_36_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_36_19_i_5_n_0,
   I1 => W_36_19_i_14_n_0,
   I2 => x86_out_26,
   I3 => x86_out_1,
   I4 => x86_out_3,
   I5 => W_36_19_i_15_n_0,
   O => W_36_19_i_9_n_0
);
W_36_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x113_out_22,
   I1 => x98_out_22,
   I2 => x112_out_8,
   I3 => x112_out_29,
   I4 => x112_out_25,
   O => W_36_23_i_10_n_0
);
W_36_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x98_out_21,
   I1 => x112_out_24,
   I2 => x112_out_28,
   I3 => x112_out_7,
   I4 => x113_out_21,
   O => W_36_23_i_11_n_0
);
W_36_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x113_out_21,
   I1 => x98_out_21,
   I2 => x112_out_7,
   I3 => x112_out_28,
   I4 => x112_out_24,
   O => W_36_23_i_12_n_0
);
W_36_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x98_out_20,
   I1 => x112_out_23,
   I2 => x112_out_27,
   I3 => x112_out_6,
   I4 => x113_out_20,
   O => W_36_23_i_13_n_0
);
W_36_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x113_out_20,
   I1 => x98_out_20,
   I2 => x112_out_6,
   I3 => x112_out_27,
   I4 => x112_out_23,
   O => W_36_23_i_14_n_0
);
W_36_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x98_out_19,
   I1 => x112_out_22,
   I2 => x112_out_26,
   I3 => x112_out_5,
   I4 => x113_out_19,
   O => W_36_23_i_15_n_0
);
W_36_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x113_out_19,
   I1 => x98_out_19,
   I2 => x112_out_5,
   I3 => x112_out_26,
   I4 => x112_out_22,
   O => W_36_23_i_16_n_0
);
W_36_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x98_out_18,
   I1 => x112_out_21,
   I2 => x112_out_25,
   I3 => x112_out_4,
   I4 => x113_out_18,
   O => W_36_23_i_17_n_0
);
W_36_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x86_out_7,
   I1 => x86_out_9,
   I2 => W_36_23_i_10_n_0,
   I3 => W_36_23_i_11_n_0,
   O => W_36_23_i_2_n_0
);
W_36_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x86_out_31,
   I1 => x86_out_6,
   I2 => x86_out_8,
   I3 => W_36_23_i_12_n_0,
   I4 => W_36_23_i_13_n_0,
   O => W_36_23_i_3_n_0
);
W_36_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x86_out_30,
   I1 => x86_out_5,
   I2 => x86_out_7,
   I3 => W_36_23_i_14_n_0,
   I4 => W_36_23_i_15_n_0,
   O => W_36_23_i_4_n_0
);
W_36_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x86_out_29,
   I1 => x86_out_4,
   I2 => x86_out_6,
   I3 => W_36_23_i_16_n_0,
   I4 => W_36_23_i_17_n_0,
   O => W_36_23_i_5_n_0
);
W_36_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x86_out_8,
   I1 => x86_out_10,
   I2 => W_36_27_i_16_n_0,
   I3 => W_36_27_i_17_n_0,
   I4 => W_36_23_i_2_n_0,
   O => W_36_23_i_6_n_0
);
W_36_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x86_out_7,
   I1 => x86_out_9,
   I2 => W_36_23_i_10_n_0,
   I3 => W_36_23_i_11_n_0,
   I4 => W_36_23_i_3_n_0,
   O => W_36_23_i_7_n_0
);
W_36_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_36_23_i_4_n_0,
   I1 => W_36_23_i_12_n_0,
   I2 => x86_out_31,
   I3 => x86_out_6,
   I4 => x86_out_8,
   I5 => W_36_23_i_13_n_0,
   O => W_36_23_i_8_n_0
);
W_36_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_36_23_i_5_n_0,
   I1 => W_36_23_i_14_n_0,
   I2 => x86_out_30,
   I3 => x86_out_5,
   I4 => x86_out_7,
   I5 => W_36_23_i_15_n_0,
   O => W_36_23_i_9_n_0
);
W_36_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x113_out_26,
   I1 => x98_out_26,
   I2 => x112_out_12,
   I3 => x112_out_1,
   I4 => x112_out_29,
   O => W_36_27_i_10_n_0
);
W_36_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x98_out_25,
   I1 => x112_out_28,
   I2 => x112_out_0,
   I3 => x112_out_11,
   I4 => x113_out_25,
   O => W_36_27_i_11_n_0
);
W_36_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x113_out_25,
   I1 => x98_out_25,
   I2 => x112_out_11,
   I3 => x112_out_0,
   I4 => x112_out_28,
   O => W_36_27_i_12_n_0
);
W_36_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x98_out_24,
   I1 => x112_out_27,
   I2 => x112_out_31,
   I3 => x112_out_10,
   I4 => x113_out_24,
   O => W_36_27_i_13_n_0
);
W_36_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x113_out_24,
   I1 => x98_out_24,
   I2 => x112_out_10,
   I3 => x112_out_31,
   I4 => x112_out_27,
   O => W_36_27_i_14_n_0
);
W_36_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x98_out_23,
   I1 => x112_out_26,
   I2 => x112_out_30,
   I3 => x112_out_9,
   I4 => x113_out_23,
   O => W_36_27_i_15_n_0
);
W_36_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x113_out_23,
   I1 => x98_out_23,
   I2 => x112_out_9,
   I3 => x112_out_30,
   I4 => x112_out_26,
   O => W_36_27_i_16_n_0
);
W_36_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x98_out_22,
   I1 => x112_out_25,
   I2 => x112_out_29,
   I3 => x112_out_8,
   I4 => x113_out_22,
   O => W_36_27_i_17_n_0
);
W_36_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x86_out_11,
   I1 => x86_out_13,
   I2 => W_36_27_i_10_n_0,
   I3 => W_36_27_i_11_n_0,
   O => W_36_27_i_2_n_0
);
W_36_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x86_out_10,
   I1 => x86_out_12,
   I2 => W_36_27_i_12_n_0,
   I3 => W_36_27_i_13_n_0,
   O => W_36_27_i_3_n_0
);
W_36_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x86_out_9,
   I1 => x86_out_11,
   I2 => W_36_27_i_14_n_0,
   I3 => W_36_27_i_15_n_0,
   O => W_36_27_i_4_n_0
);
W_36_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x86_out_8,
   I1 => x86_out_10,
   I2 => W_36_27_i_16_n_0,
   I3 => W_36_27_i_17_n_0,
   O => W_36_27_i_5_n_0
);
W_36_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x86_out_12,
   I1 => x86_out_14,
   I2 => W_36_31_i_13_n_0,
   I3 => W_36_31_i_14_n_0,
   I4 => W_36_27_i_2_n_0,
   O => W_36_27_i_6_n_0
);
W_36_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x86_out_11,
   I1 => x86_out_13,
   I2 => W_36_27_i_10_n_0,
   I3 => W_36_27_i_11_n_0,
   I4 => W_36_27_i_3_n_0,
   O => W_36_27_i_7_n_0
);
W_36_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x86_out_10,
   I1 => x86_out_12,
   I2 => W_36_27_i_12_n_0,
   I3 => W_36_27_i_13_n_0,
   I4 => W_36_27_i_4_n_0,
   O => W_36_27_i_8_n_0
);
W_36_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x86_out_9,
   I1 => x86_out_11,
   I2 => W_36_27_i_14_n_0,
   I3 => W_36_27_i_15_n_0,
   I4 => W_36_27_i_5_n_0,
   O => W_36_27_i_9_n_0
);
W_36_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x98_out_28,
   I1 => x112_out_31,
   I2 => x112_out_3,
   I3 => x112_out_14,
   I4 => x113_out_28,
   O => W_36_31_i_10_n_0
);
W_36_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x113_out_28,
   I1 => x98_out_28,
   I2 => x112_out_14,
   I3 => x112_out_3,
   I4 => x112_out_31,
   O => W_36_31_i_11_n_0
);
W_36_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x98_out_27,
   I1 => x112_out_30,
   I2 => x112_out_2,
   I3 => x112_out_13,
   I4 => x113_out_27,
   O => W_36_31_i_12_n_0
);
W_36_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x113_out_27,
   I1 => x98_out_27,
   I2 => x112_out_13,
   I3 => x112_out_2,
   I4 => x112_out_30,
   O => W_36_31_i_13_n_0
);
W_36_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x98_out_26,
   I1 => x112_out_29,
   I2 => x112_out_1,
   I3 => x112_out_12,
   I4 => x113_out_26,
   O => W_36_31_i_14_n_0
);
W_36_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x98_out_29,
   I1 => x112_out_4,
   I2 => x112_out_15,
   I3 => x113_out_29,
   O => W_36_31_i_15_n_0
);
W_36_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x86_out_17,
   I1 => x86_out_15,
   O => SIGMA_LCASE_1227_out_0_30
);
W_36_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => x112_out_6,
   I1 => x112_out_17,
   I2 => x98_out_31,
   I3 => x113_out_31,
   I4 => x86_out_16,
   I5 => x86_out_18,
   O => W_36_31_i_17_n_0
);
W_36_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x112_out_16,
   I1 => x112_out_5,
   O => SIGMA_LCASE_0223_out_30
);
W_36_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x113_out_30,
   I1 => x98_out_30,
   I2 => x112_out_16,
   I3 => x112_out_5,
   O => W_36_31_i_19_n_0
);
W_36_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x86_out_14,
   I1 => x86_out_16,
   I2 => W_36_31_i_9_n_0,
   I3 => W_36_31_i_10_n_0,
   O => W_36_31_i_2_n_0
);
W_36_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x86_out_13,
   I1 => x86_out_15,
   I2 => W_36_31_i_11_n_0,
   I3 => W_36_31_i_12_n_0,
   O => W_36_31_i_3_n_0
);
W_36_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x86_out_12,
   I1 => x86_out_14,
   I2 => W_36_31_i_13_n_0,
   I3 => W_36_31_i_14_n_0,
   O => W_36_31_i_4_n_0
);
W_36_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_36_31_i_15_n_0,
   I1 => SIGMA_LCASE_1227_out_0_30,
   I2 => W_36_31_i_17_n_0,
   I3 => x98_out_30,
   I4 => SIGMA_LCASE_0223_out_30,
   I5 => x113_out_30,
   O => W_36_31_i_5_n_0
);
W_36_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_36_31_i_2_n_0,
   I1 => W_36_31_i_19_n_0,
   I2 => x86_out_15,
   I3 => x86_out_17,
   I4 => W_36_31_i_15_n_0,
   O => W_36_31_i_6_n_0
);
W_36_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x86_out_14,
   I1 => x86_out_16,
   I2 => W_36_31_i_9_n_0,
   I3 => W_36_31_i_10_n_0,
   I4 => W_36_31_i_3_n_0,
   O => W_36_31_i_7_n_0
);
W_36_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x86_out_13,
   I1 => x86_out_15,
   I2 => W_36_31_i_11_n_0,
   I3 => W_36_31_i_12_n_0,
   I4 => W_36_31_i_4_n_0,
   O => W_36_31_i_8_n_0
);
W_36_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x113_out_29,
   I1 => x98_out_29,
   I2 => x112_out_15,
   I3 => x112_out_4,
   O => W_36_31_i_9_n_0
);
W_36_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x113_out_2,
   I1 => x98_out_2,
   I2 => x112_out_20,
   I3 => x112_out_9,
   I4 => x112_out_5,
   O => W_36_3_i_10_n_0
);
W_36_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x98_out_1,
   I1 => x112_out_4,
   I2 => x112_out_8,
   I3 => x112_out_19,
   I4 => x113_out_1,
   O => W_36_3_i_11_n_0
);
W_36_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x112_out_19,
   I1 => x112_out_8,
   I2 => x112_out_4,
   O => SIGMA_LCASE_0223_out_1
);
W_36_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x86_out_21,
   I1 => x86_out_19,
   I2 => x86_out_12,
   O => SIGMA_LCASE_1227_out_0_2
);
W_36_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x86_out_20,
   I1 => x86_out_18,
   I2 => x86_out_11,
   O => SIGMA_LCASE_1227_out_1
);
W_36_3_i_15 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x113_out_1,
   I1 => x98_out_1,
   I2 => x112_out_19,
   I3 => x112_out_8,
   I4 => x112_out_4,
   O => W_36_3_i_15_n_0
);
W_36_3_i_16 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x112_out_18,
   I1 => x112_out_7,
   I2 => x112_out_3,
   O => SIGMA_LCASE_0223_out_0
);
W_36_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x86_out_12,
   I1 => x86_out_19,
   I2 => x86_out_21,
   I3 => W_36_3_i_10_n_0,
   I4 => W_36_3_i_11_n_0,
   O => W_36_3_i_2_n_0
);
W_36_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_36_3_i_11_n_0,
   I1 => x86_out_21,
   I2 => x86_out_19,
   I3 => x86_out_12,
   I4 => W_36_3_i_10_n_0,
   O => W_36_3_i_3_n_0
);
W_36_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_0223_out_1,
   I1 => x98_out_1,
   I2 => x113_out_1,
   I3 => x86_out_11,
   I4 => x86_out_18,
   I5 => x86_out_20,
   O => W_36_3_i_4_n_0
);
W_36_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x113_out_0,
   I1 => x98_out_0,
   I2 => x112_out_18,
   I3 => x112_out_7,
   I4 => x112_out_3,
   O => W_36_3_i_5_n_0
);
W_36_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_36_3_i_2_n_0,
   I1 => W_36_7_i_16_n_0,
   I2 => x86_out_13,
   I3 => x86_out_20,
   I4 => x86_out_22,
   I5 => W_36_7_i_17_n_0,
   O => W_36_3_i_6_n_0
);
W_36_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_36_3_i_10_n_0,
   I1 => SIGMA_LCASE_1227_out_0_2,
   I2 => x113_out_1,
   I3 => x98_out_1,
   I4 => SIGMA_LCASE_0223_out_1,
   I5 => SIGMA_LCASE_1227_out_1,
   O => W_36_3_i_7_n_0
);
W_36_3_i_8 : LUT5
  generic map(
   INIT => X"99969666"
  )
 port map (
   I0 => SIGMA_LCASE_1227_out_1,
   I1 => W_36_3_i_15_n_0,
   I2 => x113_out_0,
   I3 => SIGMA_LCASE_0223_out_0,
   I4 => x98_out_0,
   O => W_36_3_i_8_n_0
);
W_36_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_36_3_i_5_n_0,
   I1 => x86_out_10,
   I2 => x86_out_17,
   I3 => x86_out_19,
   O => W_36_3_i_9_n_0
);
W_36_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x113_out_6,
   I1 => x98_out_6,
   I2 => x112_out_24,
   I3 => x112_out_13,
   I4 => x112_out_9,
   O => W_36_7_i_10_n_0
);
W_36_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x98_out_5,
   I1 => x112_out_8,
   I2 => x112_out_12,
   I3 => x112_out_23,
   I4 => x113_out_5,
   O => W_36_7_i_11_n_0
);
W_36_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x113_out_5,
   I1 => x98_out_5,
   I2 => x112_out_23,
   I3 => x112_out_12,
   I4 => x112_out_8,
   O => W_36_7_i_12_n_0
);
W_36_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x98_out_4,
   I1 => x112_out_7,
   I2 => x112_out_11,
   I3 => x112_out_22,
   I4 => x113_out_4,
   O => W_36_7_i_13_n_0
);
W_36_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x113_out_4,
   I1 => x98_out_4,
   I2 => x112_out_22,
   I3 => x112_out_11,
   I4 => x112_out_7,
   O => W_36_7_i_14_n_0
);
W_36_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x98_out_3,
   I1 => x112_out_6,
   I2 => x112_out_10,
   I3 => x112_out_21,
   I4 => x113_out_3,
   O => W_36_7_i_15_n_0
);
W_36_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x113_out_3,
   I1 => x98_out_3,
   I2 => x112_out_21,
   I3 => x112_out_10,
   I4 => x112_out_6,
   O => W_36_7_i_16_n_0
);
W_36_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x98_out_2,
   I1 => x112_out_5,
   I2 => x112_out_9,
   I3 => x112_out_20,
   I4 => x113_out_2,
   O => W_36_7_i_17_n_0
);
W_36_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x86_out_16,
   I1 => x86_out_23,
   I2 => x86_out_25,
   I3 => W_36_7_i_10_n_0,
   I4 => W_36_7_i_11_n_0,
   O => W_36_7_i_2_n_0
);
W_36_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x86_out_15,
   I1 => x86_out_22,
   I2 => x86_out_24,
   I3 => W_36_7_i_12_n_0,
   I4 => W_36_7_i_13_n_0,
   O => W_36_7_i_3_n_0
);
W_36_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x86_out_14,
   I1 => x86_out_21,
   I2 => x86_out_23,
   I3 => W_36_7_i_14_n_0,
   I4 => W_36_7_i_15_n_0,
   O => W_36_7_i_4_n_0
);
W_36_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x86_out_13,
   I1 => x86_out_20,
   I2 => x86_out_22,
   I3 => W_36_7_i_16_n_0,
   I4 => W_36_7_i_17_n_0,
   O => W_36_7_i_5_n_0
);
W_36_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_36_7_i_2_n_0,
   I1 => W_36_11_i_16_n_0,
   I2 => x86_out_17,
   I3 => x86_out_24,
   I4 => x86_out_26,
   I5 => W_36_11_i_17_n_0,
   O => W_36_7_i_6_n_0
);
W_36_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_36_7_i_3_n_0,
   I1 => W_36_7_i_10_n_0,
   I2 => x86_out_16,
   I3 => x86_out_23,
   I4 => x86_out_25,
   I5 => W_36_7_i_11_n_0,
   O => W_36_7_i_7_n_0
);
W_36_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_36_7_i_4_n_0,
   I1 => W_36_7_i_12_n_0,
   I2 => x86_out_15,
   I3 => x86_out_22,
   I4 => x86_out_24,
   I5 => W_36_7_i_13_n_0,
   O => W_36_7_i_8_n_0
);
W_36_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_36_7_i_5_n_0,
   I1 => W_36_7_i_14_n_0,
   I2 => x86_out_14,
   I3 => x86_out_21,
   I4 => x86_out_23,
   I5 => W_36_7_i_15_n_0,
   O => W_36_7_i_9_n_0
);
W_37_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x112_out_10,
   I1 => x96_out_10,
   I2 => x111_out_28,
   I3 => x111_out_17,
   I4 => x111_out_13,
   O => W_37_11_i_10_n_0
);
W_37_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x96_out_9,
   I1 => x111_out_12,
   I2 => x111_out_16,
   I3 => x111_out_27,
   I4 => x112_out_9,
   O => W_37_11_i_11_n_0
);
W_37_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x112_out_9,
   I1 => x96_out_9,
   I2 => x111_out_27,
   I3 => x111_out_16,
   I4 => x111_out_12,
   O => W_37_11_i_12_n_0
);
W_37_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x96_out_8,
   I1 => x111_out_11,
   I2 => x111_out_15,
   I3 => x111_out_26,
   I4 => x112_out_8,
   O => W_37_11_i_13_n_0
);
W_37_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x112_out_8,
   I1 => x96_out_8,
   I2 => x111_out_26,
   I3 => x111_out_15,
   I4 => x111_out_11,
   O => W_37_11_i_14_n_0
);
W_37_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x96_out_7,
   I1 => x111_out_10,
   I2 => x111_out_14,
   I3 => x111_out_25,
   I4 => x112_out_7,
   O => W_37_11_i_15_n_0
);
W_37_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x112_out_7,
   I1 => x96_out_7,
   I2 => x111_out_25,
   I3 => x111_out_14,
   I4 => x111_out_10,
   O => W_37_11_i_16_n_0
);
W_37_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x96_out_6,
   I1 => x111_out_9,
   I2 => x111_out_13,
   I3 => x111_out_24,
   I4 => x112_out_6,
   O => W_37_11_i_17_n_0
);
W_37_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x83_out_20,
   I1 => x83_out_27,
   I2 => x83_out_29,
   I3 => W_37_11_i_10_n_0,
   I4 => W_37_11_i_11_n_0,
   O => W_37_11_i_2_n_0
);
W_37_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x83_out_19,
   I1 => x83_out_26,
   I2 => x83_out_28,
   I3 => W_37_11_i_12_n_0,
   I4 => W_37_11_i_13_n_0,
   O => W_37_11_i_3_n_0
);
W_37_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x83_out_18,
   I1 => x83_out_25,
   I2 => x83_out_27,
   I3 => W_37_11_i_14_n_0,
   I4 => W_37_11_i_15_n_0,
   O => W_37_11_i_4_n_0
);
W_37_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x83_out_17,
   I1 => x83_out_24,
   I2 => x83_out_26,
   I3 => W_37_11_i_16_n_0,
   I4 => W_37_11_i_17_n_0,
   O => W_37_11_i_5_n_0
);
W_37_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_37_11_i_2_n_0,
   I1 => W_37_15_i_16_n_0,
   I2 => x83_out_21,
   I3 => x83_out_28,
   I4 => x83_out_30,
   I5 => W_37_15_i_17_n_0,
   O => W_37_11_i_6_n_0
);
W_37_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_37_11_i_3_n_0,
   I1 => W_37_11_i_10_n_0,
   I2 => x83_out_20,
   I3 => x83_out_27,
   I4 => x83_out_29,
   I5 => W_37_11_i_11_n_0,
   O => W_37_11_i_7_n_0
);
W_37_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_37_11_i_4_n_0,
   I1 => W_37_11_i_12_n_0,
   I2 => x83_out_19,
   I3 => x83_out_26,
   I4 => x83_out_28,
   I5 => W_37_11_i_13_n_0,
   O => W_37_11_i_8_n_0
);
W_37_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_37_11_i_5_n_0,
   I1 => W_37_11_i_14_n_0,
   I2 => x83_out_18,
   I3 => x83_out_25,
   I4 => x83_out_27,
   I5 => W_37_11_i_15_n_0,
   O => W_37_11_i_9_n_0
);
W_37_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x112_out_14,
   I1 => x96_out_14,
   I2 => x111_out_0,
   I3 => x111_out_21,
   I4 => x111_out_17,
   O => W_37_15_i_10_n_0
);
W_37_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x96_out_13,
   I1 => x111_out_16,
   I2 => x111_out_20,
   I3 => x111_out_31,
   I4 => x112_out_13,
   O => W_37_15_i_11_n_0
);
W_37_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x112_out_13,
   I1 => x96_out_13,
   I2 => x111_out_31,
   I3 => x111_out_20,
   I4 => x111_out_16,
   O => W_37_15_i_12_n_0
);
W_37_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x96_out_12,
   I1 => x111_out_15,
   I2 => x111_out_19,
   I3 => x111_out_30,
   I4 => x112_out_12,
   O => W_37_15_i_13_n_0
);
W_37_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x112_out_12,
   I1 => x96_out_12,
   I2 => x111_out_30,
   I3 => x111_out_19,
   I4 => x111_out_15,
   O => W_37_15_i_14_n_0
);
W_37_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x96_out_11,
   I1 => x111_out_14,
   I2 => x111_out_18,
   I3 => x111_out_29,
   I4 => x112_out_11,
   O => W_37_15_i_15_n_0
);
W_37_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x112_out_11,
   I1 => x96_out_11,
   I2 => x111_out_29,
   I3 => x111_out_18,
   I4 => x111_out_14,
   O => W_37_15_i_16_n_0
);
W_37_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x96_out_10,
   I1 => x111_out_13,
   I2 => x111_out_17,
   I3 => x111_out_28,
   I4 => x112_out_10,
   O => W_37_15_i_17_n_0
);
W_37_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x83_out_24,
   I1 => x83_out_31,
   I2 => x83_out_1,
   I3 => W_37_15_i_10_n_0,
   I4 => W_37_15_i_11_n_0,
   O => W_37_15_i_2_n_0
);
W_37_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x83_out_23,
   I1 => x83_out_30,
   I2 => x83_out_0,
   I3 => W_37_15_i_12_n_0,
   I4 => W_37_15_i_13_n_0,
   O => W_37_15_i_3_n_0
);
W_37_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x83_out_22,
   I1 => x83_out_29,
   I2 => x83_out_31,
   I3 => W_37_15_i_14_n_0,
   I4 => W_37_15_i_15_n_0,
   O => W_37_15_i_4_n_0
);
W_37_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x83_out_21,
   I1 => x83_out_28,
   I2 => x83_out_30,
   I3 => W_37_15_i_16_n_0,
   I4 => W_37_15_i_17_n_0,
   O => W_37_15_i_5_n_0
);
W_37_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_37_15_i_2_n_0,
   I1 => W_37_19_i_16_n_0,
   I2 => x83_out_25,
   I3 => x83_out_0,
   I4 => x83_out_2,
   I5 => W_37_19_i_17_n_0,
   O => W_37_15_i_6_n_0
);
W_37_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_37_15_i_3_n_0,
   I1 => W_37_15_i_10_n_0,
   I2 => x83_out_24,
   I3 => x83_out_31,
   I4 => x83_out_1,
   I5 => W_37_15_i_11_n_0,
   O => W_37_15_i_7_n_0
);
W_37_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_37_15_i_4_n_0,
   I1 => W_37_15_i_12_n_0,
   I2 => x83_out_23,
   I3 => x83_out_30,
   I4 => x83_out_0,
   I5 => W_37_15_i_13_n_0,
   O => W_37_15_i_8_n_0
);
W_37_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_37_15_i_5_n_0,
   I1 => W_37_15_i_14_n_0,
   I2 => x83_out_22,
   I3 => x83_out_29,
   I4 => x83_out_31,
   I5 => W_37_15_i_15_n_0,
   O => W_37_15_i_9_n_0
);
W_37_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x112_out_18,
   I1 => x96_out_18,
   I2 => x111_out_4,
   I3 => x111_out_25,
   I4 => x111_out_21,
   O => W_37_19_i_10_n_0
);
W_37_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x96_out_17,
   I1 => x111_out_20,
   I2 => x111_out_24,
   I3 => x111_out_3,
   I4 => x112_out_17,
   O => W_37_19_i_11_n_0
);
W_37_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x112_out_17,
   I1 => x96_out_17,
   I2 => x111_out_3,
   I3 => x111_out_24,
   I4 => x111_out_20,
   O => W_37_19_i_12_n_0
);
W_37_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x96_out_16,
   I1 => x111_out_19,
   I2 => x111_out_23,
   I3 => x111_out_2,
   I4 => x112_out_16,
   O => W_37_19_i_13_n_0
);
W_37_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x112_out_16,
   I1 => x96_out_16,
   I2 => x111_out_2,
   I3 => x111_out_23,
   I4 => x111_out_19,
   O => W_37_19_i_14_n_0
);
W_37_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x96_out_15,
   I1 => x111_out_18,
   I2 => x111_out_22,
   I3 => x111_out_1,
   I4 => x112_out_15,
   O => W_37_19_i_15_n_0
);
W_37_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x112_out_15,
   I1 => x96_out_15,
   I2 => x111_out_1,
   I3 => x111_out_22,
   I4 => x111_out_18,
   O => W_37_19_i_16_n_0
);
W_37_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x96_out_14,
   I1 => x111_out_17,
   I2 => x111_out_21,
   I3 => x111_out_0,
   I4 => x112_out_14,
   O => W_37_19_i_17_n_0
);
W_37_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x83_out_28,
   I1 => x83_out_3,
   I2 => x83_out_5,
   I3 => W_37_19_i_10_n_0,
   I4 => W_37_19_i_11_n_0,
   O => W_37_19_i_2_n_0
);
W_37_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x83_out_27,
   I1 => x83_out_2,
   I2 => x83_out_4,
   I3 => W_37_19_i_12_n_0,
   I4 => W_37_19_i_13_n_0,
   O => W_37_19_i_3_n_0
);
W_37_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x83_out_26,
   I1 => x83_out_1,
   I2 => x83_out_3,
   I3 => W_37_19_i_14_n_0,
   I4 => W_37_19_i_15_n_0,
   O => W_37_19_i_4_n_0
);
W_37_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x83_out_25,
   I1 => x83_out_0,
   I2 => x83_out_2,
   I3 => W_37_19_i_16_n_0,
   I4 => W_37_19_i_17_n_0,
   O => W_37_19_i_5_n_0
);
W_37_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_37_19_i_2_n_0,
   I1 => W_37_23_i_16_n_0,
   I2 => x83_out_29,
   I3 => x83_out_4,
   I4 => x83_out_6,
   I5 => W_37_23_i_17_n_0,
   O => W_37_19_i_6_n_0
);
W_37_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_37_19_i_3_n_0,
   I1 => W_37_19_i_10_n_0,
   I2 => x83_out_28,
   I3 => x83_out_3,
   I4 => x83_out_5,
   I5 => W_37_19_i_11_n_0,
   O => W_37_19_i_7_n_0
);
W_37_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_37_19_i_4_n_0,
   I1 => W_37_19_i_12_n_0,
   I2 => x83_out_27,
   I3 => x83_out_2,
   I4 => x83_out_4,
   I5 => W_37_19_i_13_n_0,
   O => W_37_19_i_8_n_0
);
W_37_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_37_19_i_5_n_0,
   I1 => W_37_19_i_14_n_0,
   I2 => x83_out_26,
   I3 => x83_out_1,
   I4 => x83_out_3,
   I5 => W_37_19_i_15_n_0,
   O => W_37_19_i_9_n_0
);
W_37_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x112_out_22,
   I1 => x96_out_22,
   I2 => x111_out_8,
   I3 => x111_out_29,
   I4 => x111_out_25,
   O => W_37_23_i_10_n_0
);
W_37_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x96_out_21,
   I1 => x111_out_24,
   I2 => x111_out_28,
   I3 => x111_out_7,
   I4 => x112_out_21,
   O => W_37_23_i_11_n_0
);
W_37_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x112_out_21,
   I1 => x96_out_21,
   I2 => x111_out_7,
   I3 => x111_out_28,
   I4 => x111_out_24,
   O => W_37_23_i_12_n_0
);
W_37_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x96_out_20,
   I1 => x111_out_23,
   I2 => x111_out_27,
   I3 => x111_out_6,
   I4 => x112_out_20,
   O => W_37_23_i_13_n_0
);
W_37_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x112_out_20,
   I1 => x96_out_20,
   I2 => x111_out_6,
   I3 => x111_out_27,
   I4 => x111_out_23,
   O => W_37_23_i_14_n_0
);
W_37_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x96_out_19,
   I1 => x111_out_22,
   I2 => x111_out_26,
   I3 => x111_out_5,
   I4 => x112_out_19,
   O => W_37_23_i_15_n_0
);
W_37_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x112_out_19,
   I1 => x96_out_19,
   I2 => x111_out_5,
   I3 => x111_out_26,
   I4 => x111_out_22,
   O => W_37_23_i_16_n_0
);
W_37_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x96_out_18,
   I1 => x111_out_21,
   I2 => x111_out_25,
   I3 => x111_out_4,
   I4 => x112_out_18,
   O => W_37_23_i_17_n_0
);
W_37_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x83_out_7,
   I1 => x83_out_9,
   I2 => W_37_23_i_10_n_0,
   I3 => W_37_23_i_11_n_0,
   O => W_37_23_i_2_n_0
);
W_37_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x83_out_31,
   I1 => x83_out_6,
   I2 => x83_out_8,
   I3 => W_37_23_i_12_n_0,
   I4 => W_37_23_i_13_n_0,
   O => W_37_23_i_3_n_0
);
W_37_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x83_out_30,
   I1 => x83_out_5,
   I2 => x83_out_7,
   I3 => W_37_23_i_14_n_0,
   I4 => W_37_23_i_15_n_0,
   O => W_37_23_i_4_n_0
);
W_37_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x83_out_29,
   I1 => x83_out_4,
   I2 => x83_out_6,
   I3 => W_37_23_i_16_n_0,
   I4 => W_37_23_i_17_n_0,
   O => W_37_23_i_5_n_0
);
W_37_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x83_out_8,
   I1 => x83_out_10,
   I2 => W_37_27_i_16_n_0,
   I3 => W_37_27_i_17_n_0,
   I4 => W_37_23_i_2_n_0,
   O => W_37_23_i_6_n_0
);
W_37_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x83_out_7,
   I1 => x83_out_9,
   I2 => W_37_23_i_10_n_0,
   I3 => W_37_23_i_11_n_0,
   I4 => W_37_23_i_3_n_0,
   O => W_37_23_i_7_n_0
);
W_37_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_37_23_i_4_n_0,
   I1 => W_37_23_i_12_n_0,
   I2 => x83_out_31,
   I3 => x83_out_6,
   I4 => x83_out_8,
   I5 => W_37_23_i_13_n_0,
   O => W_37_23_i_8_n_0
);
W_37_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_37_23_i_5_n_0,
   I1 => W_37_23_i_14_n_0,
   I2 => x83_out_30,
   I3 => x83_out_5,
   I4 => x83_out_7,
   I5 => W_37_23_i_15_n_0,
   O => W_37_23_i_9_n_0
);
W_37_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x112_out_26,
   I1 => x96_out_26,
   I2 => x111_out_12,
   I3 => x111_out_1,
   I4 => x111_out_29,
   O => W_37_27_i_10_n_0
);
W_37_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x96_out_25,
   I1 => x111_out_28,
   I2 => x111_out_0,
   I3 => x111_out_11,
   I4 => x112_out_25,
   O => W_37_27_i_11_n_0
);
W_37_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x112_out_25,
   I1 => x96_out_25,
   I2 => x111_out_11,
   I3 => x111_out_0,
   I4 => x111_out_28,
   O => W_37_27_i_12_n_0
);
W_37_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x96_out_24,
   I1 => x111_out_27,
   I2 => x111_out_31,
   I3 => x111_out_10,
   I4 => x112_out_24,
   O => W_37_27_i_13_n_0
);
W_37_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x112_out_24,
   I1 => x96_out_24,
   I2 => x111_out_10,
   I3 => x111_out_31,
   I4 => x111_out_27,
   O => W_37_27_i_14_n_0
);
W_37_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x96_out_23,
   I1 => x111_out_26,
   I2 => x111_out_30,
   I3 => x111_out_9,
   I4 => x112_out_23,
   O => W_37_27_i_15_n_0
);
W_37_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x112_out_23,
   I1 => x96_out_23,
   I2 => x111_out_9,
   I3 => x111_out_30,
   I4 => x111_out_26,
   O => W_37_27_i_16_n_0
);
W_37_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x96_out_22,
   I1 => x111_out_25,
   I2 => x111_out_29,
   I3 => x111_out_8,
   I4 => x112_out_22,
   O => W_37_27_i_17_n_0
);
W_37_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x83_out_11,
   I1 => x83_out_13,
   I2 => W_37_27_i_10_n_0,
   I3 => W_37_27_i_11_n_0,
   O => W_37_27_i_2_n_0
);
W_37_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x83_out_10,
   I1 => x83_out_12,
   I2 => W_37_27_i_12_n_0,
   I3 => W_37_27_i_13_n_0,
   O => W_37_27_i_3_n_0
);
W_37_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x83_out_9,
   I1 => x83_out_11,
   I2 => W_37_27_i_14_n_0,
   I3 => W_37_27_i_15_n_0,
   O => W_37_27_i_4_n_0
);
W_37_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x83_out_8,
   I1 => x83_out_10,
   I2 => W_37_27_i_16_n_0,
   I3 => W_37_27_i_17_n_0,
   O => W_37_27_i_5_n_0
);
W_37_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x83_out_12,
   I1 => x83_out_14,
   I2 => W_37_31_i_13_n_0,
   I3 => W_37_31_i_14_n_0,
   I4 => W_37_27_i_2_n_0,
   O => W_37_27_i_6_n_0
);
W_37_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x83_out_11,
   I1 => x83_out_13,
   I2 => W_37_27_i_10_n_0,
   I3 => W_37_27_i_11_n_0,
   I4 => W_37_27_i_3_n_0,
   O => W_37_27_i_7_n_0
);
W_37_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x83_out_10,
   I1 => x83_out_12,
   I2 => W_37_27_i_12_n_0,
   I3 => W_37_27_i_13_n_0,
   I4 => W_37_27_i_4_n_0,
   O => W_37_27_i_8_n_0
);
W_37_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x83_out_9,
   I1 => x83_out_11,
   I2 => W_37_27_i_14_n_0,
   I3 => W_37_27_i_15_n_0,
   I4 => W_37_27_i_5_n_0,
   O => W_37_27_i_9_n_0
);
W_37_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x96_out_28,
   I1 => x111_out_31,
   I2 => x111_out_3,
   I3 => x111_out_14,
   I4 => x112_out_28,
   O => W_37_31_i_10_n_0
);
W_37_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x112_out_28,
   I1 => x96_out_28,
   I2 => x111_out_14,
   I3 => x111_out_3,
   I4 => x111_out_31,
   O => W_37_31_i_11_n_0
);
W_37_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x96_out_27,
   I1 => x111_out_30,
   I2 => x111_out_2,
   I3 => x111_out_13,
   I4 => x112_out_27,
   O => W_37_31_i_12_n_0
);
W_37_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x112_out_27,
   I1 => x96_out_27,
   I2 => x111_out_13,
   I3 => x111_out_2,
   I4 => x111_out_30,
   O => W_37_31_i_13_n_0
);
W_37_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x96_out_26,
   I1 => x111_out_29,
   I2 => x111_out_1,
   I3 => x111_out_12,
   I4 => x112_out_26,
   O => W_37_31_i_14_n_0
);
W_37_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x96_out_29,
   I1 => x111_out_4,
   I2 => x111_out_15,
   I3 => x112_out_29,
   O => W_37_31_i_15_n_0
);
W_37_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x83_out_17,
   I1 => x83_out_15,
   O => SIGMA_LCASE_1219_out_0_30
);
W_37_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => x111_out_6,
   I1 => x111_out_17,
   I2 => x96_out_31,
   I3 => x112_out_31,
   I4 => x83_out_16,
   I5 => x83_out_18,
   O => W_37_31_i_17_n_0
);
W_37_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x111_out_16,
   I1 => x111_out_5,
   O => SIGMA_LCASE_0215_out_30
);
W_37_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x112_out_30,
   I1 => x96_out_30,
   I2 => x111_out_16,
   I3 => x111_out_5,
   O => W_37_31_i_19_n_0
);
W_37_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x83_out_14,
   I1 => x83_out_16,
   I2 => W_37_31_i_9_n_0,
   I3 => W_37_31_i_10_n_0,
   O => W_37_31_i_2_n_0
);
W_37_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x83_out_13,
   I1 => x83_out_15,
   I2 => W_37_31_i_11_n_0,
   I3 => W_37_31_i_12_n_0,
   O => W_37_31_i_3_n_0
);
W_37_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x83_out_12,
   I1 => x83_out_14,
   I2 => W_37_31_i_13_n_0,
   I3 => W_37_31_i_14_n_0,
   O => W_37_31_i_4_n_0
);
W_37_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_37_31_i_15_n_0,
   I1 => SIGMA_LCASE_1219_out_0_30,
   I2 => W_37_31_i_17_n_0,
   I3 => x96_out_30,
   I4 => SIGMA_LCASE_0215_out_30,
   I5 => x112_out_30,
   O => W_37_31_i_5_n_0
);
W_37_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_37_31_i_2_n_0,
   I1 => W_37_31_i_19_n_0,
   I2 => x83_out_15,
   I3 => x83_out_17,
   I4 => W_37_31_i_15_n_0,
   O => W_37_31_i_6_n_0
);
W_37_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x83_out_14,
   I1 => x83_out_16,
   I2 => W_37_31_i_9_n_0,
   I3 => W_37_31_i_10_n_0,
   I4 => W_37_31_i_3_n_0,
   O => W_37_31_i_7_n_0
);
W_37_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x83_out_13,
   I1 => x83_out_15,
   I2 => W_37_31_i_11_n_0,
   I3 => W_37_31_i_12_n_0,
   I4 => W_37_31_i_4_n_0,
   O => W_37_31_i_8_n_0
);
W_37_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x112_out_29,
   I1 => x96_out_29,
   I2 => x111_out_15,
   I3 => x111_out_4,
   O => W_37_31_i_9_n_0
);
W_37_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x112_out_2,
   I1 => x96_out_2,
   I2 => x111_out_20,
   I3 => x111_out_9,
   I4 => x111_out_5,
   O => W_37_3_i_10_n_0
);
W_37_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x96_out_1,
   I1 => x111_out_4,
   I2 => x111_out_8,
   I3 => x111_out_19,
   I4 => x112_out_1,
   O => W_37_3_i_11_n_0
);
W_37_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x111_out_19,
   I1 => x111_out_8,
   I2 => x111_out_4,
   O => SIGMA_LCASE_0215_out_1
);
W_37_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x83_out_21,
   I1 => x83_out_19,
   I2 => x83_out_12,
   O => SIGMA_LCASE_1219_out_0_2
);
W_37_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x83_out_20,
   I1 => x83_out_18,
   I2 => x83_out_11,
   O => SIGMA_LCASE_1219_out_1
);
W_37_3_i_15 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x112_out_1,
   I1 => x96_out_1,
   I2 => x111_out_19,
   I3 => x111_out_8,
   I4 => x111_out_4,
   O => W_37_3_i_15_n_0
);
W_37_3_i_16 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x111_out_18,
   I1 => x111_out_7,
   I2 => x111_out_3,
   O => SIGMA_LCASE_0215_out_0
);
W_37_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x83_out_12,
   I1 => x83_out_19,
   I2 => x83_out_21,
   I3 => W_37_3_i_10_n_0,
   I4 => W_37_3_i_11_n_0,
   O => W_37_3_i_2_n_0
);
W_37_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_37_3_i_11_n_0,
   I1 => x83_out_21,
   I2 => x83_out_19,
   I3 => x83_out_12,
   I4 => W_37_3_i_10_n_0,
   O => W_37_3_i_3_n_0
);
W_37_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_0215_out_1,
   I1 => x96_out_1,
   I2 => x112_out_1,
   I3 => x83_out_11,
   I4 => x83_out_18,
   I5 => x83_out_20,
   O => W_37_3_i_4_n_0
);
W_37_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x112_out_0,
   I1 => x96_out_0,
   I2 => x111_out_18,
   I3 => x111_out_7,
   I4 => x111_out_3,
   O => W_37_3_i_5_n_0
);
W_37_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_37_3_i_2_n_0,
   I1 => W_37_7_i_16_n_0,
   I2 => x83_out_13,
   I3 => x83_out_20,
   I4 => x83_out_22,
   I5 => W_37_7_i_17_n_0,
   O => W_37_3_i_6_n_0
);
W_37_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_37_3_i_10_n_0,
   I1 => SIGMA_LCASE_1219_out_0_2,
   I2 => x112_out_1,
   I3 => x96_out_1,
   I4 => SIGMA_LCASE_0215_out_1,
   I5 => SIGMA_LCASE_1219_out_1,
   O => W_37_3_i_7_n_0
);
W_37_3_i_8 : LUT5
  generic map(
   INIT => X"99969666"
  )
 port map (
   I0 => SIGMA_LCASE_1219_out_1,
   I1 => W_37_3_i_15_n_0,
   I2 => x112_out_0,
   I3 => SIGMA_LCASE_0215_out_0,
   I4 => x96_out_0,
   O => W_37_3_i_8_n_0
);
W_37_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_37_3_i_5_n_0,
   I1 => x83_out_10,
   I2 => x83_out_17,
   I3 => x83_out_19,
   O => W_37_3_i_9_n_0
);
W_37_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x112_out_6,
   I1 => x96_out_6,
   I2 => x111_out_24,
   I3 => x111_out_13,
   I4 => x111_out_9,
   O => W_37_7_i_10_n_0
);
W_37_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x96_out_5,
   I1 => x111_out_8,
   I2 => x111_out_12,
   I3 => x111_out_23,
   I4 => x112_out_5,
   O => W_37_7_i_11_n_0
);
W_37_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x112_out_5,
   I1 => x96_out_5,
   I2 => x111_out_23,
   I3 => x111_out_12,
   I4 => x111_out_8,
   O => W_37_7_i_12_n_0
);
W_37_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x96_out_4,
   I1 => x111_out_7,
   I2 => x111_out_11,
   I3 => x111_out_22,
   I4 => x112_out_4,
   O => W_37_7_i_13_n_0
);
W_37_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x112_out_4,
   I1 => x96_out_4,
   I2 => x111_out_22,
   I3 => x111_out_11,
   I4 => x111_out_7,
   O => W_37_7_i_14_n_0
);
W_37_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x96_out_3,
   I1 => x111_out_6,
   I2 => x111_out_10,
   I3 => x111_out_21,
   I4 => x112_out_3,
   O => W_37_7_i_15_n_0
);
W_37_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x112_out_3,
   I1 => x96_out_3,
   I2 => x111_out_21,
   I3 => x111_out_10,
   I4 => x111_out_6,
   O => W_37_7_i_16_n_0
);
W_37_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x96_out_2,
   I1 => x111_out_5,
   I2 => x111_out_9,
   I3 => x111_out_20,
   I4 => x112_out_2,
   O => W_37_7_i_17_n_0
);
W_37_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x83_out_16,
   I1 => x83_out_23,
   I2 => x83_out_25,
   I3 => W_37_7_i_10_n_0,
   I4 => W_37_7_i_11_n_0,
   O => W_37_7_i_2_n_0
);
W_37_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x83_out_15,
   I1 => x83_out_22,
   I2 => x83_out_24,
   I3 => W_37_7_i_12_n_0,
   I4 => W_37_7_i_13_n_0,
   O => W_37_7_i_3_n_0
);
W_37_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x83_out_14,
   I1 => x83_out_21,
   I2 => x83_out_23,
   I3 => W_37_7_i_14_n_0,
   I4 => W_37_7_i_15_n_0,
   O => W_37_7_i_4_n_0
);
W_37_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x83_out_13,
   I1 => x83_out_20,
   I2 => x83_out_22,
   I3 => W_37_7_i_16_n_0,
   I4 => W_37_7_i_17_n_0,
   O => W_37_7_i_5_n_0
);
W_37_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_37_7_i_2_n_0,
   I1 => W_37_11_i_16_n_0,
   I2 => x83_out_17,
   I3 => x83_out_24,
   I4 => x83_out_26,
   I5 => W_37_11_i_17_n_0,
   O => W_37_7_i_6_n_0
);
W_37_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_37_7_i_3_n_0,
   I1 => W_37_7_i_10_n_0,
   I2 => x83_out_16,
   I3 => x83_out_23,
   I4 => x83_out_25,
   I5 => W_37_7_i_11_n_0,
   O => W_37_7_i_7_n_0
);
W_37_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_37_7_i_4_n_0,
   I1 => W_37_7_i_12_n_0,
   I2 => x83_out_15,
   I3 => x83_out_22,
   I4 => x83_out_24,
   I5 => W_37_7_i_13_n_0,
   O => W_37_7_i_8_n_0
);
W_37_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_37_7_i_5_n_0,
   I1 => W_37_7_i_14_n_0,
   I2 => x83_out_14,
   I3 => x83_out_21,
   I4 => x83_out_23,
   I5 => W_37_7_i_15_n_0,
   O => W_37_7_i_9_n_0
);
W_38_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x111_out_10,
   I1 => x94_out_10,
   I2 => x110_out_28,
   I3 => x110_out_17,
   I4 => x110_out_13,
   O => W_38_11_i_10_n_0
);
W_38_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x94_out_9,
   I1 => x110_out_12,
   I2 => x110_out_16,
   I3 => x110_out_27,
   I4 => x111_out_9,
   O => W_38_11_i_11_n_0
);
W_38_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x111_out_9,
   I1 => x94_out_9,
   I2 => x110_out_27,
   I3 => x110_out_16,
   I4 => x110_out_12,
   O => W_38_11_i_12_n_0
);
W_38_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x94_out_8,
   I1 => x110_out_11,
   I2 => x110_out_15,
   I3 => x110_out_26,
   I4 => x111_out_8,
   O => W_38_11_i_13_n_0
);
W_38_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x111_out_8,
   I1 => x94_out_8,
   I2 => x110_out_26,
   I3 => x110_out_15,
   I4 => x110_out_11,
   O => W_38_11_i_14_n_0
);
W_38_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x94_out_7,
   I1 => x110_out_10,
   I2 => x110_out_14,
   I3 => x110_out_25,
   I4 => x111_out_7,
   O => W_38_11_i_15_n_0
);
W_38_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x111_out_7,
   I1 => x94_out_7,
   I2 => x110_out_25,
   I3 => x110_out_14,
   I4 => x110_out_10,
   O => W_38_11_i_16_n_0
);
W_38_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x94_out_6,
   I1 => x110_out_9,
   I2 => x110_out_13,
   I3 => x110_out_24,
   I4 => x111_out_6,
   O => W_38_11_i_17_n_0
);
W_38_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x80_out_20,
   I1 => x80_out_27,
   I2 => x80_out_29,
   I3 => W_38_11_i_10_n_0,
   I4 => W_38_11_i_11_n_0,
   O => W_38_11_i_2_n_0
);
W_38_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x80_out_19,
   I1 => x80_out_26,
   I2 => x80_out_28,
   I3 => W_38_11_i_12_n_0,
   I4 => W_38_11_i_13_n_0,
   O => W_38_11_i_3_n_0
);
W_38_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x80_out_18,
   I1 => x80_out_25,
   I2 => x80_out_27,
   I3 => W_38_11_i_14_n_0,
   I4 => W_38_11_i_15_n_0,
   O => W_38_11_i_4_n_0
);
W_38_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x80_out_17,
   I1 => x80_out_24,
   I2 => x80_out_26,
   I3 => W_38_11_i_16_n_0,
   I4 => W_38_11_i_17_n_0,
   O => W_38_11_i_5_n_0
);
W_38_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_38_11_i_2_n_0,
   I1 => W_38_15_i_16_n_0,
   I2 => x80_out_21,
   I3 => x80_out_28,
   I4 => x80_out_30,
   I5 => W_38_15_i_17_n_0,
   O => W_38_11_i_6_n_0
);
W_38_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_38_11_i_3_n_0,
   I1 => W_38_11_i_10_n_0,
   I2 => x80_out_20,
   I3 => x80_out_27,
   I4 => x80_out_29,
   I5 => W_38_11_i_11_n_0,
   O => W_38_11_i_7_n_0
);
W_38_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_38_11_i_4_n_0,
   I1 => W_38_11_i_12_n_0,
   I2 => x80_out_19,
   I3 => x80_out_26,
   I4 => x80_out_28,
   I5 => W_38_11_i_13_n_0,
   O => W_38_11_i_8_n_0
);
W_38_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_38_11_i_5_n_0,
   I1 => W_38_11_i_14_n_0,
   I2 => x80_out_18,
   I3 => x80_out_25,
   I4 => x80_out_27,
   I5 => W_38_11_i_15_n_0,
   O => W_38_11_i_9_n_0
);
W_38_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x111_out_14,
   I1 => x94_out_14,
   I2 => x110_out_0,
   I3 => x110_out_21,
   I4 => x110_out_17,
   O => W_38_15_i_10_n_0
);
W_38_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x94_out_13,
   I1 => x110_out_16,
   I2 => x110_out_20,
   I3 => x110_out_31,
   I4 => x111_out_13,
   O => W_38_15_i_11_n_0
);
W_38_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x111_out_13,
   I1 => x94_out_13,
   I2 => x110_out_31,
   I3 => x110_out_20,
   I4 => x110_out_16,
   O => W_38_15_i_12_n_0
);
W_38_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x94_out_12,
   I1 => x110_out_15,
   I2 => x110_out_19,
   I3 => x110_out_30,
   I4 => x111_out_12,
   O => W_38_15_i_13_n_0
);
W_38_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x111_out_12,
   I1 => x94_out_12,
   I2 => x110_out_30,
   I3 => x110_out_19,
   I4 => x110_out_15,
   O => W_38_15_i_14_n_0
);
W_38_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x94_out_11,
   I1 => x110_out_14,
   I2 => x110_out_18,
   I3 => x110_out_29,
   I4 => x111_out_11,
   O => W_38_15_i_15_n_0
);
W_38_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x111_out_11,
   I1 => x94_out_11,
   I2 => x110_out_29,
   I3 => x110_out_18,
   I4 => x110_out_14,
   O => W_38_15_i_16_n_0
);
W_38_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x94_out_10,
   I1 => x110_out_13,
   I2 => x110_out_17,
   I3 => x110_out_28,
   I4 => x111_out_10,
   O => W_38_15_i_17_n_0
);
W_38_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x80_out_24,
   I1 => x80_out_31,
   I2 => x80_out_1,
   I3 => W_38_15_i_10_n_0,
   I4 => W_38_15_i_11_n_0,
   O => W_38_15_i_2_n_0
);
W_38_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x80_out_23,
   I1 => x80_out_30,
   I2 => x80_out_0,
   I3 => W_38_15_i_12_n_0,
   I4 => W_38_15_i_13_n_0,
   O => W_38_15_i_3_n_0
);
W_38_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x80_out_22,
   I1 => x80_out_29,
   I2 => x80_out_31,
   I3 => W_38_15_i_14_n_0,
   I4 => W_38_15_i_15_n_0,
   O => W_38_15_i_4_n_0
);
W_38_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x80_out_21,
   I1 => x80_out_28,
   I2 => x80_out_30,
   I3 => W_38_15_i_16_n_0,
   I4 => W_38_15_i_17_n_0,
   O => W_38_15_i_5_n_0
);
W_38_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_38_15_i_2_n_0,
   I1 => W_38_19_i_16_n_0,
   I2 => x80_out_25,
   I3 => x80_out_0,
   I4 => x80_out_2,
   I5 => W_38_19_i_17_n_0,
   O => W_38_15_i_6_n_0
);
W_38_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_38_15_i_3_n_0,
   I1 => W_38_15_i_10_n_0,
   I2 => x80_out_24,
   I3 => x80_out_31,
   I4 => x80_out_1,
   I5 => W_38_15_i_11_n_0,
   O => W_38_15_i_7_n_0
);
W_38_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_38_15_i_4_n_0,
   I1 => W_38_15_i_12_n_0,
   I2 => x80_out_23,
   I3 => x80_out_30,
   I4 => x80_out_0,
   I5 => W_38_15_i_13_n_0,
   O => W_38_15_i_8_n_0
);
W_38_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_38_15_i_5_n_0,
   I1 => W_38_15_i_14_n_0,
   I2 => x80_out_22,
   I3 => x80_out_29,
   I4 => x80_out_31,
   I5 => W_38_15_i_15_n_0,
   O => W_38_15_i_9_n_0
);
W_38_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x111_out_18,
   I1 => x94_out_18,
   I2 => x110_out_4,
   I3 => x110_out_25,
   I4 => x110_out_21,
   O => W_38_19_i_10_n_0
);
W_38_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x94_out_17,
   I1 => x110_out_20,
   I2 => x110_out_24,
   I3 => x110_out_3,
   I4 => x111_out_17,
   O => W_38_19_i_11_n_0
);
W_38_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x111_out_17,
   I1 => x94_out_17,
   I2 => x110_out_3,
   I3 => x110_out_24,
   I4 => x110_out_20,
   O => W_38_19_i_12_n_0
);
W_38_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x94_out_16,
   I1 => x110_out_19,
   I2 => x110_out_23,
   I3 => x110_out_2,
   I4 => x111_out_16,
   O => W_38_19_i_13_n_0
);
W_38_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x111_out_16,
   I1 => x94_out_16,
   I2 => x110_out_2,
   I3 => x110_out_23,
   I4 => x110_out_19,
   O => W_38_19_i_14_n_0
);
W_38_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x94_out_15,
   I1 => x110_out_18,
   I2 => x110_out_22,
   I3 => x110_out_1,
   I4 => x111_out_15,
   O => W_38_19_i_15_n_0
);
W_38_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x111_out_15,
   I1 => x94_out_15,
   I2 => x110_out_1,
   I3 => x110_out_22,
   I4 => x110_out_18,
   O => W_38_19_i_16_n_0
);
W_38_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x94_out_14,
   I1 => x110_out_17,
   I2 => x110_out_21,
   I3 => x110_out_0,
   I4 => x111_out_14,
   O => W_38_19_i_17_n_0
);
W_38_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x80_out_28,
   I1 => x80_out_3,
   I2 => x80_out_5,
   I3 => W_38_19_i_10_n_0,
   I4 => W_38_19_i_11_n_0,
   O => W_38_19_i_2_n_0
);
W_38_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x80_out_27,
   I1 => x80_out_2,
   I2 => x80_out_4,
   I3 => W_38_19_i_12_n_0,
   I4 => W_38_19_i_13_n_0,
   O => W_38_19_i_3_n_0
);
W_38_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x80_out_26,
   I1 => x80_out_1,
   I2 => x80_out_3,
   I3 => W_38_19_i_14_n_0,
   I4 => W_38_19_i_15_n_0,
   O => W_38_19_i_4_n_0
);
W_38_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x80_out_25,
   I1 => x80_out_0,
   I2 => x80_out_2,
   I3 => W_38_19_i_16_n_0,
   I4 => W_38_19_i_17_n_0,
   O => W_38_19_i_5_n_0
);
W_38_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_38_19_i_2_n_0,
   I1 => W_38_23_i_16_n_0,
   I2 => x80_out_29,
   I3 => x80_out_4,
   I4 => x80_out_6,
   I5 => W_38_23_i_17_n_0,
   O => W_38_19_i_6_n_0
);
W_38_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_38_19_i_3_n_0,
   I1 => W_38_19_i_10_n_0,
   I2 => x80_out_28,
   I3 => x80_out_3,
   I4 => x80_out_5,
   I5 => W_38_19_i_11_n_0,
   O => W_38_19_i_7_n_0
);
W_38_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_38_19_i_4_n_0,
   I1 => W_38_19_i_12_n_0,
   I2 => x80_out_27,
   I3 => x80_out_2,
   I4 => x80_out_4,
   I5 => W_38_19_i_13_n_0,
   O => W_38_19_i_8_n_0
);
W_38_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_38_19_i_5_n_0,
   I1 => W_38_19_i_14_n_0,
   I2 => x80_out_26,
   I3 => x80_out_1,
   I4 => x80_out_3,
   I5 => W_38_19_i_15_n_0,
   O => W_38_19_i_9_n_0
);
W_38_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x111_out_22,
   I1 => x94_out_22,
   I2 => x110_out_8,
   I3 => x110_out_29,
   I4 => x110_out_25,
   O => W_38_23_i_10_n_0
);
W_38_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x94_out_21,
   I1 => x110_out_24,
   I2 => x110_out_28,
   I3 => x110_out_7,
   I4 => x111_out_21,
   O => W_38_23_i_11_n_0
);
W_38_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x111_out_21,
   I1 => x94_out_21,
   I2 => x110_out_7,
   I3 => x110_out_28,
   I4 => x110_out_24,
   O => W_38_23_i_12_n_0
);
W_38_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x94_out_20,
   I1 => x110_out_23,
   I2 => x110_out_27,
   I3 => x110_out_6,
   I4 => x111_out_20,
   O => W_38_23_i_13_n_0
);
W_38_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x111_out_20,
   I1 => x94_out_20,
   I2 => x110_out_6,
   I3 => x110_out_27,
   I4 => x110_out_23,
   O => W_38_23_i_14_n_0
);
W_38_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x94_out_19,
   I1 => x110_out_22,
   I2 => x110_out_26,
   I3 => x110_out_5,
   I4 => x111_out_19,
   O => W_38_23_i_15_n_0
);
W_38_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x111_out_19,
   I1 => x94_out_19,
   I2 => x110_out_5,
   I3 => x110_out_26,
   I4 => x110_out_22,
   O => W_38_23_i_16_n_0
);
W_38_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x94_out_18,
   I1 => x110_out_21,
   I2 => x110_out_25,
   I3 => x110_out_4,
   I4 => x111_out_18,
   O => W_38_23_i_17_n_0
);
W_38_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x80_out_7,
   I1 => x80_out_9,
   I2 => W_38_23_i_10_n_0,
   I3 => W_38_23_i_11_n_0,
   O => W_38_23_i_2_n_0
);
W_38_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x80_out_31,
   I1 => x80_out_6,
   I2 => x80_out_8,
   I3 => W_38_23_i_12_n_0,
   I4 => W_38_23_i_13_n_0,
   O => W_38_23_i_3_n_0
);
W_38_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x80_out_30,
   I1 => x80_out_5,
   I2 => x80_out_7,
   I3 => W_38_23_i_14_n_0,
   I4 => W_38_23_i_15_n_0,
   O => W_38_23_i_4_n_0
);
W_38_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x80_out_29,
   I1 => x80_out_4,
   I2 => x80_out_6,
   I3 => W_38_23_i_16_n_0,
   I4 => W_38_23_i_17_n_0,
   O => W_38_23_i_5_n_0
);
W_38_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x80_out_8,
   I1 => x80_out_10,
   I2 => W_38_27_i_16_n_0,
   I3 => W_38_27_i_17_n_0,
   I4 => W_38_23_i_2_n_0,
   O => W_38_23_i_6_n_0
);
W_38_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x80_out_7,
   I1 => x80_out_9,
   I2 => W_38_23_i_10_n_0,
   I3 => W_38_23_i_11_n_0,
   I4 => W_38_23_i_3_n_0,
   O => W_38_23_i_7_n_0
);
W_38_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_38_23_i_4_n_0,
   I1 => W_38_23_i_12_n_0,
   I2 => x80_out_31,
   I3 => x80_out_6,
   I4 => x80_out_8,
   I5 => W_38_23_i_13_n_0,
   O => W_38_23_i_8_n_0
);
W_38_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_38_23_i_5_n_0,
   I1 => W_38_23_i_14_n_0,
   I2 => x80_out_30,
   I3 => x80_out_5,
   I4 => x80_out_7,
   I5 => W_38_23_i_15_n_0,
   O => W_38_23_i_9_n_0
);
W_38_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x111_out_26,
   I1 => x94_out_26,
   I2 => x110_out_12,
   I3 => x110_out_1,
   I4 => x110_out_29,
   O => W_38_27_i_10_n_0
);
W_38_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x94_out_25,
   I1 => x110_out_28,
   I2 => x110_out_0,
   I3 => x110_out_11,
   I4 => x111_out_25,
   O => W_38_27_i_11_n_0
);
W_38_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x111_out_25,
   I1 => x94_out_25,
   I2 => x110_out_11,
   I3 => x110_out_0,
   I4 => x110_out_28,
   O => W_38_27_i_12_n_0
);
W_38_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x94_out_24,
   I1 => x110_out_27,
   I2 => x110_out_31,
   I3 => x110_out_10,
   I4 => x111_out_24,
   O => W_38_27_i_13_n_0
);
W_38_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x111_out_24,
   I1 => x94_out_24,
   I2 => x110_out_10,
   I3 => x110_out_31,
   I4 => x110_out_27,
   O => W_38_27_i_14_n_0
);
W_38_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x94_out_23,
   I1 => x110_out_26,
   I2 => x110_out_30,
   I3 => x110_out_9,
   I4 => x111_out_23,
   O => W_38_27_i_15_n_0
);
W_38_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x111_out_23,
   I1 => x94_out_23,
   I2 => x110_out_9,
   I3 => x110_out_30,
   I4 => x110_out_26,
   O => W_38_27_i_16_n_0
);
W_38_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x94_out_22,
   I1 => x110_out_25,
   I2 => x110_out_29,
   I3 => x110_out_8,
   I4 => x111_out_22,
   O => W_38_27_i_17_n_0
);
W_38_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x80_out_11,
   I1 => x80_out_13,
   I2 => W_38_27_i_10_n_0,
   I3 => W_38_27_i_11_n_0,
   O => W_38_27_i_2_n_0
);
W_38_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x80_out_10,
   I1 => x80_out_12,
   I2 => W_38_27_i_12_n_0,
   I3 => W_38_27_i_13_n_0,
   O => W_38_27_i_3_n_0
);
W_38_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x80_out_9,
   I1 => x80_out_11,
   I2 => W_38_27_i_14_n_0,
   I3 => W_38_27_i_15_n_0,
   O => W_38_27_i_4_n_0
);
W_38_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x80_out_8,
   I1 => x80_out_10,
   I2 => W_38_27_i_16_n_0,
   I3 => W_38_27_i_17_n_0,
   O => W_38_27_i_5_n_0
);
W_38_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x80_out_12,
   I1 => x80_out_14,
   I2 => W_38_31_i_13_n_0,
   I3 => W_38_31_i_14_n_0,
   I4 => W_38_27_i_2_n_0,
   O => W_38_27_i_6_n_0
);
W_38_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x80_out_11,
   I1 => x80_out_13,
   I2 => W_38_27_i_10_n_0,
   I3 => W_38_27_i_11_n_0,
   I4 => W_38_27_i_3_n_0,
   O => W_38_27_i_7_n_0
);
W_38_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x80_out_10,
   I1 => x80_out_12,
   I2 => W_38_27_i_12_n_0,
   I3 => W_38_27_i_13_n_0,
   I4 => W_38_27_i_4_n_0,
   O => W_38_27_i_8_n_0
);
W_38_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x80_out_9,
   I1 => x80_out_11,
   I2 => W_38_27_i_14_n_0,
   I3 => W_38_27_i_15_n_0,
   I4 => W_38_27_i_5_n_0,
   O => W_38_27_i_9_n_0
);
W_38_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x94_out_28,
   I1 => x110_out_31,
   I2 => x110_out_3,
   I3 => x110_out_14,
   I4 => x111_out_28,
   O => W_38_31_i_10_n_0
);
W_38_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x111_out_28,
   I1 => x94_out_28,
   I2 => x110_out_14,
   I3 => x110_out_3,
   I4 => x110_out_31,
   O => W_38_31_i_11_n_0
);
W_38_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x94_out_27,
   I1 => x110_out_30,
   I2 => x110_out_2,
   I3 => x110_out_13,
   I4 => x111_out_27,
   O => W_38_31_i_12_n_0
);
W_38_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x111_out_27,
   I1 => x94_out_27,
   I2 => x110_out_13,
   I3 => x110_out_2,
   I4 => x110_out_30,
   O => W_38_31_i_13_n_0
);
W_38_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x94_out_26,
   I1 => x110_out_29,
   I2 => x110_out_1,
   I3 => x110_out_12,
   I4 => x111_out_26,
   O => W_38_31_i_14_n_0
);
W_38_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x94_out_29,
   I1 => x110_out_4,
   I2 => x110_out_15,
   I3 => x111_out_29,
   O => W_38_31_i_15_n_0
);
W_38_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x80_out_17,
   I1 => x80_out_15,
   O => SIGMA_LCASE_1211_out_0_30
);
W_38_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => x110_out_6,
   I1 => x110_out_17,
   I2 => x94_out_31,
   I3 => x111_out_31,
   I4 => x80_out_16,
   I5 => x80_out_18,
   O => W_38_31_i_17_n_0
);
W_38_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x110_out_16,
   I1 => x110_out_5,
   O => SIGMA_LCASE_0207_out_30
);
W_38_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x111_out_30,
   I1 => x94_out_30,
   I2 => x110_out_16,
   I3 => x110_out_5,
   O => W_38_31_i_19_n_0
);
W_38_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x80_out_14,
   I1 => x80_out_16,
   I2 => W_38_31_i_9_n_0,
   I3 => W_38_31_i_10_n_0,
   O => W_38_31_i_2_n_0
);
W_38_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x80_out_13,
   I1 => x80_out_15,
   I2 => W_38_31_i_11_n_0,
   I3 => W_38_31_i_12_n_0,
   O => W_38_31_i_3_n_0
);
W_38_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x80_out_12,
   I1 => x80_out_14,
   I2 => W_38_31_i_13_n_0,
   I3 => W_38_31_i_14_n_0,
   O => W_38_31_i_4_n_0
);
W_38_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_38_31_i_15_n_0,
   I1 => SIGMA_LCASE_1211_out_0_30,
   I2 => W_38_31_i_17_n_0,
   I3 => x94_out_30,
   I4 => SIGMA_LCASE_0207_out_30,
   I5 => x111_out_30,
   O => W_38_31_i_5_n_0
);
W_38_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_38_31_i_2_n_0,
   I1 => W_38_31_i_19_n_0,
   I2 => x80_out_15,
   I3 => x80_out_17,
   I4 => W_38_31_i_15_n_0,
   O => W_38_31_i_6_n_0
);
W_38_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x80_out_14,
   I1 => x80_out_16,
   I2 => W_38_31_i_9_n_0,
   I3 => W_38_31_i_10_n_0,
   I4 => W_38_31_i_3_n_0,
   O => W_38_31_i_7_n_0
);
W_38_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x80_out_13,
   I1 => x80_out_15,
   I2 => W_38_31_i_11_n_0,
   I3 => W_38_31_i_12_n_0,
   I4 => W_38_31_i_4_n_0,
   O => W_38_31_i_8_n_0
);
W_38_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x111_out_29,
   I1 => x94_out_29,
   I2 => x110_out_15,
   I3 => x110_out_4,
   O => W_38_31_i_9_n_0
);
W_38_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x111_out_2,
   I1 => x94_out_2,
   I2 => x110_out_20,
   I3 => x110_out_9,
   I4 => x110_out_5,
   O => W_38_3_i_10_n_0
);
W_38_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x94_out_1,
   I1 => x110_out_4,
   I2 => x110_out_8,
   I3 => x110_out_19,
   I4 => x111_out_1,
   O => W_38_3_i_11_n_0
);
W_38_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x110_out_19,
   I1 => x110_out_8,
   I2 => x110_out_4,
   O => SIGMA_LCASE_0207_out_1
);
W_38_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x80_out_21,
   I1 => x80_out_19,
   I2 => x80_out_12,
   O => SIGMA_LCASE_1211_out_0_2
);
W_38_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x80_out_20,
   I1 => x80_out_18,
   I2 => x80_out_11,
   O => SIGMA_LCASE_1211_out_1
);
W_38_3_i_15 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x111_out_1,
   I1 => x94_out_1,
   I2 => x110_out_19,
   I3 => x110_out_8,
   I4 => x110_out_4,
   O => W_38_3_i_15_n_0
);
W_38_3_i_16 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x110_out_18,
   I1 => x110_out_7,
   I2 => x110_out_3,
   O => SIGMA_LCASE_0207_out_0
);
W_38_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x80_out_12,
   I1 => x80_out_19,
   I2 => x80_out_21,
   I3 => W_38_3_i_10_n_0,
   I4 => W_38_3_i_11_n_0,
   O => W_38_3_i_2_n_0
);
W_38_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_38_3_i_11_n_0,
   I1 => x80_out_21,
   I2 => x80_out_19,
   I3 => x80_out_12,
   I4 => W_38_3_i_10_n_0,
   O => W_38_3_i_3_n_0
);
W_38_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_0207_out_1,
   I1 => x94_out_1,
   I2 => x111_out_1,
   I3 => x80_out_11,
   I4 => x80_out_18,
   I5 => x80_out_20,
   O => W_38_3_i_4_n_0
);
W_38_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x111_out_0,
   I1 => x94_out_0,
   I2 => x110_out_18,
   I3 => x110_out_7,
   I4 => x110_out_3,
   O => W_38_3_i_5_n_0
);
W_38_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_38_3_i_2_n_0,
   I1 => W_38_7_i_16_n_0,
   I2 => x80_out_13,
   I3 => x80_out_20,
   I4 => x80_out_22,
   I5 => W_38_7_i_17_n_0,
   O => W_38_3_i_6_n_0
);
W_38_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_38_3_i_10_n_0,
   I1 => SIGMA_LCASE_1211_out_0_2,
   I2 => x111_out_1,
   I3 => x94_out_1,
   I4 => SIGMA_LCASE_0207_out_1,
   I5 => SIGMA_LCASE_1211_out_1,
   O => W_38_3_i_7_n_0
);
W_38_3_i_8 : LUT5
  generic map(
   INIT => X"99969666"
  )
 port map (
   I0 => SIGMA_LCASE_1211_out_1,
   I1 => W_38_3_i_15_n_0,
   I2 => x111_out_0,
   I3 => SIGMA_LCASE_0207_out_0,
   I4 => x94_out_0,
   O => W_38_3_i_8_n_0
);
W_38_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_38_3_i_5_n_0,
   I1 => x80_out_10,
   I2 => x80_out_17,
   I3 => x80_out_19,
   O => W_38_3_i_9_n_0
);
W_38_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x111_out_6,
   I1 => x94_out_6,
   I2 => x110_out_24,
   I3 => x110_out_13,
   I4 => x110_out_9,
   O => W_38_7_i_10_n_0
);
W_38_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x94_out_5,
   I1 => x110_out_8,
   I2 => x110_out_12,
   I3 => x110_out_23,
   I4 => x111_out_5,
   O => W_38_7_i_11_n_0
);
W_38_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x111_out_5,
   I1 => x94_out_5,
   I2 => x110_out_23,
   I3 => x110_out_12,
   I4 => x110_out_8,
   O => W_38_7_i_12_n_0
);
W_38_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x94_out_4,
   I1 => x110_out_7,
   I2 => x110_out_11,
   I3 => x110_out_22,
   I4 => x111_out_4,
   O => W_38_7_i_13_n_0
);
W_38_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x111_out_4,
   I1 => x94_out_4,
   I2 => x110_out_22,
   I3 => x110_out_11,
   I4 => x110_out_7,
   O => W_38_7_i_14_n_0
);
W_38_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x94_out_3,
   I1 => x110_out_6,
   I2 => x110_out_10,
   I3 => x110_out_21,
   I4 => x111_out_3,
   O => W_38_7_i_15_n_0
);
W_38_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x111_out_3,
   I1 => x94_out_3,
   I2 => x110_out_21,
   I3 => x110_out_10,
   I4 => x110_out_6,
   O => W_38_7_i_16_n_0
);
W_38_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x94_out_2,
   I1 => x110_out_5,
   I2 => x110_out_9,
   I3 => x110_out_20,
   I4 => x111_out_2,
   O => W_38_7_i_17_n_0
);
W_38_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x80_out_16,
   I1 => x80_out_23,
   I2 => x80_out_25,
   I3 => W_38_7_i_10_n_0,
   I4 => W_38_7_i_11_n_0,
   O => W_38_7_i_2_n_0
);
W_38_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x80_out_15,
   I1 => x80_out_22,
   I2 => x80_out_24,
   I3 => W_38_7_i_12_n_0,
   I4 => W_38_7_i_13_n_0,
   O => W_38_7_i_3_n_0
);
W_38_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x80_out_14,
   I1 => x80_out_21,
   I2 => x80_out_23,
   I3 => W_38_7_i_14_n_0,
   I4 => W_38_7_i_15_n_0,
   O => W_38_7_i_4_n_0
);
W_38_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x80_out_13,
   I1 => x80_out_20,
   I2 => x80_out_22,
   I3 => W_38_7_i_16_n_0,
   I4 => W_38_7_i_17_n_0,
   O => W_38_7_i_5_n_0
);
W_38_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_38_7_i_2_n_0,
   I1 => W_38_11_i_16_n_0,
   I2 => x80_out_17,
   I3 => x80_out_24,
   I4 => x80_out_26,
   I5 => W_38_11_i_17_n_0,
   O => W_38_7_i_6_n_0
);
W_38_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_38_7_i_3_n_0,
   I1 => W_38_7_i_10_n_0,
   I2 => x80_out_16,
   I3 => x80_out_23,
   I4 => x80_out_25,
   I5 => W_38_7_i_11_n_0,
   O => W_38_7_i_7_n_0
);
W_38_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_38_7_i_4_n_0,
   I1 => W_38_7_i_12_n_0,
   I2 => x80_out_15,
   I3 => x80_out_22,
   I4 => x80_out_24,
   I5 => W_38_7_i_13_n_0,
   O => W_38_7_i_8_n_0
);
W_38_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_38_7_i_5_n_0,
   I1 => W_38_7_i_14_n_0,
   I2 => x80_out_14,
   I3 => x80_out_21,
   I4 => x80_out_23,
   I5 => W_38_7_i_15_n_0,
   O => W_38_7_i_9_n_0
);
W_39_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x110_out_10,
   I1 => x92_out_10,
   I2 => x108_out_28,
   I3 => x108_out_17,
   I4 => x108_out_13,
   O => W_39_11_i_10_n_0
);
W_39_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x92_out_9,
   I1 => x108_out_12,
   I2 => x108_out_16,
   I3 => x108_out_27,
   I4 => x110_out_9,
   O => W_39_11_i_11_n_0
);
W_39_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x110_out_9,
   I1 => x92_out_9,
   I2 => x108_out_27,
   I3 => x108_out_16,
   I4 => x108_out_12,
   O => W_39_11_i_12_n_0
);
W_39_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x92_out_8,
   I1 => x108_out_11,
   I2 => x108_out_15,
   I3 => x108_out_26,
   I4 => x110_out_8,
   O => W_39_11_i_13_n_0
);
W_39_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x110_out_8,
   I1 => x92_out_8,
   I2 => x108_out_26,
   I3 => x108_out_15,
   I4 => x108_out_11,
   O => W_39_11_i_14_n_0
);
W_39_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x92_out_7,
   I1 => x108_out_10,
   I2 => x108_out_14,
   I3 => x108_out_25,
   I4 => x110_out_7,
   O => W_39_11_i_15_n_0
);
W_39_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x110_out_7,
   I1 => x92_out_7,
   I2 => x108_out_25,
   I3 => x108_out_14,
   I4 => x108_out_10,
   O => W_39_11_i_16_n_0
);
W_39_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x92_out_6,
   I1 => x108_out_9,
   I2 => x108_out_13,
   I3 => x108_out_24,
   I4 => x110_out_6,
   O => W_39_11_i_17_n_0
);
W_39_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x77_out_20,
   I1 => x77_out_27,
   I2 => x77_out_29,
   I3 => W_39_11_i_10_n_0,
   I4 => W_39_11_i_11_n_0,
   O => W_39_11_i_2_n_0
);
W_39_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x77_out_19,
   I1 => x77_out_26,
   I2 => x77_out_28,
   I3 => W_39_11_i_12_n_0,
   I4 => W_39_11_i_13_n_0,
   O => W_39_11_i_3_n_0
);
W_39_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x77_out_18,
   I1 => x77_out_25,
   I2 => x77_out_27,
   I3 => W_39_11_i_14_n_0,
   I4 => W_39_11_i_15_n_0,
   O => W_39_11_i_4_n_0
);
W_39_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x77_out_17,
   I1 => x77_out_24,
   I2 => x77_out_26,
   I3 => W_39_11_i_16_n_0,
   I4 => W_39_11_i_17_n_0,
   O => W_39_11_i_5_n_0
);
W_39_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_39_11_i_2_n_0,
   I1 => W_39_15_i_16_n_0,
   I2 => x77_out_21,
   I3 => x77_out_28,
   I4 => x77_out_30,
   I5 => W_39_15_i_17_n_0,
   O => W_39_11_i_6_n_0
);
W_39_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_39_11_i_3_n_0,
   I1 => W_39_11_i_10_n_0,
   I2 => x77_out_20,
   I3 => x77_out_27,
   I4 => x77_out_29,
   I5 => W_39_11_i_11_n_0,
   O => W_39_11_i_7_n_0
);
W_39_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_39_11_i_4_n_0,
   I1 => W_39_11_i_12_n_0,
   I2 => x77_out_19,
   I3 => x77_out_26,
   I4 => x77_out_28,
   I5 => W_39_11_i_13_n_0,
   O => W_39_11_i_8_n_0
);
W_39_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_39_11_i_5_n_0,
   I1 => W_39_11_i_14_n_0,
   I2 => x77_out_18,
   I3 => x77_out_25,
   I4 => x77_out_27,
   I5 => W_39_11_i_15_n_0,
   O => W_39_11_i_9_n_0
);
W_39_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x110_out_14,
   I1 => x92_out_14,
   I2 => x108_out_0,
   I3 => x108_out_21,
   I4 => x108_out_17,
   O => W_39_15_i_10_n_0
);
W_39_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x92_out_13,
   I1 => x108_out_16,
   I2 => x108_out_20,
   I3 => x108_out_31,
   I4 => x110_out_13,
   O => W_39_15_i_11_n_0
);
W_39_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x110_out_13,
   I1 => x92_out_13,
   I2 => x108_out_31,
   I3 => x108_out_20,
   I4 => x108_out_16,
   O => W_39_15_i_12_n_0
);
W_39_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x92_out_12,
   I1 => x108_out_15,
   I2 => x108_out_19,
   I3 => x108_out_30,
   I4 => x110_out_12,
   O => W_39_15_i_13_n_0
);
W_39_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x110_out_12,
   I1 => x92_out_12,
   I2 => x108_out_30,
   I3 => x108_out_19,
   I4 => x108_out_15,
   O => W_39_15_i_14_n_0
);
W_39_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x92_out_11,
   I1 => x108_out_14,
   I2 => x108_out_18,
   I3 => x108_out_29,
   I4 => x110_out_11,
   O => W_39_15_i_15_n_0
);
W_39_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x110_out_11,
   I1 => x92_out_11,
   I2 => x108_out_29,
   I3 => x108_out_18,
   I4 => x108_out_14,
   O => W_39_15_i_16_n_0
);
W_39_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x92_out_10,
   I1 => x108_out_13,
   I2 => x108_out_17,
   I3 => x108_out_28,
   I4 => x110_out_10,
   O => W_39_15_i_17_n_0
);
W_39_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x77_out_24,
   I1 => x77_out_31,
   I2 => x77_out_1,
   I3 => W_39_15_i_10_n_0,
   I4 => W_39_15_i_11_n_0,
   O => W_39_15_i_2_n_0
);
W_39_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x77_out_23,
   I1 => x77_out_30,
   I2 => x77_out_0,
   I3 => W_39_15_i_12_n_0,
   I4 => W_39_15_i_13_n_0,
   O => W_39_15_i_3_n_0
);
W_39_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x77_out_22,
   I1 => x77_out_29,
   I2 => x77_out_31,
   I3 => W_39_15_i_14_n_0,
   I4 => W_39_15_i_15_n_0,
   O => W_39_15_i_4_n_0
);
W_39_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x77_out_21,
   I1 => x77_out_28,
   I2 => x77_out_30,
   I3 => W_39_15_i_16_n_0,
   I4 => W_39_15_i_17_n_0,
   O => W_39_15_i_5_n_0
);
W_39_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_39_15_i_2_n_0,
   I1 => W_39_19_i_16_n_0,
   I2 => x77_out_25,
   I3 => x77_out_0,
   I4 => x77_out_2,
   I5 => W_39_19_i_17_n_0,
   O => W_39_15_i_6_n_0
);
W_39_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_39_15_i_3_n_0,
   I1 => W_39_15_i_10_n_0,
   I2 => x77_out_24,
   I3 => x77_out_31,
   I4 => x77_out_1,
   I5 => W_39_15_i_11_n_0,
   O => W_39_15_i_7_n_0
);
W_39_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_39_15_i_4_n_0,
   I1 => W_39_15_i_12_n_0,
   I2 => x77_out_23,
   I3 => x77_out_30,
   I4 => x77_out_0,
   I5 => W_39_15_i_13_n_0,
   O => W_39_15_i_8_n_0
);
W_39_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_39_15_i_5_n_0,
   I1 => W_39_15_i_14_n_0,
   I2 => x77_out_22,
   I3 => x77_out_29,
   I4 => x77_out_31,
   I5 => W_39_15_i_15_n_0,
   O => W_39_15_i_9_n_0
);
W_39_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x110_out_18,
   I1 => x92_out_18,
   I2 => x108_out_4,
   I3 => x108_out_25,
   I4 => x108_out_21,
   O => W_39_19_i_10_n_0
);
W_39_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x92_out_17,
   I1 => x108_out_20,
   I2 => x108_out_24,
   I3 => x108_out_3,
   I4 => x110_out_17,
   O => W_39_19_i_11_n_0
);
W_39_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x110_out_17,
   I1 => x92_out_17,
   I2 => x108_out_3,
   I3 => x108_out_24,
   I4 => x108_out_20,
   O => W_39_19_i_12_n_0
);
W_39_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x92_out_16,
   I1 => x108_out_19,
   I2 => x108_out_23,
   I3 => x108_out_2,
   I4 => x110_out_16,
   O => W_39_19_i_13_n_0
);
W_39_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x110_out_16,
   I1 => x92_out_16,
   I2 => x108_out_2,
   I3 => x108_out_23,
   I4 => x108_out_19,
   O => W_39_19_i_14_n_0
);
W_39_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x92_out_15,
   I1 => x108_out_18,
   I2 => x108_out_22,
   I3 => x108_out_1,
   I4 => x110_out_15,
   O => W_39_19_i_15_n_0
);
W_39_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x110_out_15,
   I1 => x92_out_15,
   I2 => x108_out_1,
   I3 => x108_out_22,
   I4 => x108_out_18,
   O => W_39_19_i_16_n_0
);
W_39_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x92_out_14,
   I1 => x108_out_17,
   I2 => x108_out_21,
   I3 => x108_out_0,
   I4 => x110_out_14,
   O => W_39_19_i_17_n_0
);
W_39_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x77_out_28,
   I1 => x77_out_3,
   I2 => x77_out_5,
   I3 => W_39_19_i_10_n_0,
   I4 => W_39_19_i_11_n_0,
   O => W_39_19_i_2_n_0
);
W_39_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x77_out_27,
   I1 => x77_out_2,
   I2 => x77_out_4,
   I3 => W_39_19_i_12_n_0,
   I4 => W_39_19_i_13_n_0,
   O => W_39_19_i_3_n_0
);
W_39_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x77_out_26,
   I1 => x77_out_1,
   I2 => x77_out_3,
   I3 => W_39_19_i_14_n_0,
   I4 => W_39_19_i_15_n_0,
   O => W_39_19_i_4_n_0
);
W_39_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x77_out_25,
   I1 => x77_out_0,
   I2 => x77_out_2,
   I3 => W_39_19_i_16_n_0,
   I4 => W_39_19_i_17_n_0,
   O => W_39_19_i_5_n_0
);
W_39_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_39_19_i_2_n_0,
   I1 => W_39_23_i_16_n_0,
   I2 => x77_out_29,
   I3 => x77_out_4,
   I4 => x77_out_6,
   I5 => W_39_23_i_17_n_0,
   O => W_39_19_i_6_n_0
);
W_39_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_39_19_i_3_n_0,
   I1 => W_39_19_i_10_n_0,
   I2 => x77_out_28,
   I3 => x77_out_3,
   I4 => x77_out_5,
   I5 => W_39_19_i_11_n_0,
   O => W_39_19_i_7_n_0
);
W_39_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_39_19_i_4_n_0,
   I1 => W_39_19_i_12_n_0,
   I2 => x77_out_27,
   I3 => x77_out_2,
   I4 => x77_out_4,
   I5 => W_39_19_i_13_n_0,
   O => W_39_19_i_8_n_0
);
W_39_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_39_19_i_5_n_0,
   I1 => W_39_19_i_14_n_0,
   I2 => x77_out_26,
   I3 => x77_out_1,
   I4 => x77_out_3,
   I5 => W_39_19_i_15_n_0,
   O => W_39_19_i_9_n_0
);
W_39_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x110_out_22,
   I1 => x92_out_22,
   I2 => x108_out_8,
   I3 => x108_out_29,
   I4 => x108_out_25,
   O => W_39_23_i_10_n_0
);
W_39_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x92_out_21,
   I1 => x108_out_24,
   I2 => x108_out_28,
   I3 => x108_out_7,
   I4 => x110_out_21,
   O => W_39_23_i_11_n_0
);
W_39_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x110_out_21,
   I1 => x92_out_21,
   I2 => x108_out_7,
   I3 => x108_out_28,
   I4 => x108_out_24,
   O => W_39_23_i_12_n_0
);
W_39_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x92_out_20,
   I1 => x108_out_23,
   I2 => x108_out_27,
   I3 => x108_out_6,
   I4 => x110_out_20,
   O => W_39_23_i_13_n_0
);
W_39_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x110_out_20,
   I1 => x92_out_20,
   I2 => x108_out_6,
   I3 => x108_out_27,
   I4 => x108_out_23,
   O => W_39_23_i_14_n_0
);
W_39_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x92_out_19,
   I1 => x108_out_22,
   I2 => x108_out_26,
   I3 => x108_out_5,
   I4 => x110_out_19,
   O => W_39_23_i_15_n_0
);
W_39_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x110_out_19,
   I1 => x92_out_19,
   I2 => x108_out_5,
   I3 => x108_out_26,
   I4 => x108_out_22,
   O => W_39_23_i_16_n_0
);
W_39_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x92_out_18,
   I1 => x108_out_21,
   I2 => x108_out_25,
   I3 => x108_out_4,
   I4 => x110_out_18,
   O => W_39_23_i_17_n_0
);
W_39_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x77_out_7,
   I1 => x77_out_9,
   I2 => W_39_23_i_10_n_0,
   I3 => W_39_23_i_11_n_0,
   O => W_39_23_i_2_n_0
);
W_39_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x77_out_31,
   I1 => x77_out_6,
   I2 => x77_out_8,
   I3 => W_39_23_i_12_n_0,
   I4 => W_39_23_i_13_n_0,
   O => W_39_23_i_3_n_0
);
W_39_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x77_out_30,
   I1 => x77_out_5,
   I2 => x77_out_7,
   I3 => W_39_23_i_14_n_0,
   I4 => W_39_23_i_15_n_0,
   O => W_39_23_i_4_n_0
);
W_39_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x77_out_29,
   I1 => x77_out_4,
   I2 => x77_out_6,
   I3 => W_39_23_i_16_n_0,
   I4 => W_39_23_i_17_n_0,
   O => W_39_23_i_5_n_0
);
W_39_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x77_out_8,
   I1 => x77_out_10,
   I2 => W_39_27_i_16_n_0,
   I3 => W_39_27_i_17_n_0,
   I4 => W_39_23_i_2_n_0,
   O => W_39_23_i_6_n_0
);
W_39_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x77_out_7,
   I1 => x77_out_9,
   I2 => W_39_23_i_10_n_0,
   I3 => W_39_23_i_11_n_0,
   I4 => W_39_23_i_3_n_0,
   O => W_39_23_i_7_n_0
);
W_39_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_39_23_i_4_n_0,
   I1 => W_39_23_i_12_n_0,
   I2 => x77_out_31,
   I3 => x77_out_6,
   I4 => x77_out_8,
   I5 => W_39_23_i_13_n_0,
   O => W_39_23_i_8_n_0
);
W_39_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_39_23_i_5_n_0,
   I1 => W_39_23_i_14_n_0,
   I2 => x77_out_30,
   I3 => x77_out_5,
   I4 => x77_out_7,
   I5 => W_39_23_i_15_n_0,
   O => W_39_23_i_9_n_0
);
W_39_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x110_out_26,
   I1 => x92_out_26,
   I2 => x108_out_12,
   I3 => x108_out_1,
   I4 => x108_out_29,
   O => W_39_27_i_10_n_0
);
W_39_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x92_out_25,
   I1 => x108_out_28,
   I2 => x108_out_0,
   I3 => x108_out_11,
   I4 => x110_out_25,
   O => W_39_27_i_11_n_0
);
W_39_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x110_out_25,
   I1 => x92_out_25,
   I2 => x108_out_11,
   I3 => x108_out_0,
   I4 => x108_out_28,
   O => W_39_27_i_12_n_0
);
W_39_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x92_out_24,
   I1 => x108_out_27,
   I2 => x108_out_31,
   I3 => x108_out_10,
   I4 => x110_out_24,
   O => W_39_27_i_13_n_0
);
W_39_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x110_out_24,
   I1 => x92_out_24,
   I2 => x108_out_10,
   I3 => x108_out_31,
   I4 => x108_out_27,
   O => W_39_27_i_14_n_0
);
W_39_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x92_out_23,
   I1 => x108_out_26,
   I2 => x108_out_30,
   I3 => x108_out_9,
   I4 => x110_out_23,
   O => W_39_27_i_15_n_0
);
W_39_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x110_out_23,
   I1 => x92_out_23,
   I2 => x108_out_9,
   I3 => x108_out_30,
   I4 => x108_out_26,
   O => W_39_27_i_16_n_0
);
W_39_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x92_out_22,
   I1 => x108_out_25,
   I2 => x108_out_29,
   I3 => x108_out_8,
   I4 => x110_out_22,
   O => W_39_27_i_17_n_0
);
W_39_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x77_out_11,
   I1 => x77_out_13,
   I2 => W_39_27_i_10_n_0,
   I3 => W_39_27_i_11_n_0,
   O => W_39_27_i_2_n_0
);
W_39_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x77_out_10,
   I1 => x77_out_12,
   I2 => W_39_27_i_12_n_0,
   I3 => W_39_27_i_13_n_0,
   O => W_39_27_i_3_n_0
);
W_39_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x77_out_9,
   I1 => x77_out_11,
   I2 => W_39_27_i_14_n_0,
   I3 => W_39_27_i_15_n_0,
   O => W_39_27_i_4_n_0
);
W_39_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x77_out_8,
   I1 => x77_out_10,
   I2 => W_39_27_i_16_n_0,
   I3 => W_39_27_i_17_n_0,
   O => W_39_27_i_5_n_0
);
W_39_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x77_out_12,
   I1 => x77_out_14,
   I2 => W_39_31_i_13_n_0,
   I3 => W_39_31_i_14_n_0,
   I4 => W_39_27_i_2_n_0,
   O => W_39_27_i_6_n_0
);
W_39_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x77_out_11,
   I1 => x77_out_13,
   I2 => W_39_27_i_10_n_0,
   I3 => W_39_27_i_11_n_0,
   I4 => W_39_27_i_3_n_0,
   O => W_39_27_i_7_n_0
);
W_39_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x77_out_10,
   I1 => x77_out_12,
   I2 => W_39_27_i_12_n_0,
   I3 => W_39_27_i_13_n_0,
   I4 => W_39_27_i_4_n_0,
   O => W_39_27_i_8_n_0
);
W_39_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x77_out_9,
   I1 => x77_out_11,
   I2 => W_39_27_i_14_n_0,
   I3 => W_39_27_i_15_n_0,
   I4 => W_39_27_i_5_n_0,
   O => W_39_27_i_9_n_0
);
W_39_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x92_out_28,
   I1 => x108_out_31,
   I2 => x108_out_3,
   I3 => x108_out_14,
   I4 => x110_out_28,
   O => W_39_31_i_10_n_0
);
W_39_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x110_out_28,
   I1 => x92_out_28,
   I2 => x108_out_14,
   I3 => x108_out_3,
   I4 => x108_out_31,
   O => W_39_31_i_11_n_0
);
W_39_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x92_out_27,
   I1 => x108_out_30,
   I2 => x108_out_2,
   I3 => x108_out_13,
   I4 => x110_out_27,
   O => W_39_31_i_12_n_0
);
W_39_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x110_out_27,
   I1 => x92_out_27,
   I2 => x108_out_13,
   I3 => x108_out_2,
   I4 => x108_out_30,
   O => W_39_31_i_13_n_0
);
W_39_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x92_out_26,
   I1 => x108_out_29,
   I2 => x108_out_1,
   I3 => x108_out_12,
   I4 => x110_out_26,
   O => W_39_31_i_14_n_0
);
W_39_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x92_out_29,
   I1 => x108_out_4,
   I2 => x108_out_15,
   I3 => x110_out_29,
   O => W_39_31_i_15_n_0
);
W_39_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x77_out_17,
   I1 => x77_out_15,
   O => SIGMA_LCASE_1203_out_0_30
);
W_39_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => x108_out_6,
   I1 => x108_out_17,
   I2 => x92_out_31,
   I3 => x110_out_31,
   I4 => x77_out_16,
   I5 => x77_out_18,
   O => W_39_31_i_17_n_0
);
W_39_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x108_out_16,
   I1 => x108_out_5,
   O => SIGMA_LCASE_0199_out_30
);
W_39_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x110_out_30,
   I1 => x92_out_30,
   I2 => x108_out_16,
   I3 => x108_out_5,
   O => W_39_31_i_19_n_0
);
W_39_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x77_out_14,
   I1 => x77_out_16,
   I2 => W_39_31_i_9_n_0,
   I3 => W_39_31_i_10_n_0,
   O => W_39_31_i_2_n_0
);
W_39_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x77_out_13,
   I1 => x77_out_15,
   I2 => W_39_31_i_11_n_0,
   I3 => W_39_31_i_12_n_0,
   O => W_39_31_i_3_n_0
);
W_39_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x77_out_12,
   I1 => x77_out_14,
   I2 => W_39_31_i_13_n_0,
   I3 => W_39_31_i_14_n_0,
   O => W_39_31_i_4_n_0
);
W_39_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_39_31_i_15_n_0,
   I1 => SIGMA_LCASE_1203_out_0_30,
   I2 => W_39_31_i_17_n_0,
   I3 => x92_out_30,
   I4 => SIGMA_LCASE_0199_out_30,
   I5 => x110_out_30,
   O => W_39_31_i_5_n_0
);
W_39_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_39_31_i_2_n_0,
   I1 => W_39_31_i_19_n_0,
   I2 => x77_out_15,
   I3 => x77_out_17,
   I4 => W_39_31_i_15_n_0,
   O => W_39_31_i_6_n_0
);
W_39_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x77_out_14,
   I1 => x77_out_16,
   I2 => W_39_31_i_9_n_0,
   I3 => W_39_31_i_10_n_0,
   I4 => W_39_31_i_3_n_0,
   O => W_39_31_i_7_n_0
);
W_39_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x77_out_13,
   I1 => x77_out_15,
   I2 => W_39_31_i_11_n_0,
   I3 => W_39_31_i_12_n_0,
   I4 => W_39_31_i_4_n_0,
   O => W_39_31_i_8_n_0
);
W_39_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x110_out_29,
   I1 => x92_out_29,
   I2 => x108_out_15,
   I3 => x108_out_4,
   O => W_39_31_i_9_n_0
);
W_39_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x110_out_2,
   I1 => x92_out_2,
   I2 => x108_out_20,
   I3 => x108_out_9,
   I4 => x108_out_5,
   O => W_39_3_i_10_n_0
);
W_39_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x92_out_1,
   I1 => x108_out_4,
   I2 => x108_out_8,
   I3 => x108_out_19,
   I4 => x110_out_1,
   O => W_39_3_i_11_n_0
);
W_39_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x108_out_19,
   I1 => x108_out_8,
   I2 => x108_out_4,
   O => SIGMA_LCASE_0199_out_1
);
W_39_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x77_out_21,
   I1 => x77_out_19,
   I2 => x77_out_12,
   O => SIGMA_LCASE_1203_out_0_2
);
W_39_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x77_out_20,
   I1 => x77_out_18,
   I2 => x77_out_11,
   O => SIGMA_LCASE_1203_out_1
);
W_39_3_i_15 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x110_out_1,
   I1 => x92_out_1,
   I2 => x108_out_19,
   I3 => x108_out_8,
   I4 => x108_out_4,
   O => W_39_3_i_15_n_0
);
W_39_3_i_16 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x108_out_18,
   I1 => x108_out_7,
   I2 => x108_out_3,
   O => SIGMA_LCASE_0199_out_0
);
W_39_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x77_out_12,
   I1 => x77_out_19,
   I2 => x77_out_21,
   I3 => W_39_3_i_10_n_0,
   I4 => W_39_3_i_11_n_0,
   O => W_39_3_i_2_n_0
);
W_39_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_39_3_i_11_n_0,
   I1 => x77_out_21,
   I2 => x77_out_19,
   I3 => x77_out_12,
   I4 => W_39_3_i_10_n_0,
   O => W_39_3_i_3_n_0
);
W_39_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_0199_out_1,
   I1 => x92_out_1,
   I2 => x110_out_1,
   I3 => x77_out_11,
   I4 => x77_out_18,
   I5 => x77_out_20,
   O => W_39_3_i_4_n_0
);
W_39_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x110_out_0,
   I1 => x92_out_0,
   I2 => x108_out_18,
   I3 => x108_out_7,
   I4 => x108_out_3,
   O => W_39_3_i_5_n_0
);
W_39_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_39_3_i_2_n_0,
   I1 => W_39_7_i_16_n_0,
   I2 => x77_out_13,
   I3 => x77_out_20,
   I4 => x77_out_22,
   I5 => W_39_7_i_17_n_0,
   O => W_39_3_i_6_n_0
);
W_39_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_39_3_i_10_n_0,
   I1 => SIGMA_LCASE_1203_out_0_2,
   I2 => x110_out_1,
   I3 => x92_out_1,
   I4 => SIGMA_LCASE_0199_out_1,
   I5 => SIGMA_LCASE_1203_out_1,
   O => W_39_3_i_7_n_0
);
W_39_3_i_8 : LUT5
  generic map(
   INIT => X"99969666"
  )
 port map (
   I0 => SIGMA_LCASE_1203_out_1,
   I1 => W_39_3_i_15_n_0,
   I2 => x110_out_0,
   I3 => SIGMA_LCASE_0199_out_0,
   I4 => x92_out_0,
   O => W_39_3_i_8_n_0
);
W_39_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_39_3_i_5_n_0,
   I1 => x77_out_10,
   I2 => x77_out_17,
   I3 => x77_out_19,
   O => W_39_3_i_9_n_0
);
W_39_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x110_out_6,
   I1 => x92_out_6,
   I2 => x108_out_24,
   I3 => x108_out_13,
   I4 => x108_out_9,
   O => W_39_7_i_10_n_0
);
W_39_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x92_out_5,
   I1 => x108_out_8,
   I2 => x108_out_12,
   I3 => x108_out_23,
   I4 => x110_out_5,
   O => W_39_7_i_11_n_0
);
W_39_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x110_out_5,
   I1 => x92_out_5,
   I2 => x108_out_23,
   I3 => x108_out_12,
   I4 => x108_out_8,
   O => W_39_7_i_12_n_0
);
W_39_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x92_out_4,
   I1 => x108_out_7,
   I2 => x108_out_11,
   I3 => x108_out_22,
   I4 => x110_out_4,
   O => W_39_7_i_13_n_0
);
W_39_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x110_out_4,
   I1 => x92_out_4,
   I2 => x108_out_22,
   I3 => x108_out_11,
   I4 => x108_out_7,
   O => W_39_7_i_14_n_0
);
W_39_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x92_out_3,
   I1 => x108_out_6,
   I2 => x108_out_10,
   I3 => x108_out_21,
   I4 => x110_out_3,
   O => W_39_7_i_15_n_0
);
W_39_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x110_out_3,
   I1 => x92_out_3,
   I2 => x108_out_21,
   I3 => x108_out_10,
   I4 => x108_out_6,
   O => W_39_7_i_16_n_0
);
W_39_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x92_out_2,
   I1 => x108_out_5,
   I2 => x108_out_9,
   I3 => x108_out_20,
   I4 => x110_out_2,
   O => W_39_7_i_17_n_0
);
W_39_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x77_out_16,
   I1 => x77_out_23,
   I2 => x77_out_25,
   I3 => W_39_7_i_10_n_0,
   I4 => W_39_7_i_11_n_0,
   O => W_39_7_i_2_n_0
);
W_39_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x77_out_15,
   I1 => x77_out_22,
   I2 => x77_out_24,
   I3 => W_39_7_i_12_n_0,
   I4 => W_39_7_i_13_n_0,
   O => W_39_7_i_3_n_0
);
W_39_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x77_out_14,
   I1 => x77_out_21,
   I2 => x77_out_23,
   I3 => W_39_7_i_14_n_0,
   I4 => W_39_7_i_15_n_0,
   O => W_39_7_i_4_n_0
);
W_39_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x77_out_13,
   I1 => x77_out_20,
   I2 => x77_out_22,
   I3 => W_39_7_i_16_n_0,
   I4 => W_39_7_i_17_n_0,
   O => W_39_7_i_5_n_0
);
W_39_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_39_7_i_2_n_0,
   I1 => W_39_11_i_16_n_0,
   I2 => x77_out_17,
   I3 => x77_out_24,
   I4 => x77_out_26,
   I5 => W_39_11_i_17_n_0,
   O => W_39_7_i_6_n_0
);
W_39_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_39_7_i_3_n_0,
   I1 => W_39_7_i_10_n_0,
   I2 => x77_out_16,
   I3 => x77_out_23,
   I4 => x77_out_25,
   I5 => W_39_7_i_11_n_0,
   O => W_39_7_i_7_n_0
);
W_39_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_39_7_i_4_n_0,
   I1 => W_39_7_i_12_n_0,
   I2 => x77_out_15,
   I3 => x77_out_22,
   I4 => x77_out_24,
   I5 => W_39_7_i_13_n_0,
   O => W_39_7_i_8_n_0
);
W_39_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_39_7_i_5_n_0,
   I1 => W_39_7_i_14_n_0,
   I2 => x77_out_14,
   I3 => x77_out_21,
   I4 => x77_out_23,
   I5 => W_39_7_i_15_n_0,
   O => W_39_7_i_9_n_0
);
W_40_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x108_out_10,
   I1 => x89_out_10,
   I2 => x106_out_28,
   I3 => x106_out_17,
   I4 => x106_out_13,
   O => W_40_11_i_10_n_0
);
W_40_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x89_out_9,
   I1 => x106_out_12,
   I2 => x106_out_16,
   I3 => x106_out_27,
   I4 => x108_out_9,
   O => W_40_11_i_11_n_0
);
W_40_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x108_out_9,
   I1 => x89_out_9,
   I2 => x106_out_27,
   I3 => x106_out_16,
   I4 => x106_out_12,
   O => W_40_11_i_12_n_0
);
W_40_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x89_out_8,
   I1 => x106_out_11,
   I2 => x106_out_15,
   I3 => x106_out_26,
   I4 => x108_out_8,
   O => W_40_11_i_13_n_0
);
W_40_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x108_out_8,
   I1 => x89_out_8,
   I2 => x106_out_26,
   I3 => x106_out_15,
   I4 => x106_out_11,
   O => W_40_11_i_14_n_0
);
W_40_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x89_out_7,
   I1 => x106_out_10,
   I2 => x106_out_14,
   I3 => x106_out_25,
   I4 => x108_out_7,
   O => W_40_11_i_15_n_0
);
W_40_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x108_out_7,
   I1 => x89_out_7,
   I2 => x106_out_25,
   I3 => x106_out_14,
   I4 => x106_out_10,
   O => W_40_11_i_16_n_0
);
W_40_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x89_out_6,
   I1 => x106_out_9,
   I2 => x106_out_13,
   I3 => x106_out_24,
   I4 => x108_out_6,
   O => W_40_11_i_17_n_0
);
W_40_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x74_out_20,
   I1 => x74_out_27,
   I2 => x74_out_29,
   I3 => W_40_11_i_10_n_0,
   I4 => W_40_11_i_11_n_0,
   O => W_40_11_i_2_n_0
);
W_40_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x74_out_19,
   I1 => x74_out_26,
   I2 => x74_out_28,
   I3 => W_40_11_i_12_n_0,
   I4 => W_40_11_i_13_n_0,
   O => W_40_11_i_3_n_0
);
W_40_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x74_out_18,
   I1 => x74_out_25,
   I2 => x74_out_27,
   I3 => W_40_11_i_14_n_0,
   I4 => W_40_11_i_15_n_0,
   O => W_40_11_i_4_n_0
);
W_40_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x74_out_17,
   I1 => x74_out_24,
   I2 => x74_out_26,
   I3 => W_40_11_i_16_n_0,
   I4 => W_40_11_i_17_n_0,
   O => W_40_11_i_5_n_0
);
W_40_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_40_11_i_2_n_0,
   I1 => W_40_15_i_16_n_0,
   I2 => x74_out_21,
   I3 => x74_out_28,
   I4 => x74_out_30,
   I5 => W_40_15_i_17_n_0,
   O => W_40_11_i_6_n_0
);
W_40_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_40_11_i_3_n_0,
   I1 => W_40_11_i_10_n_0,
   I2 => x74_out_20,
   I3 => x74_out_27,
   I4 => x74_out_29,
   I5 => W_40_11_i_11_n_0,
   O => W_40_11_i_7_n_0
);
W_40_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_40_11_i_4_n_0,
   I1 => W_40_11_i_12_n_0,
   I2 => x74_out_19,
   I3 => x74_out_26,
   I4 => x74_out_28,
   I5 => W_40_11_i_13_n_0,
   O => W_40_11_i_8_n_0
);
W_40_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_40_11_i_5_n_0,
   I1 => W_40_11_i_14_n_0,
   I2 => x74_out_18,
   I3 => x74_out_25,
   I4 => x74_out_27,
   I5 => W_40_11_i_15_n_0,
   O => W_40_11_i_9_n_0
);
W_40_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x108_out_14,
   I1 => x89_out_14,
   I2 => x106_out_0,
   I3 => x106_out_21,
   I4 => x106_out_17,
   O => W_40_15_i_10_n_0
);
W_40_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x89_out_13,
   I1 => x106_out_16,
   I2 => x106_out_20,
   I3 => x106_out_31,
   I4 => x108_out_13,
   O => W_40_15_i_11_n_0
);
W_40_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x108_out_13,
   I1 => x89_out_13,
   I2 => x106_out_31,
   I3 => x106_out_20,
   I4 => x106_out_16,
   O => W_40_15_i_12_n_0
);
W_40_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x89_out_12,
   I1 => x106_out_15,
   I2 => x106_out_19,
   I3 => x106_out_30,
   I4 => x108_out_12,
   O => W_40_15_i_13_n_0
);
W_40_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x108_out_12,
   I1 => x89_out_12,
   I2 => x106_out_30,
   I3 => x106_out_19,
   I4 => x106_out_15,
   O => W_40_15_i_14_n_0
);
W_40_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x89_out_11,
   I1 => x106_out_14,
   I2 => x106_out_18,
   I3 => x106_out_29,
   I4 => x108_out_11,
   O => W_40_15_i_15_n_0
);
W_40_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x108_out_11,
   I1 => x89_out_11,
   I2 => x106_out_29,
   I3 => x106_out_18,
   I4 => x106_out_14,
   O => W_40_15_i_16_n_0
);
W_40_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x89_out_10,
   I1 => x106_out_13,
   I2 => x106_out_17,
   I3 => x106_out_28,
   I4 => x108_out_10,
   O => W_40_15_i_17_n_0
);
W_40_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x74_out_24,
   I1 => x74_out_31,
   I2 => x74_out_1,
   I3 => W_40_15_i_10_n_0,
   I4 => W_40_15_i_11_n_0,
   O => W_40_15_i_2_n_0
);
W_40_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x74_out_23,
   I1 => x74_out_30,
   I2 => x74_out_0,
   I3 => W_40_15_i_12_n_0,
   I4 => W_40_15_i_13_n_0,
   O => W_40_15_i_3_n_0
);
W_40_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x74_out_22,
   I1 => x74_out_29,
   I2 => x74_out_31,
   I3 => W_40_15_i_14_n_0,
   I4 => W_40_15_i_15_n_0,
   O => W_40_15_i_4_n_0
);
W_40_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x74_out_21,
   I1 => x74_out_28,
   I2 => x74_out_30,
   I3 => W_40_15_i_16_n_0,
   I4 => W_40_15_i_17_n_0,
   O => W_40_15_i_5_n_0
);
W_40_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_40_15_i_2_n_0,
   I1 => W_40_19_i_16_n_0,
   I2 => x74_out_25,
   I3 => x74_out_0,
   I4 => x74_out_2,
   I5 => W_40_19_i_17_n_0,
   O => W_40_15_i_6_n_0
);
W_40_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_40_15_i_3_n_0,
   I1 => W_40_15_i_10_n_0,
   I2 => x74_out_24,
   I3 => x74_out_31,
   I4 => x74_out_1,
   I5 => W_40_15_i_11_n_0,
   O => W_40_15_i_7_n_0
);
W_40_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_40_15_i_4_n_0,
   I1 => W_40_15_i_12_n_0,
   I2 => x74_out_23,
   I3 => x74_out_30,
   I4 => x74_out_0,
   I5 => W_40_15_i_13_n_0,
   O => W_40_15_i_8_n_0
);
W_40_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_40_15_i_5_n_0,
   I1 => W_40_15_i_14_n_0,
   I2 => x74_out_22,
   I3 => x74_out_29,
   I4 => x74_out_31,
   I5 => W_40_15_i_15_n_0,
   O => W_40_15_i_9_n_0
);
W_40_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x108_out_18,
   I1 => x89_out_18,
   I2 => x106_out_4,
   I3 => x106_out_25,
   I4 => x106_out_21,
   O => W_40_19_i_10_n_0
);
W_40_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x89_out_17,
   I1 => x106_out_20,
   I2 => x106_out_24,
   I3 => x106_out_3,
   I4 => x108_out_17,
   O => W_40_19_i_11_n_0
);
W_40_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x108_out_17,
   I1 => x89_out_17,
   I2 => x106_out_3,
   I3 => x106_out_24,
   I4 => x106_out_20,
   O => W_40_19_i_12_n_0
);
W_40_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x89_out_16,
   I1 => x106_out_19,
   I2 => x106_out_23,
   I3 => x106_out_2,
   I4 => x108_out_16,
   O => W_40_19_i_13_n_0
);
W_40_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x108_out_16,
   I1 => x89_out_16,
   I2 => x106_out_2,
   I3 => x106_out_23,
   I4 => x106_out_19,
   O => W_40_19_i_14_n_0
);
W_40_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x89_out_15,
   I1 => x106_out_18,
   I2 => x106_out_22,
   I3 => x106_out_1,
   I4 => x108_out_15,
   O => W_40_19_i_15_n_0
);
W_40_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x108_out_15,
   I1 => x89_out_15,
   I2 => x106_out_1,
   I3 => x106_out_22,
   I4 => x106_out_18,
   O => W_40_19_i_16_n_0
);
W_40_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x89_out_14,
   I1 => x106_out_17,
   I2 => x106_out_21,
   I3 => x106_out_0,
   I4 => x108_out_14,
   O => W_40_19_i_17_n_0
);
W_40_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x74_out_28,
   I1 => x74_out_3,
   I2 => x74_out_5,
   I3 => W_40_19_i_10_n_0,
   I4 => W_40_19_i_11_n_0,
   O => W_40_19_i_2_n_0
);
W_40_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x74_out_27,
   I1 => x74_out_2,
   I2 => x74_out_4,
   I3 => W_40_19_i_12_n_0,
   I4 => W_40_19_i_13_n_0,
   O => W_40_19_i_3_n_0
);
W_40_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x74_out_26,
   I1 => x74_out_1,
   I2 => x74_out_3,
   I3 => W_40_19_i_14_n_0,
   I4 => W_40_19_i_15_n_0,
   O => W_40_19_i_4_n_0
);
W_40_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x74_out_25,
   I1 => x74_out_0,
   I2 => x74_out_2,
   I3 => W_40_19_i_16_n_0,
   I4 => W_40_19_i_17_n_0,
   O => W_40_19_i_5_n_0
);
W_40_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_40_19_i_2_n_0,
   I1 => W_40_23_i_16_n_0,
   I2 => x74_out_29,
   I3 => x74_out_4,
   I4 => x74_out_6,
   I5 => W_40_23_i_17_n_0,
   O => W_40_19_i_6_n_0
);
W_40_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_40_19_i_3_n_0,
   I1 => W_40_19_i_10_n_0,
   I2 => x74_out_28,
   I3 => x74_out_3,
   I4 => x74_out_5,
   I5 => W_40_19_i_11_n_0,
   O => W_40_19_i_7_n_0
);
W_40_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_40_19_i_4_n_0,
   I1 => W_40_19_i_12_n_0,
   I2 => x74_out_27,
   I3 => x74_out_2,
   I4 => x74_out_4,
   I5 => W_40_19_i_13_n_0,
   O => W_40_19_i_8_n_0
);
W_40_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_40_19_i_5_n_0,
   I1 => W_40_19_i_14_n_0,
   I2 => x74_out_26,
   I3 => x74_out_1,
   I4 => x74_out_3,
   I5 => W_40_19_i_15_n_0,
   O => W_40_19_i_9_n_0
);
W_40_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x108_out_22,
   I1 => x89_out_22,
   I2 => x106_out_8,
   I3 => x106_out_29,
   I4 => x106_out_25,
   O => W_40_23_i_10_n_0
);
W_40_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x89_out_21,
   I1 => x106_out_24,
   I2 => x106_out_28,
   I3 => x106_out_7,
   I4 => x108_out_21,
   O => W_40_23_i_11_n_0
);
W_40_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x108_out_21,
   I1 => x89_out_21,
   I2 => x106_out_7,
   I3 => x106_out_28,
   I4 => x106_out_24,
   O => W_40_23_i_12_n_0
);
W_40_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x89_out_20,
   I1 => x106_out_23,
   I2 => x106_out_27,
   I3 => x106_out_6,
   I4 => x108_out_20,
   O => W_40_23_i_13_n_0
);
W_40_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x108_out_20,
   I1 => x89_out_20,
   I2 => x106_out_6,
   I3 => x106_out_27,
   I4 => x106_out_23,
   O => W_40_23_i_14_n_0
);
W_40_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x89_out_19,
   I1 => x106_out_22,
   I2 => x106_out_26,
   I3 => x106_out_5,
   I4 => x108_out_19,
   O => W_40_23_i_15_n_0
);
W_40_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x108_out_19,
   I1 => x89_out_19,
   I2 => x106_out_5,
   I3 => x106_out_26,
   I4 => x106_out_22,
   O => W_40_23_i_16_n_0
);
W_40_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x89_out_18,
   I1 => x106_out_21,
   I2 => x106_out_25,
   I3 => x106_out_4,
   I4 => x108_out_18,
   O => W_40_23_i_17_n_0
);
W_40_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x74_out_7,
   I1 => x74_out_9,
   I2 => W_40_23_i_10_n_0,
   I3 => W_40_23_i_11_n_0,
   O => W_40_23_i_2_n_0
);
W_40_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x74_out_31,
   I1 => x74_out_6,
   I2 => x74_out_8,
   I3 => W_40_23_i_12_n_0,
   I4 => W_40_23_i_13_n_0,
   O => W_40_23_i_3_n_0
);
W_40_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x74_out_30,
   I1 => x74_out_5,
   I2 => x74_out_7,
   I3 => W_40_23_i_14_n_0,
   I4 => W_40_23_i_15_n_0,
   O => W_40_23_i_4_n_0
);
W_40_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x74_out_29,
   I1 => x74_out_4,
   I2 => x74_out_6,
   I3 => W_40_23_i_16_n_0,
   I4 => W_40_23_i_17_n_0,
   O => W_40_23_i_5_n_0
);
W_40_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x74_out_8,
   I1 => x74_out_10,
   I2 => W_40_27_i_16_n_0,
   I3 => W_40_27_i_17_n_0,
   I4 => W_40_23_i_2_n_0,
   O => W_40_23_i_6_n_0
);
W_40_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x74_out_7,
   I1 => x74_out_9,
   I2 => W_40_23_i_10_n_0,
   I3 => W_40_23_i_11_n_0,
   I4 => W_40_23_i_3_n_0,
   O => W_40_23_i_7_n_0
);
W_40_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_40_23_i_4_n_0,
   I1 => W_40_23_i_12_n_0,
   I2 => x74_out_31,
   I3 => x74_out_6,
   I4 => x74_out_8,
   I5 => W_40_23_i_13_n_0,
   O => W_40_23_i_8_n_0
);
W_40_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_40_23_i_5_n_0,
   I1 => W_40_23_i_14_n_0,
   I2 => x74_out_30,
   I3 => x74_out_5,
   I4 => x74_out_7,
   I5 => W_40_23_i_15_n_0,
   O => W_40_23_i_9_n_0
);
W_40_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x108_out_26,
   I1 => x89_out_26,
   I2 => x106_out_12,
   I3 => x106_out_1,
   I4 => x106_out_29,
   O => W_40_27_i_10_n_0
);
W_40_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x89_out_25,
   I1 => x106_out_28,
   I2 => x106_out_0,
   I3 => x106_out_11,
   I4 => x108_out_25,
   O => W_40_27_i_11_n_0
);
W_40_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x108_out_25,
   I1 => x89_out_25,
   I2 => x106_out_11,
   I3 => x106_out_0,
   I4 => x106_out_28,
   O => W_40_27_i_12_n_0
);
W_40_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x89_out_24,
   I1 => x106_out_27,
   I2 => x106_out_31,
   I3 => x106_out_10,
   I4 => x108_out_24,
   O => W_40_27_i_13_n_0
);
W_40_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x108_out_24,
   I1 => x89_out_24,
   I2 => x106_out_10,
   I3 => x106_out_31,
   I4 => x106_out_27,
   O => W_40_27_i_14_n_0
);
W_40_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x89_out_23,
   I1 => x106_out_26,
   I2 => x106_out_30,
   I3 => x106_out_9,
   I4 => x108_out_23,
   O => W_40_27_i_15_n_0
);
W_40_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x108_out_23,
   I1 => x89_out_23,
   I2 => x106_out_9,
   I3 => x106_out_30,
   I4 => x106_out_26,
   O => W_40_27_i_16_n_0
);
W_40_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x89_out_22,
   I1 => x106_out_25,
   I2 => x106_out_29,
   I3 => x106_out_8,
   I4 => x108_out_22,
   O => W_40_27_i_17_n_0
);
W_40_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x74_out_11,
   I1 => x74_out_13,
   I2 => W_40_27_i_10_n_0,
   I3 => W_40_27_i_11_n_0,
   O => W_40_27_i_2_n_0
);
W_40_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x74_out_10,
   I1 => x74_out_12,
   I2 => W_40_27_i_12_n_0,
   I3 => W_40_27_i_13_n_0,
   O => W_40_27_i_3_n_0
);
W_40_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x74_out_9,
   I1 => x74_out_11,
   I2 => W_40_27_i_14_n_0,
   I3 => W_40_27_i_15_n_0,
   O => W_40_27_i_4_n_0
);
W_40_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x74_out_8,
   I1 => x74_out_10,
   I2 => W_40_27_i_16_n_0,
   I3 => W_40_27_i_17_n_0,
   O => W_40_27_i_5_n_0
);
W_40_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x74_out_12,
   I1 => x74_out_14,
   I2 => W_40_31_i_13_n_0,
   I3 => W_40_31_i_14_n_0,
   I4 => W_40_27_i_2_n_0,
   O => W_40_27_i_6_n_0
);
W_40_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x74_out_11,
   I1 => x74_out_13,
   I2 => W_40_27_i_10_n_0,
   I3 => W_40_27_i_11_n_0,
   I4 => W_40_27_i_3_n_0,
   O => W_40_27_i_7_n_0
);
W_40_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x74_out_10,
   I1 => x74_out_12,
   I2 => W_40_27_i_12_n_0,
   I3 => W_40_27_i_13_n_0,
   I4 => W_40_27_i_4_n_0,
   O => W_40_27_i_8_n_0
);
W_40_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x74_out_9,
   I1 => x74_out_11,
   I2 => W_40_27_i_14_n_0,
   I3 => W_40_27_i_15_n_0,
   I4 => W_40_27_i_5_n_0,
   O => W_40_27_i_9_n_0
);
W_40_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x89_out_28,
   I1 => x106_out_31,
   I2 => x106_out_3,
   I3 => x106_out_14,
   I4 => x108_out_28,
   O => W_40_31_i_10_n_0
);
W_40_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x108_out_28,
   I1 => x89_out_28,
   I2 => x106_out_14,
   I3 => x106_out_3,
   I4 => x106_out_31,
   O => W_40_31_i_11_n_0
);
W_40_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x89_out_27,
   I1 => x106_out_30,
   I2 => x106_out_2,
   I3 => x106_out_13,
   I4 => x108_out_27,
   O => W_40_31_i_12_n_0
);
W_40_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x108_out_27,
   I1 => x89_out_27,
   I2 => x106_out_13,
   I3 => x106_out_2,
   I4 => x106_out_30,
   O => W_40_31_i_13_n_0
);
W_40_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x89_out_26,
   I1 => x106_out_29,
   I2 => x106_out_1,
   I3 => x106_out_12,
   I4 => x108_out_26,
   O => W_40_31_i_14_n_0
);
W_40_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x89_out_29,
   I1 => x106_out_4,
   I2 => x106_out_15,
   I3 => x108_out_29,
   O => W_40_31_i_15_n_0
);
W_40_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x74_out_17,
   I1 => x74_out_15,
   O => SIGMA_LCASE_1195_out_0_30
);
W_40_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => x106_out_6,
   I1 => x106_out_17,
   I2 => x89_out_31,
   I3 => x108_out_31,
   I4 => x74_out_16,
   I5 => x74_out_18,
   O => W_40_31_i_17_n_0
);
W_40_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x106_out_16,
   I1 => x106_out_5,
   O => SIGMA_LCASE_0191_out_30
);
W_40_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x108_out_30,
   I1 => x89_out_30,
   I2 => x106_out_16,
   I3 => x106_out_5,
   O => W_40_31_i_19_n_0
);
W_40_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x74_out_14,
   I1 => x74_out_16,
   I2 => W_40_31_i_9_n_0,
   I3 => W_40_31_i_10_n_0,
   O => W_40_31_i_2_n_0
);
W_40_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x74_out_13,
   I1 => x74_out_15,
   I2 => W_40_31_i_11_n_0,
   I3 => W_40_31_i_12_n_0,
   O => W_40_31_i_3_n_0
);
W_40_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x74_out_12,
   I1 => x74_out_14,
   I2 => W_40_31_i_13_n_0,
   I3 => W_40_31_i_14_n_0,
   O => W_40_31_i_4_n_0
);
W_40_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_40_31_i_15_n_0,
   I1 => SIGMA_LCASE_1195_out_0_30,
   I2 => W_40_31_i_17_n_0,
   I3 => x89_out_30,
   I4 => SIGMA_LCASE_0191_out_30,
   I5 => x108_out_30,
   O => W_40_31_i_5_n_0
);
W_40_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_40_31_i_2_n_0,
   I1 => W_40_31_i_19_n_0,
   I2 => x74_out_15,
   I3 => x74_out_17,
   I4 => W_40_31_i_15_n_0,
   O => W_40_31_i_6_n_0
);
W_40_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x74_out_14,
   I1 => x74_out_16,
   I2 => W_40_31_i_9_n_0,
   I3 => W_40_31_i_10_n_0,
   I4 => W_40_31_i_3_n_0,
   O => W_40_31_i_7_n_0
);
W_40_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x74_out_13,
   I1 => x74_out_15,
   I2 => W_40_31_i_11_n_0,
   I3 => W_40_31_i_12_n_0,
   I4 => W_40_31_i_4_n_0,
   O => W_40_31_i_8_n_0
);
W_40_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x108_out_29,
   I1 => x89_out_29,
   I2 => x106_out_15,
   I3 => x106_out_4,
   O => W_40_31_i_9_n_0
);
W_40_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x108_out_2,
   I1 => x89_out_2,
   I2 => x106_out_20,
   I3 => x106_out_9,
   I4 => x106_out_5,
   O => W_40_3_i_10_n_0
);
W_40_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x89_out_1,
   I1 => x106_out_4,
   I2 => x106_out_8,
   I3 => x106_out_19,
   I4 => x108_out_1,
   O => W_40_3_i_11_n_0
);
W_40_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x106_out_19,
   I1 => x106_out_8,
   I2 => x106_out_4,
   O => SIGMA_LCASE_0191_out_1
);
W_40_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x74_out_21,
   I1 => x74_out_19,
   I2 => x74_out_12,
   O => SIGMA_LCASE_1195_out_0_2
);
W_40_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x74_out_20,
   I1 => x74_out_18,
   I2 => x74_out_11,
   O => SIGMA_LCASE_1195_out_1
);
W_40_3_i_15 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x108_out_1,
   I1 => x89_out_1,
   I2 => x106_out_19,
   I3 => x106_out_8,
   I4 => x106_out_4,
   O => W_40_3_i_15_n_0
);
W_40_3_i_16 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x106_out_18,
   I1 => x106_out_7,
   I2 => x106_out_3,
   O => SIGMA_LCASE_0191_out_0
);
W_40_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x74_out_12,
   I1 => x74_out_19,
   I2 => x74_out_21,
   I3 => W_40_3_i_10_n_0,
   I4 => W_40_3_i_11_n_0,
   O => W_40_3_i_2_n_0
);
W_40_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_40_3_i_11_n_0,
   I1 => x74_out_21,
   I2 => x74_out_19,
   I3 => x74_out_12,
   I4 => W_40_3_i_10_n_0,
   O => W_40_3_i_3_n_0
);
W_40_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_0191_out_1,
   I1 => x89_out_1,
   I2 => x108_out_1,
   I3 => x74_out_11,
   I4 => x74_out_18,
   I5 => x74_out_20,
   O => W_40_3_i_4_n_0
);
W_40_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x108_out_0,
   I1 => x89_out_0,
   I2 => x106_out_18,
   I3 => x106_out_7,
   I4 => x106_out_3,
   O => W_40_3_i_5_n_0
);
W_40_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_40_3_i_2_n_0,
   I1 => W_40_7_i_16_n_0,
   I2 => x74_out_13,
   I3 => x74_out_20,
   I4 => x74_out_22,
   I5 => W_40_7_i_17_n_0,
   O => W_40_3_i_6_n_0
);
W_40_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_40_3_i_10_n_0,
   I1 => SIGMA_LCASE_1195_out_0_2,
   I2 => x108_out_1,
   I3 => x89_out_1,
   I4 => SIGMA_LCASE_0191_out_1,
   I5 => SIGMA_LCASE_1195_out_1,
   O => W_40_3_i_7_n_0
);
W_40_3_i_8 : LUT5
  generic map(
   INIT => X"99969666"
  )
 port map (
   I0 => SIGMA_LCASE_1195_out_1,
   I1 => W_40_3_i_15_n_0,
   I2 => x108_out_0,
   I3 => SIGMA_LCASE_0191_out_0,
   I4 => x89_out_0,
   O => W_40_3_i_8_n_0
);
W_40_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_40_3_i_5_n_0,
   I1 => x74_out_10,
   I2 => x74_out_17,
   I3 => x74_out_19,
   O => W_40_3_i_9_n_0
);
W_40_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x108_out_6,
   I1 => x89_out_6,
   I2 => x106_out_24,
   I3 => x106_out_13,
   I4 => x106_out_9,
   O => W_40_7_i_10_n_0
);
W_40_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x89_out_5,
   I1 => x106_out_8,
   I2 => x106_out_12,
   I3 => x106_out_23,
   I4 => x108_out_5,
   O => W_40_7_i_11_n_0
);
W_40_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x108_out_5,
   I1 => x89_out_5,
   I2 => x106_out_23,
   I3 => x106_out_12,
   I4 => x106_out_8,
   O => W_40_7_i_12_n_0
);
W_40_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x89_out_4,
   I1 => x106_out_7,
   I2 => x106_out_11,
   I3 => x106_out_22,
   I4 => x108_out_4,
   O => W_40_7_i_13_n_0
);
W_40_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x108_out_4,
   I1 => x89_out_4,
   I2 => x106_out_22,
   I3 => x106_out_11,
   I4 => x106_out_7,
   O => W_40_7_i_14_n_0
);
W_40_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x89_out_3,
   I1 => x106_out_6,
   I2 => x106_out_10,
   I3 => x106_out_21,
   I4 => x108_out_3,
   O => W_40_7_i_15_n_0
);
W_40_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x108_out_3,
   I1 => x89_out_3,
   I2 => x106_out_21,
   I3 => x106_out_10,
   I4 => x106_out_6,
   O => W_40_7_i_16_n_0
);
W_40_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x89_out_2,
   I1 => x106_out_5,
   I2 => x106_out_9,
   I3 => x106_out_20,
   I4 => x108_out_2,
   O => W_40_7_i_17_n_0
);
W_40_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x74_out_16,
   I1 => x74_out_23,
   I2 => x74_out_25,
   I3 => W_40_7_i_10_n_0,
   I4 => W_40_7_i_11_n_0,
   O => W_40_7_i_2_n_0
);
W_40_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x74_out_15,
   I1 => x74_out_22,
   I2 => x74_out_24,
   I3 => W_40_7_i_12_n_0,
   I4 => W_40_7_i_13_n_0,
   O => W_40_7_i_3_n_0
);
W_40_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x74_out_14,
   I1 => x74_out_21,
   I2 => x74_out_23,
   I3 => W_40_7_i_14_n_0,
   I4 => W_40_7_i_15_n_0,
   O => W_40_7_i_4_n_0
);
W_40_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x74_out_13,
   I1 => x74_out_20,
   I2 => x74_out_22,
   I3 => W_40_7_i_16_n_0,
   I4 => W_40_7_i_17_n_0,
   O => W_40_7_i_5_n_0
);
W_40_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_40_7_i_2_n_0,
   I1 => W_40_11_i_16_n_0,
   I2 => x74_out_17,
   I3 => x74_out_24,
   I4 => x74_out_26,
   I5 => W_40_11_i_17_n_0,
   O => W_40_7_i_6_n_0
);
W_40_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_40_7_i_3_n_0,
   I1 => W_40_7_i_10_n_0,
   I2 => x74_out_16,
   I3 => x74_out_23,
   I4 => x74_out_25,
   I5 => W_40_7_i_11_n_0,
   O => W_40_7_i_7_n_0
);
W_40_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_40_7_i_4_n_0,
   I1 => W_40_7_i_12_n_0,
   I2 => x74_out_15,
   I3 => x74_out_22,
   I4 => x74_out_24,
   I5 => W_40_7_i_13_n_0,
   O => W_40_7_i_8_n_0
);
W_40_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_40_7_i_5_n_0,
   I1 => W_40_7_i_14_n_0,
   I2 => x74_out_14,
   I3 => x74_out_21,
   I4 => x74_out_23,
   I5 => W_40_7_i_15_n_0,
   O => W_40_7_i_9_n_0
);
W_41_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x106_out_10,
   I1 => x86_out_10,
   I2 => x104_out_28,
   I3 => x104_out_17,
   I4 => x104_out_13,
   O => W_41_11_i_10_n_0
);
W_41_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x86_out_9,
   I1 => x104_out_12,
   I2 => x104_out_16,
   I3 => x104_out_27,
   I4 => x106_out_9,
   O => W_41_11_i_11_n_0
);
W_41_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x106_out_9,
   I1 => x86_out_9,
   I2 => x104_out_27,
   I3 => x104_out_16,
   I4 => x104_out_12,
   O => W_41_11_i_12_n_0
);
W_41_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x86_out_8,
   I1 => x104_out_11,
   I2 => x104_out_15,
   I3 => x104_out_26,
   I4 => x106_out_8,
   O => W_41_11_i_13_n_0
);
W_41_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x106_out_8,
   I1 => x86_out_8,
   I2 => x104_out_26,
   I3 => x104_out_15,
   I4 => x104_out_11,
   O => W_41_11_i_14_n_0
);
W_41_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x86_out_7,
   I1 => x104_out_10,
   I2 => x104_out_14,
   I3 => x104_out_25,
   I4 => x106_out_7,
   O => W_41_11_i_15_n_0
);
W_41_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x106_out_7,
   I1 => x86_out_7,
   I2 => x104_out_25,
   I3 => x104_out_14,
   I4 => x104_out_10,
   O => W_41_11_i_16_n_0
);
W_41_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x86_out_6,
   I1 => x104_out_9,
   I2 => x104_out_13,
   I3 => x104_out_24,
   I4 => x106_out_6,
   O => W_41_11_i_17_n_0
);
W_41_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x71_out_20,
   I1 => x71_out_27,
   I2 => x71_out_29,
   I3 => W_41_11_i_10_n_0,
   I4 => W_41_11_i_11_n_0,
   O => W_41_11_i_2_n_0
);
W_41_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x71_out_19,
   I1 => x71_out_26,
   I2 => x71_out_28,
   I3 => W_41_11_i_12_n_0,
   I4 => W_41_11_i_13_n_0,
   O => W_41_11_i_3_n_0
);
W_41_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x71_out_18,
   I1 => x71_out_25,
   I2 => x71_out_27,
   I3 => W_41_11_i_14_n_0,
   I4 => W_41_11_i_15_n_0,
   O => W_41_11_i_4_n_0
);
W_41_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x71_out_17,
   I1 => x71_out_24,
   I2 => x71_out_26,
   I3 => W_41_11_i_16_n_0,
   I4 => W_41_11_i_17_n_0,
   O => W_41_11_i_5_n_0
);
W_41_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_41_11_i_2_n_0,
   I1 => W_41_15_i_16_n_0,
   I2 => x71_out_21,
   I3 => x71_out_28,
   I4 => x71_out_30,
   I5 => W_41_15_i_17_n_0,
   O => W_41_11_i_6_n_0
);
W_41_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_41_11_i_3_n_0,
   I1 => W_41_11_i_10_n_0,
   I2 => x71_out_20,
   I3 => x71_out_27,
   I4 => x71_out_29,
   I5 => W_41_11_i_11_n_0,
   O => W_41_11_i_7_n_0
);
W_41_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_41_11_i_4_n_0,
   I1 => W_41_11_i_12_n_0,
   I2 => x71_out_19,
   I3 => x71_out_26,
   I4 => x71_out_28,
   I5 => W_41_11_i_13_n_0,
   O => W_41_11_i_8_n_0
);
W_41_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_41_11_i_5_n_0,
   I1 => W_41_11_i_14_n_0,
   I2 => x71_out_18,
   I3 => x71_out_25,
   I4 => x71_out_27,
   I5 => W_41_11_i_15_n_0,
   O => W_41_11_i_9_n_0
);
W_41_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x106_out_14,
   I1 => x86_out_14,
   I2 => x104_out_0,
   I3 => x104_out_21,
   I4 => x104_out_17,
   O => W_41_15_i_10_n_0
);
W_41_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x86_out_13,
   I1 => x104_out_16,
   I2 => x104_out_20,
   I3 => x104_out_31,
   I4 => x106_out_13,
   O => W_41_15_i_11_n_0
);
W_41_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x106_out_13,
   I1 => x86_out_13,
   I2 => x104_out_31,
   I3 => x104_out_20,
   I4 => x104_out_16,
   O => W_41_15_i_12_n_0
);
W_41_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x86_out_12,
   I1 => x104_out_15,
   I2 => x104_out_19,
   I3 => x104_out_30,
   I4 => x106_out_12,
   O => W_41_15_i_13_n_0
);
W_41_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x106_out_12,
   I1 => x86_out_12,
   I2 => x104_out_30,
   I3 => x104_out_19,
   I4 => x104_out_15,
   O => W_41_15_i_14_n_0
);
W_41_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x86_out_11,
   I1 => x104_out_14,
   I2 => x104_out_18,
   I3 => x104_out_29,
   I4 => x106_out_11,
   O => W_41_15_i_15_n_0
);
W_41_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x106_out_11,
   I1 => x86_out_11,
   I2 => x104_out_29,
   I3 => x104_out_18,
   I4 => x104_out_14,
   O => W_41_15_i_16_n_0
);
W_41_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x86_out_10,
   I1 => x104_out_13,
   I2 => x104_out_17,
   I3 => x104_out_28,
   I4 => x106_out_10,
   O => W_41_15_i_17_n_0
);
W_41_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x71_out_24,
   I1 => x71_out_31,
   I2 => x71_out_1,
   I3 => W_41_15_i_10_n_0,
   I4 => W_41_15_i_11_n_0,
   O => W_41_15_i_2_n_0
);
W_41_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x71_out_23,
   I1 => x71_out_30,
   I2 => x71_out_0,
   I3 => W_41_15_i_12_n_0,
   I4 => W_41_15_i_13_n_0,
   O => W_41_15_i_3_n_0
);
W_41_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x71_out_22,
   I1 => x71_out_29,
   I2 => x71_out_31,
   I3 => W_41_15_i_14_n_0,
   I4 => W_41_15_i_15_n_0,
   O => W_41_15_i_4_n_0
);
W_41_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x71_out_21,
   I1 => x71_out_28,
   I2 => x71_out_30,
   I3 => W_41_15_i_16_n_0,
   I4 => W_41_15_i_17_n_0,
   O => W_41_15_i_5_n_0
);
W_41_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_41_15_i_2_n_0,
   I1 => W_41_19_i_16_n_0,
   I2 => x71_out_25,
   I3 => x71_out_0,
   I4 => x71_out_2,
   I5 => W_41_19_i_17_n_0,
   O => W_41_15_i_6_n_0
);
W_41_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_41_15_i_3_n_0,
   I1 => W_41_15_i_10_n_0,
   I2 => x71_out_24,
   I3 => x71_out_31,
   I4 => x71_out_1,
   I5 => W_41_15_i_11_n_0,
   O => W_41_15_i_7_n_0
);
W_41_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_41_15_i_4_n_0,
   I1 => W_41_15_i_12_n_0,
   I2 => x71_out_23,
   I3 => x71_out_30,
   I4 => x71_out_0,
   I5 => W_41_15_i_13_n_0,
   O => W_41_15_i_8_n_0
);
W_41_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_41_15_i_5_n_0,
   I1 => W_41_15_i_14_n_0,
   I2 => x71_out_22,
   I3 => x71_out_29,
   I4 => x71_out_31,
   I5 => W_41_15_i_15_n_0,
   O => W_41_15_i_9_n_0
);
W_41_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x106_out_18,
   I1 => x86_out_18,
   I2 => x104_out_4,
   I3 => x104_out_25,
   I4 => x104_out_21,
   O => W_41_19_i_10_n_0
);
W_41_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x86_out_17,
   I1 => x104_out_20,
   I2 => x104_out_24,
   I3 => x104_out_3,
   I4 => x106_out_17,
   O => W_41_19_i_11_n_0
);
W_41_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x106_out_17,
   I1 => x86_out_17,
   I2 => x104_out_3,
   I3 => x104_out_24,
   I4 => x104_out_20,
   O => W_41_19_i_12_n_0
);
W_41_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x86_out_16,
   I1 => x104_out_19,
   I2 => x104_out_23,
   I3 => x104_out_2,
   I4 => x106_out_16,
   O => W_41_19_i_13_n_0
);
W_41_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x106_out_16,
   I1 => x86_out_16,
   I2 => x104_out_2,
   I3 => x104_out_23,
   I4 => x104_out_19,
   O => W_41_19_i_14_n_0
);
W_41_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x86_out_15,
   I1 => x104_out_18,
   I2 => x104_out_22,
   I3 => x104_out_1,
   I4 => x106_out_15,
   O => W_41_19_i_15_n_0
);
W_41_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x106_out_15,
   I1 => x86_out_15,
   I2 => x104_out_1,
   I3 => x104_out_22,
   I4 => x104_out_18,
   O => W_41_19_i_16_n_0
);
W_41_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x86_out_14,
   I1 => x104_out_17,
   I2 => x104_out_21,
   I3 => x104_out_0,
   I4 => x106_out_14,
   O => W_41_19_i_17_n_0
);
W_41_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x71_out_28,
   I1 => x71_out_3,
   I2 => x71_out_5,
   I3 => W_41_19_i_10_n_0,
   I4 => W_41_19_i_11_n_0,
   O => W_41_19_i_2_n_0
);
W_41_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x71_out_27,
   I1 => x71_out_2,
   I2 => x71_out_4,
   I3 => W_41_19_i_12_n_0,
   I4 => W_41_19_i_13_n_0,
   O => W_41_19_i_3_n_0
);
W_41_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x71_out_26,
   I1 => x71_out_1,
   I2 => x71_out_3,
   I3 => W_41_19_i_14_n_0,
   I4 => W_41_19_i_15_n_0,
   O => W_41_19_i_4_n_0
);
W_41_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x71_out_25,
   I1 => x71_out_0,
   I2 => x71_out_2,
   I3 => W_41_19_i_16_n_0,
   I4 => W_41_19_i_17_n_0,
   O => W_41_19_i_5_n_0
);
W_41_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_41_19_i_2_n_0,
   I1 => W_41_23_i_16_n_0,
   I2 => x71_out_29,
   I3 => x71_out_4,
   I4 => x71_out_6,
   I5 => W_41_23_i_17_n_0,
   O => W_41_19_i_6_n_0
);
W_41_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_41_19_i_3_n_0,
   I1 => W_41_19_i_10_n_0,
   I2 => x71_out_28,
   I3 => x71_out_3,
   I4 => x71_out_5,
   I5 => W_41_19_i_11_n_0,
   O => W_41_19_i_7_n_0
);
W_41_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_41_19_i_4_n_0,
   I1 => W_41_19_i_12_n_0,
   I2 => x71_out_27,
   I3 => x71_out_2,
   I4 => x71_out_4,
   I5 => W_41_19_i_13_n_0,
   O => W_41_19_i_8_n_0
);
W_41_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_41_19_i_5_n_0,
   I1 => W_41_19_i_14_n_0,
   I2 => x71_out_26,
   I3 => x71_out_1,
   I4 => x71_out_3,
   I5 => W_41_19_i_15_n_0,
   O => W_41_19_i_9_n_0
);
W_41_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x106_out_22,
   I1 => x86_out_22,
   I2 => x104_out_8,
   I3 => x104_out_29,
   I4 => x104_out_25,
   O => W_41_23_i_10_n_0
);
W_41_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x86_out_21,
   I1 => x104_out_24,
   I2 => x104_out_28,
   I3 => x104_out_7,
   I4 => x106_out_21,
   O => W_41_23_i_11_n_0
);
W_41_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x106_out_21,
   I1 => x86_out_21,
   I2 => x104_out_7,
   I3 => x104_out_28,
   I4 => x104_out_24,
   O => W_41_23_i_12_n_0
);
W_41_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x86_out_20,
   I1 => x104_out_23,
   I2 => x104_out_27,
   I3 => x104_out_6,
   I4 => x106_out_20,
   O => W_41_23_i_13_n_0
);
W_41_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x106_out_20,
   I1 => x86_out_20,
   I2 => x104_out_6,
   I3 => x104_out_27,
   I4 => x104_out_23,
   O => W_41_23_i_14_n_0
);
W_41_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x86_out_19,
   I1 => x104_out_22,
   I2 => x104_out_26,
   I3 => x104_out_5,
   I4 => x106_out_19,
   O => W_41_23_i_15_n_0
);
W_41_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x106_out_19,
   I1 => x86_out_19,
   I2 => x104_out_5,
   I3 => x104_out_26,
   I4 => x104_out_22,
   O => W_41_23_i_16_n_0
);
W_41_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x86_out_18,
   I1 => x104_out_21,
   I2 => x104_out_25,
   I3 => x104_out_4,
   I4 => x106_out_18,
   O => W_41_23_i_17_n_0
);
W_41_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x71_out_7,
   I1 => x71_out_9,
   I2 => W_41_23_i_10_n_0,
   I3 => W_41_23_i_11_n_0,
   O => W_41_23_i_2_n_0
);
W_41_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x71_out_31,
   I1 => x71_out_6,
   I2 => x71_out_8,
   I3 => W_41_23_i_12_n_0,
   I4 => W_41_23_i_13_n_0,
   O => W_41_23_i_3_n_0
);
W_41_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x71_out_30,
   I1 => x71_out_5,
   I2 => x71_out_7,
   I3 => W_41_23_i_14_n_0,
   I4 => W_41_23_i_15_n_0,
   O => W_41_23_i_4_n_0
);
W_41_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x71_out_29,
   I1 => x71_out_4,
   I2 => x71_out_6,
   I3 => W_41_23_i_16_n_0,
   I4 => W_41_23_i_17_n_0,
   O => W_41_23_i_5_n_0
);
W_41_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x71_out_8,
   I1 => x71_out_10,
   I2 => W_41_27_i_16_n_0,
   I3 => W_41_27_i_17_n_0,
   I4 => W_41_23_i_2_n_0,
   O => W_41_23_i_6_n_0
);
W_41_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x71_out_7,
   I1 => x71_out_9,
   I2 => W_41_23_i_10_n_0,
   I3 => W_41_23_i_11_n_0,
   I4 => W_41_23_i_3_n_0,
   O => W_41_23_i_7_n_0
);
W_41_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_41_23_i_4_n_0,
   I1 => W_41_23_i_12_n_0,
   I2 => x71_out_31,
   I3 => x71_out_6,
   I4 => x71_out_8,
   I5 => W_41_23_i_13_n_0,
   O => W_41_23_i_8_n_0
);
W_41_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_41_23_i_5_n_0,
   I1 => W_41_23_i_14_n_0,
   I2 => x71_out_30,
   I3 => x71_out_5,
   I4 => x71_out_7,
   I5 => W_41_23_i_15_n_0,
   O => W_41_23_i_9_n_0
);
W_41_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x106_out_26,
   I1 => x86_out_26,
   I2 => x104_out_12,
   I3 => x104_out_1,
   I4 => x104_out_29,
   O => W_41_27_i_10_n_0
);
W_41_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x86_out_25,
   I1 => x104_out_28,
   I2 => x104_out_0,
   I3 => x104_out_11,
   I4 => x106_out_25,
   O => W_41_27_i_11_n_0
);
W_41_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x106_out_25,
   I1 => x86_out_25,
   I2 => x104_out_11,
   I3 => x104_out_0,
   I4 => x104_out_28,
   O => W_41_27_i_12_n_0
);
W_41_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x86_out_24,
   I1 => x104_out_27,
   I2 => x104_out_31,
   I3 => x104_out_10,
   I4 => x106_out_24,
   O => W_41_27_i_13_n_0
);
W_41_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x106_out_24,
   I1 => x86_out_24,
   I2 => x104_out_10,
   I3 => x104_out_31,
   I4 => x104_out_27,
   O => W_41_27_i_14_n_0
);
W_41_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x86_out_23,
   I1 => x104_out_26,
   I2 => x104_out_30,
   I3 => x104_out_9,
   I4 => x106_out_23,
   O => W_41_27_i_15_n_0
);
W_41_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x106_out_23,
   I1 => x86_out_23,
   I2 => x104_out_9,
   I3 => x104_out_30,
   I4 => x104_out_26,
   O => W_41_27_i_16_n_0
);
W_41_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x86_out_22,
   I1 => x104_out_25,
   I2 => x104_out_29,
   I3 => x104_out_8,
   I4 => x106_out_22,
   O => W_41_27_i_17_n_0
);
W_41_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x71_out_11,
   I1 => x71_out_13,
   I2 => W_41_27_i_10_n_0,
   I3 => W_41_27_i_11_n_0,
   O => W_41_27_i_2_n_0
);
W_41_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x71_out_10,
   I1 => x71_out_12,
   I2 => W_41_27_i_12_n_0,
   I3 => W_41_27_i_13_n_0,
   O => W_41_27_i_3_n_0
);
W_41_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x71_out_9,
   I1 => x71_out_11,
   I2 => W_41_27_i_14_n_0,
   I3 => W_41_27_i_15_n_0,
   O => W_41_27_i_4_n_0
);
W_41_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x71_out_8,
   I1 => x71_out_10,
   I2 => W_41_27_i_16_n_0,
   I3 => W_41_27_i_17_n_0,
   O => W_41_27_i_5_n_0
);
W_41_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x71_out_12,
   I1 => x71_out_14,
   I2 => W_41_31_i_13_n_0,
   I3 => W_41_31_i_14_n_0,
   I4 => W_41_27_i_2_n_0,
   O => W_41_27_i_6_n_0
);
W_41_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x71_out_11,
   I1 => x71_out_13,
   I2 => W_41_27_i_10_n_0,
   I3 => W_41_27_i_11_n_0,
   I4 => W_41_27_i_3_n_0,
   O => W_41_27_i_7_n_0
);
W_41_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x71_out_10,
   I1 => x71_out_12,
   I2 => W_41_27_i_12_n_0,
   I3 => W_41_27_i_13_n_0,
   I4 => W_41_27_i_4_n_0,
   O => W_41_27_i_8_n_0
);
W_41_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x71_out_9,
   I1 => x71_out_11,
   I2 => W_41_27_i_14_n_0,
   I3 => W_41_27_i_15_n_0,
   I4 => W_41_27_i_5_n_0,
   O => W_41_27_i_9_n_0
);
W_41_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x86_out_28,
   I1 => x104_out_31,
   I2 => x104_out_3,
   I3 => x104_out_14,
   I4 => x106_out_28,
   O => W_41_31_i_10_n_0
);
W_41_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x106_out_28,
   I1 => x86_out_28,
   I2 => x104_out_14,
   I3 => x104_out_3,
   I4 => x104_out_31,
   O => W_41_31_i_11_n_0
);
W_41_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x86_out_27,
   I1 => x104_out_30,
   I2 => x104_out_2,
   I3 => x104_out_13,
   I4 => x106_out_27,
   O => W_41_31_i_12_n_0
);
W_41_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x106_out_27,
   I1 => x86_out_27,
   I2 => x104_out_13,
   I3 => x104_out_2,
   I4 => x104_out_30,
   O => W_41_31_i_13_n_0
);
W_41_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x86_out_26,
   I1 => x104_out_29,
   I2 => x104_out_1,
   I3 => x104_out_12,
   I4 => x106_out_26,
   O => W_41_31_i_14_n_0
);
W_41_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x86_out_29,
   I1 => x104_out_4,
   I2 => x104_out_15,
   I3 => x106_out_29,
   O => W_41_31_i_15_n_0
);
W_41_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x71_out_17,
   I1 => x71_out_15,
   O => SIGMA_LCASE_1187_out_0_30
);
W_41_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => x104_out_6,
   I1 => x104_out_17,
   I2 => x86_out_31,
   I3 => x106_out_31,
   I4 => x71_out_16,
   I5 => x71_out_18,
   O => W_41_31_i_17_n_0
);
W_41_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x104_out_16,
   I1 => x104_out_5,
   O => SIGMA_LCASE_0183_out_30
);
W_41_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x106_out_30,
   I1 => x86_out_30,
   I2 => x104_out_16,
   I3 => x104_out_5,
   O => W_41_31_i_19_n_0
);
W_41_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x71_out_14,
   I1 => x71_out_16,
   I2 => W_41_31_i_9_n_0,
   I3 => W_41_31_i_10_n_0,
   O => W_41_31_i_2_n_0
);
W_41_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x71_out_13,
   I1 => x71_out_15,
   I2 => W_41_31_i_11_n_0,
   I3 => W_41_31_i_12_n_0,
   O => W_41_31_i_3_n_0
);
W_41_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x71_out_12,
   I1 => x71_out_14,
   I2 => W_41_31_i_13_n_0,
   I3 => W_41_31_i_14_n_0,
   O => W_41_31_i_4_n_0
);
W_41_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_41_31_i_15_n_0,
   I1 => SIGMA_LCASE_1187_out_0_30,
   I2 => W_41_31_i_17_n_0,
   I3 => x86_out_30,
   I4 => SIGMA_LCASE_0183_out_30,
   I5 => x106_out_30,
   O => W_41_31_i_5_n_0
);
W_41_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_41_31_i_2_n_0,
   I1 => W_41_31_i_19_n_0,
   I2 => x71_out_15,
   I3 => x71_out_17,
   I4 => W_41_31_i_15_n_0,
   O => W_41_31_i_6_n_0
);
W_41_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x71_out_14,
   I1 => x71_out_16,
   I2 => W_41_31_i_9_n_0,
   I3 => W_41_31_i_10_n_0,
   I4 => W_41_31_i_3_n_0,
   O => W_41_31_i_7_n_0
);
W_41_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x71_out_13,
   I1 => x71_out_15,
   I2 => W_41_31_i_11_n_0,
   I3 => W_41_31_i_12_n_0,
   I4 => W_41_31_i_4_n_0,
   O => W_41_31_i_8_n_0
);
W_41_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x106_out_29,
   I1 => x86_out_29,
   I2 => x104_out_15,
   I3 => x104_out_4,
   O => W_41_31_i_9_n_0
);
W_41_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x106_out_2,
   I1 => x86_out_2,
   I2 => x104_out_20,
   I3 => x104_out_9,
   I4 => x104_out_5,
   O => W_41_3_i_10_n_0
);
W_41_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x86_out_1,
   I1 => x104_out_4,
   I2 => x104_out_8,
   I3 => x104_out_19,
   I4 => x106_out_1,
   O => W_41_3_i_11_n_0
);
W_41_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x104_out_19,
   I1 => x104_out_8,
   I2 => x104_out_4,
   O => SIGMA_LCASE_0183_out_1
);
W_41_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x71_out_21,
   I1 => x71_out_19,
   I2 => x71_out_12,
   O => SIGMA_LCASE_1187_out_0_2
);
W_41_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x71_out_20,
   I1 => x71_out_18,
   I2 => x71_out_11,
   O => SIGMA_LCASE_1187_out_1
);
W_41_3_i_15 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x106_out_1,
   I1 => x86_out_1,
   I2 => x104_out_19,
   I3 => x104_out_8,
   I4 => x104_out_4,
   O => W_41_3_i_15_n_0
);
W_41_3_i_16 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x104_out_18,
   I1 => x104_out_7,
   I2 => x104_out_3,
   O => SIGMA_LCASE_0183_out_0
);
W_41_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x71_out_12,
   I1 => x71_out_19,
   I2 => x71_out_21,
   I3 => W_41_3_i_10_n_0,
   I4 => W_41_3_i_11_n_0,
   O => W_41_3_i_2_n_0
);
W_41_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_41_3_i_11_n_0,
   I1 => x71_out_21,
   I2 => x71_out_19,
   I3 => x71_out_12,
   I4 => W_41_3_i_10_n_0,
   O => W_41_3_i_3_n_0
);
W_41_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_0183_out_1,
   I1 => x86_out_1,
   I2 => x106_out_1,
   I3 => x71_out_11,
   I4 => x71_out_18,
   I5 => x71_out_20,
   O => W_41_3_i_4_n_0
);
W_41_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x106_out_0,
   I1 => x86_out_0,
   I2 => x104_out_18,
   I3 => x104_out_7,
   I4 => x104_out_3,
   O => W_41_3_i_5_n_0
);
W_41_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_41_3_i_2_n_0,
   I1 => W_41_7_i_16_n_0,
   I2 => x71_out_13,
   I3 => x71_out_20,
   I4 => x71_out_22,
   I5 => W_41_7_i_17_n_0,
   O => W_41_3_i_6_n_0
);
W_41_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_41_3_i_10_n_0,
   I1 => SIGMA_LCASE_1187_out_0_2,
   I2 => x106_out_1,
   I3 => x86_out_1,
   I4 => SIGMA_LCASE_0183_out_1,
   I5 => SIGMA_LCASE_1187_out_1,
   O => W_41_3_i_7_n_0
);
W_41_3_i_8 : LUT5
  generic map(
   INIT => X"99969666"
  )
 port map (
   I0 => SIGMA_LCASE_1187_out_1,
   I1 => W_41_3_i_15_n_0,
   I2 => x106_out_0,
   I3 => SIGMA_LCASE_0183_out_0,
   I4 => x86_out_0,
   O => W_41_3_i_8_n_0
);
W_41_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_41_3_i_5_n_0,
   I1 => x71_out_10,
   I2 => x71_out_17,
   I3 => x71_out_19,
   O => W_41_3_i_9_n_0
);
W_41_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x106_out_6,
   I1 => x86_out_6,
   I2 => x104_out_24,
   I3 => x104_out_13,
   I4 => x104_out_9,
   O => W_41_7_i_10_n_0
);
W_41_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x86_out_5,
   I1 => x104_out_8,
   I2 => x104_out_12,
   I3 => x104_out_23,
   I4 => x106_out_5,
   O => W_41_7_i_11_n_0
);
W_41_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x106_out_5,
   I1 => x86_out_5,
   I2 => x104_out_23,
   I3 => x104_out_12,
   I4 => x104_out_8,
   O => W_41_7_i_12_n_0
);
W_41_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x86_out_4,
   I1 => x104_out_7,
   I2 => x104_out_11,
   I3 => x104_out_22,
   I4 => x106_out_4,
   O => W_41_7_i_13_n_0
);
W_41_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x106_out_4,
   I1 => x86_out_4,
   I2 => x104_out_22,
   I3 => x104_out_11,
   I4 => x104_out_7,
   O => W_41_7_i_14_n_0
);
W_41_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x86_out_3,
   I1 => x104_out_6,
   I2 => x104_out_10,
   I3 => x104_out_21,
   I4 => x106_out_3,
   O => W_41_7_i_15_n_0
);
W_41_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x106_out_3,
   I1 => x86_out_3,
   I2 => x104_out_21,
   I3 => x104_out_10,
   I4 => x104_out_6,
   O => W_41_7_i_16_n_0
);
W_41_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x86_out_2,
   I1 => x104_out_5,
   I2 => x104_out_9,
   I3 => x104_out_20,
   I4 => x106_out_2,
   O => W_41_7_i_17_n_0
);
W_41_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x71_out_16,
   I1 => x71_out_23,
   I2 => x71_out_25,
   I3 => W_41_7_i_10_n_0,
   I4 => W_41_7_i_11_n_0,
   O => W_41_7_i_2_n_0
);
W_41_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x71_out_15,
   I1 => x71_out_22,
   I2 => x71_out_24,
   I3 => W_41_7_i_12_n_0,
   I4 => W_41_7_i_13_n_0,
   O => W_41_7_i_3_n_0
);
W_41_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x71_out_14,
   I1 => x71_out_21,
   I2 => x71_out_23,
   I3 => W_41_7_i_14_n_0,
   I4 => W_41_7_i_15_n_0,
   O => W_41_7_i_4_n_0
);
W_41_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x71_out_13,
   I1 => x71_out_20,
   I2 => x71_out_22,
   I3 => W_41_7_i_16_n_0,
   I4 => W_41_7_i_17_n_0,
   O => W_41_7_i_5_n_0
);
W_41_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_41_7_i_2_n_0,
   I1 => W_41_11_i_16_n_0,
   I2 => x71_out_17,
   I3 => x71_out_24,
   I4 => x71_out_26,
   I5 => W_41_11_i_17_n_0,
   O => W_41_7_i_6_n_0
);
W_41_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_41_7_i_3_n_0,
   I1 => W_41_7_i_10_n_0,
   I2 => x71_out_16,
   I3 => x71_out_23,
   I4 => x71_out_25,
   I5 => W_41_7_i_11_n_0,
   O => W_41_7_i_7_n_0
);
W_41_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_41_7_i_4_n_0,
   I1 => W_41_7_i_12_n_0,
   I2 => x71_out_15,
   I3 => x71_out_22,
   I4 => x71_out_24,
   I5 => W_41_7_i_13_n_0,
   O => W_41_7_i_8_n_0
);
W_41_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_41_7_i_5_n_0,
   I1 => W_41_7_i_14_n_0,
   I2 => x71_out_14,
   I3 => x71_out_21,
   I4 => x71_out_23,
   I5 => W_41_7_i_15_n_0,
   O => W_41_7_i_9_n_0
);
W_42_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x104_out_10,
   I1 => x83_out_10,
   I2 => x102_out_28,
   I3 => x102_out_17,
   I4 => x102_out_13,
   O => W_42_11_i_10_n_0
);
W_42_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x83_out_9,
   I1 => x102_out_12,
   I2 => x102_out_16,
   I3 => x102_out_27,
   I4 => x104_out_9,
   O => W_42_11_i_11_n_0
);
W_42_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x104_out_9,
   I1 => x83_out_9,
   I2 => x102_out_27,
   I3 => x102_out_16,
   I4 => x102_out_12,
   O => W_42_11_i_12_n_0
);
W_42_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x83_out_8,
   I1 => x102_out_11,
   I2 => x102_out_15,
   I3 => x102_out_26,
   I4 => x104_out_8,
   O => W_42_11_i_13_n_0
);
W_42_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x104_out_8,
   I1 => x83_out_8,
   I2 => x102_out_26,
   I3 => x102_out_15,
   I4 => x102_out_11,
   O => W_42_11_i_14_n_0
);
W_42_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x83_out_7,
   I1 => x102_out_10,
   I2 => x102_out_14,
   I3 => x102_out_25,
   I4 => x104_out_7,
   O => W_42_11_i_15_n_0
);
W_42_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x104_out_7,
   I1 => x83_out_7,
   I2 => x102_out_25,
   I3 => x102_out_14,
   I4 => x102_out_10,
   O => W_42_11_i_16_n_0
);
W_42_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x83_out_6,
   I1 => x102_out_9,
   I2 => x102_out_13,
   I3 => x102_out_24,
   I4 => x104_out_6,
   O => W_42_11_i_17_n_0
);
W_42_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x68_out_20,
   I1 => x68_out_27,
   I2 => x68_out_29,
   I3 => W_42_11_i_10_n_0,
   I4 => W_42_11_i_11_n_0,
   O => W_42_11_i_2_n_0
);
W_42_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x68_out_19,
   I1 => x68_out_26,
   I2 => x68_out_28,
   I3 => W_42_11_i_12_n_0,
   I4 => W_42_11_i_13_n_0,
   O => W_42_11_i_3_n_0
);
W_42_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x68_out_18,
   I1 => x68_out_25,
   I2 => x68_out_27,
   I3 => W_42_11_i_14_n_0,
   I4 => W_42_11_i_15_n_0,
   O => W_42_11_i_4_n_0
);
W_42_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x68_out_17,
   I1 => x68_out_24,
   I2 => x68_out_26,
   I3 => W_42_11_i_16_n_0,
   I4 => W_42_11_i_17_n_0,
   O => W_42_11_i_5_n_0
);
W_42_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_42_11_i_2_n_0,
   I1 => W_42_15_i_16_n_0,
   I2 => x68_out_21,
   I3 => x68_out_28,
   I4 => x68_out_30,
   I5 => W_42_15_i_17_n_0,
   O => W_42_11_i_6_n_0
);
W_42_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_42_11_i_3_n_0,
   I1 => W_42_11_i_10_n_0,
   I2 => x68_out_20,
   I3 => x68_out_27,
   I4 => x68_out_29,
   I5 => W_42_11_i_11_n_0,
   O => W_42_11_i_7_n_0
);
W_42_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_42_11_i_4_n_0,
   I1 => W_42_11_i_12_n_0,
   I2 => x68_out_19,
   I3 => x68_out_26,
   I4 => x68_out_28,
   I5 => W_42_11_i_13_n_0,
   O => W_42_11_i_8_n_0
);
W_42_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_42_11_i_5_n_0,
   I1 => W_42_11_i_14_n_0,
   I2 => x68_out_18,
   I3 => x68_out_25,
   I4 => x68_out_27,
   I5 => W_42_11_i_15_n_0,
   O => W_42_11_i_9_n_0
);
W_42_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x104_out_14,
   I1 => x83_out_14,
   I2 => x102_out_0,
   I3 => x102_out_21,
   I4 => x102_out_17,
   O => W_42_15_i_10_n_0
);
W_42_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x83_out_13,
   I1 => x102_out_16,
   I2 => x102_out_20,
   I3 => x102_out_31,
   I4 => x104_out_13,
   O => W_42_15_i_11_n_0
);
W_42_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x104_out_13,
   I1 => x83_out_13,
   I2 => x102_out_31,
   I3 => x102_out_20,
   I4 => x102_out_16,
   O => W_42_15_i_12_n_0
);
W_42_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x83_out_12,
   I1 => x102_out_15,
   I2 => x102_out_19,
   I3 => x102_out_30,
   I4 => x104_out_12,
   O => W_42_15_i_13_n_0
);
W_42_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x104_out_12,
   I1 => x83_out_12,
   I2 => x102_out_30,
   I3 => x102_out_19,
   I4 => x102_out_15,
   O => W_42_15_i_14_n_0
);
W_42_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x83_out_11,
   I1 => x102_out_14,
   I2 => x102_out_18,
   I3 => x102_out_29,
   I4 => x104_out_11,
   O => W_42_15_i_15_n_0
);
W_42_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x104_out_11,
   I1 => x83_out_11,
   I2 => x102_out_29,
   I3 => x102_out_18,
   I4 => x102_out_14,
   O => W_42_15_i_16_n_0
);
W_42_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x83_out_10,
   I1 => x102_out_13,
   I2 => x102_out_17,
   I3 => x102_out_28,
   I4 => x104_out_10,
   O => W_42_15_i_17_n_0
);
W_42_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x68_out_24,
   I1 => x68_out_31,
   I2 => x68_out_1,
   I3 => W_42_15_i_10_n_0,
   I4 => W_42_15_i_11_n_0,
   O => W_42_15_i_2_n_0
);
W_42_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x68_out_23,
   I1 => x68_out_30,
   I2 => x68_out_0,
   I3 => W_42_15_i_12_n_0,
   I4 => W_42_15_i_13_n_0,
   O => W_42_15_i_3_n_0
);
W_42_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x68_out_22,
   I1 => x68_out_29,
   I2 => x68_out_31,
   I3 => W_42_15_i_14_n_0,
   I4 => W_42_15_i_15_n_0,
   O => W_42_15_i_4_n_0
);
W_42_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x68_out_21,
   I1 => x68_out_28,
   I2 => x68_out_30,
   I3 => W_42_15_i_16_n_0,
   I4 => W_42_15_i_17_n_0,
   O => W_42_15_i_5_n_0
);
W_42_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_42_15_i_2_n_0,
   I1 => W_42_19_i_16_n_0,
   I2 => x68_out_25,
   I3 => x68_out_0,
   I4 => x68_out_2,
   I5 => W_42_19_i_17_n_0,
   O => W_42_15_i_6_n_0
);
W_42_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_42_15_i_3_n_0,
   I1 => W_42_15_i_10_n_0,
   I2 => x68_out_24,
   I3 => x68_out_31,
   I4 => x68_out_1,
   I5 => W_42_15_i_11_n_0,
   O => W_42_15_i_7_n_0
);
W_42_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_42_15_i_4_n_0,
   I1 => W_42_15_i_12_n_0,
   I2 => x68_out_23,
   I3 => x68_out_30,
   I4 => x68_out_0,
   I5 => W_42_15_i_13_n_0,
   O => W_42_15_i_8_n_0
);
W_42_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_42_15_i_5_n_0,
   I1 => W_42_15_i_14_n_0,
   I2 => x68_out_22,
   I3 => x68_out_29,
   I4 => x68_out_31,
   I5 => W_42_15_i_15_n_0,
   O => W_42_15_i_9_n_0
);
W_42_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x104_out_18,
   I1 => x83_out_18,
   I2 => x102_out_4,
   I3 => x102_out_25,
   I4 => x102_out_21,
   O => W_42_19_i_10_n_0
);
W_42_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x83_out_17,
   I1 => x102_out_20,
   I2 => x102_out_24,
   I3 => x102_out_3,
   I4 => x104_out_17,
   O => W_42_19_i_11_n_0
);
W_42_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x104_out_17,
   I1 => x83_out_17,
   I2 => x102_out_3,
   I3 => x102_out_24,
   I4 => x102_out_20,
   O => W_42_19_i_12_n_0
);
W_42_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x83_out_16,
   I1 => x102_out_19,
   I2 => x102_out_23,
   I3 => x102_out_2,
   I4 => x104_out_16,
   O => W_42_19_i_13_n_0
);
W_42_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x104_out_16,
   I1 => x83_out_16,
   I2 => x102_out_2,
   I3 => x102_out_23,
   I4 => x102_out_19,
   O => W_42_19_i_14_n_0
);
W_42_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x83_out_15,
   I1 => x102_out_18,
   I2 => x102_out_22,
   I3 => x102_out_1,
   I4 => x104_out_15,
   O => W_42_19_i_15_n_0
);
W_42_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x104_out_15,
   I1 => x83_out_15,
   I2 => x102_out_1,
   I3 => x102_out_22,
   I4 => x102_out_18,
   O => W_42_19_i_16_n_0
);
W_42_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x83_out_14,
   I1 => x102_out_17,
   I2 => x102_out_21,
   I3 => x102_out_0,
   I4 => x104_out_14,
   O => W_42_19_i_17_n_0
);
W_42_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x68_out_28,
   I1 => x68_out_3,
   I2 => x68_out_5,
   I3 => W_42_19_i_10_n_0,
   I4 => W_42_19_i_11_n_0,
   O => W_42_19_i_2_n_0
);
W_42_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x68_out_27,
   I1 => x68_out_2,
   I2 => x68_out_4,
   I3 => W_42_19_i_12_n_0,
   I4 => W_42_19_i_13_n_0,
   O => W_42_19_i_3_n_0
);
W_42_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x68_out_26,
   I1 => x68_out_1,
   I2 => x68_out_3,
   I3 => W_42_19_i_14_n_0,
   I4 => W_42_19_i_15_n_0,
   O => W_42_19_i_4_n_0
);
W_42_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x68_out_25,
   I1 => x68_out_0,
   I2 => x68_out_2,
   I3 => W_42_19_i_16_n_0,
   I4 => W_42_19_i_17_n_0,
   O => W_42_19_i_5_n_0
);
W_42_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_42_19_i_2_n_0,
   I1 => W_42_23_i_16_n_0,
   I2 => x68_out_29,
   I3 => x68_out_4,
   I4 => x68_out_6,
   I5 => W_42_23_i_17_n_0,
   O => W_42_19_i_6_n_0
);
W_42_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_42_19_i_3_n_0,
   I1 => W_42_19_i_10_n_0,
   I2 => x68_out_28,
   I3 => x68_out_3,
   I4 => x68_out_5,
   I5 => W_42_19_i_11_n_0,
   O => W_42_19_i_7_n_0
);
W_42_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_42_19_i_4_n_0,
   I1 => W_42_19_i_12_n_0,
   I2 => x68_out_27,
   I3 => x68_out_2,
   I4 => x68_out_4,
   I5 => W_42_19_i_13_n_0,
   O => W_42_19_i_8_n_0
);
W_42_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_42_19_i_5_n_0,
   I1 => W_42_19_i_14_n_0,
   I2 => x68_out_26,
   I3 => x68_out_1,
   I4 => x68_out_3,
   I5 => W_42_19_i_15_n_0,
   O => W_42_19_i_9_n_0
);
W_42_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x104_out_22,
   I1 => x83_out_22,
   I2 => x102_out_8,
   I3 => x102_out_29,
   I4 => x102_out_25,
   O => W_42_23_i_10_n_0
);
W_42_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x83_out_21,
   I1 => x102_out_24,
   I2 => x102_out_28,
   I3 => x102_out_7,
   I4 => x104_out_21,
   O => W_42_23_i_11_n_0
);
W_42_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x104_out_21,
   I1 => x83_out_21,
   I2 => x102_out_7,
   I3 => x102_out_28,
   I4 => x102_out_24,
   O => W_42_23_i_12_n_0
);
W_42_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x83_out_20,
   I1 => x102_out_23,
   I2 => x102_out_27,
   I3 => x102_out_6,
   I4 => x104_out_20,
   O => W_42_23_i_13_n_0
);
W_42_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x104_out_20,
   I1 => x83_out_20,
   I2 => x102_out_6,
   I3 => x102_out_27,
   I4 => x102_out_23,
   O => W_42_23_i_14_n_0
);
W_42_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x83_out_19,
   I1 => x102_out_22,
   I2 => x102_out_26,
   I3 => x102_out_5,
   I4 => x104_out_19,
   O => W_42_23_i_15_n_0
);
W_42_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x104_out_19,
   I1 => x83_out_19,
   I2 => x102_out_5,
   I3 => x102_out_26,
   I4 => x102_out_22,
   O => W_42_23_i_16_n_0
);
W_42_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x83_out_18,
   I1 => x102_out_21,
   I2 => x102_out_25,
   I3 => x102_out_4,
   I4 => x104_out_18,
   O => W_42_23_i_17_n_0
);
W_42_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x68_out_7,
   I1 => x68_out_9,
   I2 => W_42_23_i_10_n_0,
   I3 => W_42_23_i_11_n_0,
   O => W_42_23_i_2_n_0
);
W_42_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x68_out_31,
   I1 => x68_out_6,
   I2 => x68_out_8,
   I3 => W_42_23_i_12_n_0,
   I4 => W_42_23_i_13_n_0,
   O => W_42_23_i_3_n_0
);
W_42_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x68_out_30,
   I1 => x68_out_5,
   I2 => x68_out_7,
   I3 => W_42_23_i_14_n_0,
   I4 => W_42_23_i_15_n_0,
   O => W_42_23_i_4_n_0
);
W_42_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x68_out_29,
   I1 => x68_out_4,
   I2 => x68_out_6,
   I3 => W_42_23_i_16_n_0,
   I4 => W_42_23_i_17_n_0,
   O => W_42_23_i_5_n_0
);
W_42_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x68_out_8,
   I1 => x68_out_10,
   I2 => W_42_27_i_16_n_0,
   I3 => W_42_27_i_17_n_0,
   I4 => W_42_23_i_2_n_0,
   O => W_42_23_i_6_n_0
);
W_42_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x68_out_7,
   I1 => x68_out_9,
   I2 => W_42_23_i_10_n_0,
   I3 => W_42_23_i_11_n_0,
   I4 => W_42_23_i_3_n_0,
   O => W_42_23_i_7_n_0
);
W_42_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_42_23_i_4_n_0,
   I1 => W_42_23_i_12_n_0,
   I2 => x68_out_31,
   I3 => x68_out_6,
   I4 => x68_out_8,
   I5 => W_42_23_i_13_n_0,
   O => W_42_23_i_8_n_0
);
W_42_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_42_23_i_5_n_0,
   I1 => W_42_23_i_14_n_0,
   I2 => x68_out_30,
   I3 => x68_out_5,
   I4 => x68_out_7,
   I5 => W_42_23_i_15_n_0,
   O => W_42_23_i_9_n_0
);
W_42_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x104_out_26,
   I1 => x83_out_26,
   I2 => x102_out_12,
   I3 => x102_out_1,
   I4 => x102_out_29,
   O => W_42_27_i_10_n_0
);
W_42_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x83_out_25,
   I1 => x102_out_28,
   I2 => x102_out_0,
   I3 => x102_out_11,
   I4 => x104_out_25,
   O => W_42_27_i_11_n_0
);
W_42_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x104_out_25,
   I1 => x83_out_25,
   I2 => x102_out_11,
   I3 => x102_out_0,
   I4 => x102_out_28,
   O => W_42_27_i_12_n_0
);
W_42_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x83_out_24,
   I1 => x102_out_27,
   I2 => x102_out_31,
   I3 => x102_out_10,
   I4 => x104_out_24,
   O => W_42_27_i_13_n_0
);
W_42_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x104_out_24,
   I1 => x83_out_24,
   I2 => x102_out_10,
   I3 => x102_out_31,
   I4 => x102_out_27,
   O => W_42_27_i_14_n_0
);
W_42_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x83_out_23,
   I1 => x102_out_26,
   I2 => x102_out_30,
   I3 => x102_out_9,
   I4 => x104_out_23,
   O => W_42_27_i_15_n_0
);
W_42_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x104_out_23,
   I1 => x83_out_23,
   I2 => x102_out_9,
   I3 => x102_out_30,
   I4 => x102_out_26,
   O => W_42_27_i_16_n_0
);
W_42_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x83_out_22,
   I1 => x102_out_25,
   I2 => x102_out_29,
   I3 => x102_out_8,
   I4 => x104_out_22,
   O => W_42_27_i_17_n_0
);
W_42_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x68_out_11,
   I1 => x68_out_13,
   I2 => W_42_27_i_10_n_0,
   I3 => W_42_27_i_11_n_0,
   O => W_42_27_i_2_n_0
);
W_42_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x68_out_10,
   I1 => x68_out_12,
   I2 => W_42_27_i_12_n_0,
   I3 => W_42_27_i_13_n_0,
   O => W_42_27_i_3_n_0
);
W_42_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x68_out_9,
   I1 => x68_out_11,
   I2 => W_42_27_i_14_n_0,
   I3 => W_42_27_i_15_n_0,
   O => W_42_27_i_4_n_0
);
W_42_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x68_out_8,
   I1 => x68_out_10,
   I2 => W_42_27_i_16_n_0,
   I3 => W_42_27_i_17_n_0,
   O => W_42_27_i_5_n_0
);
W_42_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x68_out_12,
   I1 => x68_out_14,
   I2 => W_42_31_i_13_n_0,
   I3 => W_42_31_i_14_n_0,
   I4 => W_42_27_i_2_n_0,
   O => W_42_27_i_6_n_0
);
W_42_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x68_out_11,
   I1 => x68_out_13,
   I2 => W_42_27_i_10_n_0,
   I3 => W_42_27_i_11_n_0,
   I4 => W_42_27_i_3_n_0,
   O => W_42_27_i_7_n_0
);
W_42_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x68_out_10,
   I1 => x68_out_12,
   I2 => W_42_27_i_12_n_0,
   I3 => W_42_27_i_13_n_0,
   I4 => W_42_27_i_4_n_0,
   O => W_42_27_i_8_n_0
);
W_42_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x68_out_9,
   I1 => x68_out_11,
   I2 => W_42_27_i_14_n_0,
   I3 => W_42_27_i_15_n_0,
   I4 => W_42_27_i_5_n_0,
   O => W_42_27_i_9_n_0
);
W_42_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x83_out_28,
   I1 => x102_out_31,
   I2 => x102_out_3,
   I3 => x102_out_14,
   I4 => x104_out_28,
   O => W_42_31_i_10_n_0
);
W_42_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x104_out_28,
   I1 => x83_out_28,
   I2 => x102_out_14,
   I3 => x102_out_3,
   I4 => x102_out_31,
   O => W_42_31_i_11_n_0
);
W_42_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x83_out_27,
   I1 => x102_out_30,
   I2 => x102_out_2,
   I3 => x102_out_13,
   I4 => x104_out_27,
   O => W_42_31_i_12_n_0
);
W_42_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x104_out_27,
   I1 => x83_out_27,
   I2 => x102_out_13,
   I3 => x102_out_2,
   I4 => x102_out_30,
   O => W_42_31_i_13_n_0
);
W_42_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x83_out_26,
   I1 => x102_out_29,
   I2 => x102_out_1,
   I3 => x102_out_12,
   I4 => x104_out_26,
   O => W_42_31_i_14_n_0
);
W_42_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x83_out_29,
   I1 => x102_out_4,
   I2 => x102_out_15,
   I3 => x104_out_29,
   O => W_42_31_i_15_n_0
);
W_42_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x68_out_17,
   I1 => x68_out_15,
   O => SIGMA_LCASE_1179_out_0_30
);
W_42_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => x102_out_6,
   I1 => x102_out_17,
   I2 => x83_out_31,
   I3 => x104_out_31,
   I4 => x68_out_16,
   I5 => x68_out_18,
   O => W_42_31_i_17_n_0
);
W_42_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x102_out_16,
   I1 => x102_out_5,
   O => SIGMA_LCASE_0175_out_30
);
W_42_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x104_out_30,
   I1 => x83_out_30,
   I2 => x102_out_16,
   I3 => x102_out_5,
   O => W_42_31_i_19_n_0
);
W_42_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x68_out_14,
   I1 => x68_out_16,
   I2 => W_42_31_i_9_n_0,
   I3 => W_42_31_i_10_n_0,
   O => W_42_31_i_2_n_0
);
W_42_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x68_out_13,
   I1 => x68_out_15,
   I2 => W_42_31_i_11_n_0,
   I3 => W_42_31_i_12_n_0,
   O => W_42_31_i_3_n_0
);
W_42_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x68_out_12,
   I1 => x68_out_14,
   I2 => W_42_31_i_13_n_0,
   I3 => W_42_31_i_14_n_0,
   O => W_42_31_i_4_n_0
);
W_42_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_42_31_i_15_n_0,
   I1 => SIGMA_LCASE_1179_out_0_30,
   I2 => W_42_31_i_17_n_0,
   I3 => x83_out_30,
   I4 => SIGMA_LCASE_0175_out_30,
   I5 => x104_out_30,
   O => W_42_31_i_5_n_0
);
W_42_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_42_31_i_2_n_0,
   I1 => W_42_31_i_19_n_0,
   I2 => x68_out_15,
   I3 => x68_out_17,
   I4 => W_42_31_i_15_n_0,
   O => W_42_31_i_6_n_0
);
W_42_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x68_out_14,
   I1 => x68_out_16,
   I2 => W_42_31_i_9_n_0,
   I3 => W_42_31_i_10_n_0,
   I4 => W_42_31_i_3_n_0,
   O => W_42_31_i_7_n_0
);
W_42_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x68_out_13,
   I1 => x68_out_15,
   I2 => W_42_31_i_11_n_0,
   I3 => W_42_31_i_12_n_0,
   I4 => W_42_31_i_4_n_0,
   O => W_42_31_i_8_n_0
);
W_42_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x104_out_29,
   I1 => x83_out_29,
   I2 => x102_out_15,
   I3 => x102_out_4,
   O => W_42_31_i_9_n_0
);
W_42_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x104_out_2,
   I1 => x83_out_2,
   I2 => x102_out_20,
   I3 => x102_out_9,
   I4 => x102_out_5,
   O => W_42_3_i_10_n_0
);
W_42_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x83_out_1,
   I1 => x102_out_4,
   I2 => x102_out_8,
   I3 => x102_out_19,
   I4 => x104_out_1,
   O => W_42_3_i_11_n_0
);
W_42_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x102_out_19,
   I1 => x102_out_8,
   I2 => x102_out_4,
   O => SIGMA_LCASE_0175_out_1
);
W_42_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x68_out_21,
   I1 => x68_out_19,
   I2 => x68_out_12,
   O => SIGMA_LCASE_1179_out_0_2
);
W_42_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x68_out_20,
   I1 => x68_out_18,
   I2 => x68_out_11,
   O => SIGMA_LCASE_1179_out_1
);
W_42_3_i_15 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x104_out_1,
   I1 => x83_out_1,
   I2 => x102_out_19,
   I3 => x102_out_8,
   I4 => x102_out_4,
   O => W_42_3_i_15_n_0
);
W_42_3_i_16 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x102_out_18,
   I1 => x102_out_7,
   I2 => x102_out_3,
   O => SIGMA_LCASE_0175_out_0
);
W_42_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x68_out_12,
   I1 => x68_out_19,
   I2 => x68_out_21,
   I3 => W_42_3_i_10_n_0,
   I4 => W_42_3_i_11_n_0,
   O => W_42_3_i_2_n_0
);
W_42_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_42_3_i_11_n_0,
   I1 => x68_out_21,
   I2 => x68_out_19,
   I3 => x68_out_12,
   I4 => W_42_3_i_10_n_0,
   O => W_42_3_i_3_n_0
);
W_42_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_0175_out_1,
   I1 => x83_out_1,
   I2 => x104_out_1,
   I3 => x68_out_11,
   I4 => x68_out_18,
   I5 => x68_out_20,
   O => W_42_3_i_4_n_0
);
W_42_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x104_out_0,
   I1 => x83_out_0,
   I2 => x102_out_18,
   I3 => x102_out_7,
   I4 => x102_out_3,
   O => W_42_3_i_5_n_0
);
W_42_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_42_3_i_2_n_0,
   I1 => W_42_7_i_16_n_0,
   I2 => x68_out_13,
   I3 => x68_out_20,
   I4 => x68_out_22,
   I5 => W_42_7_i_17_n_0,
   O => W_42_3_i_6_n_0
);
W_42_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_42_3_i_10_n_0,
   I1 => SIGMA_LCASE_1179_out_0_2,
   I2 => x104_out_1,
   I3 => x83_out_1,
   I4 => SIGMA_LCASE_0175_out_1,
   I5 => SIGMA_LCASE_1179_out_1,
   O => W_42_3_i_7_n_0
);
W_42_3_i_8 : LUT5
  generic map(
   INIT => X"99969666"
  )
 port map (
   I0 => SIGMA_LCASE_1179_out_1,
   I1 => W_42_3_i_15_n_0,
   I2 => x104_out_0,
   I3 => SIGMA_LCASE_0175_out_0,
   I4 => x83_out_0,
   O => W_42_3_i_8_n_0
);
W_42_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_42_3_i_5_n_0,
   I1 => x68_out_10,
   I2 => x68_out_17,
   I3 => x68_out_19,
   O => W_42_3_i_9_n_0
);
W_42_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x104_out_6,
   I1 => x83_out_6,
   I2 => x102_out_24,
   I3 => x102_out_13,
   I4 => x102_out_9,
   O => W_42_7_i_10_n_0
);
W_42_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x83_out_5,
   I1 => x102_out_8,
   I2 => x102_out_12,
   I3 => x102_out_23,
   I4 => x104_out_5,
   O => W_42_7_i_11_n_0
);
W_42_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x104_out_5,
   I1 => x83_out_5,
   I2 => x102_out_23,
   I3 => x102_out_12,
   I4 => x102_out_8,
   O => W_42_7_i_12_n_0
);
W_42_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x83_out_4,
   I1 => x102_out_7,
   I2 => x102_out_11,
   I3 => x102_out_22,
   I4 => x104_out_4,
   O => W_42_7_i_13_n_0
);
W_42_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x104_out_4,
   I1 => x83_out_4,
   I2 => x102_out_22,
   I3 => x102_out_11,
   I4 => x102_out_7,
   O => W_42_7_i_14_n_0
);
W_42_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x83_out_3,
   I1 => x102_out_6,
   I2 => x102_out_10,
   I3 => x102_out_21,
   I4 => x104_out_3,
   O => W_42_7_i_15_n_0
);
W_42_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x104_out_3,
   I1 => x83_out_3,
   I2 => x102_out_21,
   I3 => x102_out_10,
   I4 => x102_out_6,
   O => W_42_7_i_16_n_0
);
W_42_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x83_out_2,
   I1 => x102_out_5,
   I2 => x102_out_9,
   I3 => x102_out_20,
   I4 => x104_out_2,
   O => W_42_7_i_17_n_0
);
W_42_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x68_out_16,
   I1 => x68_out_23,
   I2 => x68_out_25,
   I3 => W_42_7_i_10_n_0,
   I4 => W_42_7_i_11_n_0,
   O => W_42_7_i_2_n_0
);
W_42_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x68_out_15,
   I1 => x68_out_22,
   I2 => x68_out_24,
   I3 => W_42_7_i_12_n_0,
   I4 => W_42_7_i_13_n_0,
   O => W_42_7_i_3_n_0
);
W_42_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x68_out_14,
   I1 => x68_out_21,
   I2 => x68_out_23,
   I3 => W_42_7_i_14_n_0,
   I4 => W_42_7_i_15_n_0,
   O => W_42_7_i_4_n_0
);
W_42_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x68_out_13,
   I1 => x68_out_20,
   I2 => x68_out_22,
   I3 => W_42_7_i_16_n_0,
   I4 => W_42_7_i_17_n_0,
   O => W_42_7_i_5_n_0
);
W_42_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_42_7_i_2_n_0,
   I1 => W_42_11_i_16_n_0,
   I2 => x68_out_17,
   I3 => x68_out_24,
   I4 => x68_out_26,
   I5 => W_42_11_i_17_n_0,
   O => W_42_7_i_6_n_0
);
W_42_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_42_7_i_3_n_0,
   I1 => W_42_7_i_10_n_0,
   I2 => x68_out_16,
   I3 => x68_out_23,
   I4 => x68_out_25,
   I5 => W_42_7_i_11_n_0,
   O => W_42_7_i_7_n_0
);
W_42_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_42_7_i_4_n_0,
   I1 => W_42_7_i_12_n_0,
   I2 => x68_out_15,
   I3 => x68_out_22,
   I4 => x68_out_24,
   I5 => W_42_7_i_13_n_0,
   O => W_42_7_i_8_n_0
);
W_42_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_42_7_i_5_n_0,
   I1 => W_42_7_i_14_n_0,
   I2 => x68_out_14,
   I3 => x68_out_21,
   I4 => x68_out_23,
   I5 => W_42_7_i_15_n_0,
   O => W_42_7_i_9_n_0
);
W_43_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x102_out_10,
   I1 => x80_out_10,
   I2 => x100_out_28,
   I3 => x100_out_17,
   I4 => x100_out_13,
   O => W_43_11_i_10_n_0
);
W_43_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x80_out_9,
   I1 => x100_out_12,
   I2 => x100_out_16,
   I3 => x100_out_27,
   I4 => x102_out_9,
   O => W_43_11_i_11_n_0
);
W_43_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x102_out_9,
   I1 => x80_out_9,
   I2 => x100_out_27,
   I3 => x100_out_16,
   I4 => x100_out_12,
   O => W_43_11_i_12_n_0
);
W_43_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x80_out_8,
   I1 => x100_out_11,
   I2 => x100_out_15,
   I3 => x100_out_26,
   I4 => x102_out_8,
   O => W_43_11_i_13_n_0
);
W_43_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x102_out_8,
   I1 => x80_out_8,
   I2 => x100_out_26,
   I3 => x100_out_15,
   I4 => x100_out_11,
   O => W_43_11_i_14_n_0
);
W_43_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x80_out_7,
   I1 => x100_out_10,
   I2 => x100_out_14,
   I3 => x100_out_25,
   I4 => x102_out_7,
   O => W_43_11_i_15_n_0
);
W_43_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x102_out_7,
   I1 => x80_out_7,
   I2 => x100_out_25,
   I3 => x100_out_14,
   I4 => x100_out_10,
   O => W_43_11_i_16_n_0
);
W_43_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x80_out_6,
   I1 => x100_out_9,
   I2 => x100_out_13,
   I3 => x100_out_24,
   I4 => x102_out_6,
   O => W_43_11_i_17_n_0
);
W_43_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x65_out_20,
   I1 => x65_out_27,
   I2 => x65_out_29,
   I3 => W_43_11_i_10_n_0,
   I4 => W_43_11_i_11_n_0,
   O => W_43_11_i_2_n_0
);
W_43_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x65_out_19,
   I1 => x65_out_26,
   I2 => x65_out_28,
   I3 => W_43_11_i_12_n_0,
   I4 => W_43_11_i_13_n_0,
   O => W_43_11_i_3_n_0
);
W_43_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x65_out_18,
   I1 => x65_out_25,
   I2 => x65_out_27,
   I3 => W_43_11_i_14_n_0,
   I4 => W_43_11_i_15_n_0,
   O => W_43_11_i_4_n_0
);
W_43_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x65_out_17,
   I1 => x65_out_24,
   I2 => x65_out_26,
   I3 => W_43_11_i_16_n_0,
   I4 => W_43_11_i_17_n_0,
   O => W_43_11_i_5_n_0
);
W_43_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_43_11_i_2_n_0,
   I1 => W_43_15_i_16_n_0,
   I2 => x65_out_21,
   I3 => x65_out_28,
   I4 => x65_out_30,
   I5 => W_43_15_i_17_n_0,
   O => W_43_11_i_6_n_0
);
W_43_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_43_11_i_3_n_0,
   I1 => W_43_11_i_10_n_0,
   I2 => x65_out_20,
   I3 => x65_out_27,
   I4 => x65_out_29,
   I5 => W_43_11_i_11_n_0,
   O => W_43_11_i_7_n_0
);
W_43_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_43_11_i_4_n_0,
   I1 => W_43_11_i_12_n_0,
   I2 => x65_out_19,
   I3 => x65_out_26,
   I4 => x65_out_28,
   I5 => W_43_11_i_13_n_0,
   O => W_43_11_i_8_n_0
);
W_43_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_43_11_i_5_n_0,
   I1 => W_43_11_i_14_n_0,
   I2 => x65_out_18,
   I3 => x65_out_25,
   I4 => x65_out_27,
   I5 => W_43_11_i_15_n_0,
   O => W_43_11_i_9_n_0
);
W_43_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x102_out_14,
   I1 => x80_out_14,
   I2 => x100_out_0,
   I3 => x100_out_21,
   I4 => x100_out_17,
   O => W_43_15_i_10_n_0
);
W_43_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x80_out_13,
   I1 => x100_out_16,
   I2 => x100_out_20,
   I3 => x100_out_31,
   I4 => x102_out_13,
   O => W_43_15_i_11_n_0
);
W_43_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x102_out_13,
   I1 => x80_out_13,
   I2 => x100_out_31,
   I3 => x100_out_20,
   I4 => x100_out_16,
   O => W_43_15_i_12_n_0
);
W_43_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x80_out_12,
   I1 => x100_out_15,
   I2 => x100_out_19,
   I3 => x100_out_30,
   I4 => x102_out_12,
   O => W_43_15_i_13_n_0
);
W_43_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x102_out_12,
   I1 => x80_out_12,
   I2 => x100_out_30,
   I3 => x100_out_19,
   I4 => x100_out_15,
   O => W_43_15_i_14_n_0
);
W_43_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x80_out_11,
   I1 => x100_out_14,
   I2 => x100_out_18,
   I3 => x100_out_29,
   I4 => x102_out_11,
   O => W_43_15_i_15_n_0
);
W_43_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x102_out_11,
   I1 => x80_out_11,
   I2 => x100_out_29,
   I3 => x100_out_18,
   I4 => x100_out_14,
   O => W_43_15_i_16_n_0
);
W_43_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x80_out_10,
   I1 => x100_out_13,
   I2 => x100_out_17,
   I3 => x100_out_28,
   I4 => x102_out_10,
   O => W_43_15_i_17_n_0
);
W_43_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x65_out_24,
   I1 => x65_out_31,
   I2 => x65_out_1,
   I3 => W_43_15_i_10_n_0,
   I4 => W_43_15_i_11_n_0,
   O => W_43_15_i_2_n_0
);
W_43_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x65_out_23,
   I1 => x65_out_30,
   I2 => x65_out_0,
   I3 => W_43_15_i_12_n_0,
   I4 => W_43_15_i_13_n_0,
   O => W_43_15_i_3_n_0
);
W_43_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x65_out_22,
   I1 => x65_out_29,
   I2 => x65_out_31,
   I3 => W_43_15_i_14_n_0,
   I4 => W_43_15_i_15_n_0,
   O => W_43_15_i_4_n_0
);
W_43_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x65_out_21,
   I1 => x65_out_28,
   I2 => x65_out_30,
   I3 => W_43_15_i_16_n_0,
   I4 => W_43_15_i_17_n_0,
   O => W_43_15_i_5_n_0
);
W_43_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_43_15_i_2_n_0,
   I1 => W_43_19_i_16_n_0,
   I2 => x65_out_25,
   I3 => x65_out_0,
   I4 => x65_out_2,
   I5 => W_43_19_i_17_n_0,
   O => W_43_15_i_6_n_0
);
W_43_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_43_15_i_3_n_0,
   I1 => W_43_15_i_10_n_0,
   I2 => x65_out_24,
   I3 => x65_out_31,
   I4 => x65_out_1,
   I5 => W_43_15_i_11_n_0,
   O => W_43_15_i_7_n_0
);
W_43_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_43_15_i_4_n_0,
   I1 => W_43_15_i_12_n_0,
   I2 => x65_out_23,
   I3 => x65_out_30,
   I4 => x65_out_0,
   I5 => W_43_15_i_13_n_0,
   O => W_43_15_i_8_n_0
);
W_43_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_43_15_i_5_n_0,
   I1 => W_43_15_i_14_n_0,
   I2 => x65_out_22,
   I3 => x65_out_29,
   I4 => x65_out_31,
   I5 => W_43_15_i_15_n_0,
   O => W_43_15_i_9_n_0
);
W_43_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x102_out_18,
   I1 => x80_out_18,
   I2 => x100_out_4,
   I3 => x100_out_25,
   I4 => x100_out_21,
   O => W_43_19_i_10_n_0
);
W_43_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x80_out_17,
   I1 => x100_out_20,
   I2 => x100_out_24,
   I3 => x100_out_3,
   I4 => x102_out_17,
   O => W_43_19_i_11_n_0
);
W_43_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x102_out_17,
   I1 => x80_out_17,
   I2 => x100_out_3,
   I3 => x100_out_24,
   I4 => x100_out_20,
   O => W_43_19_i_12_n_0
);
W_43_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x80_out_16,
   I1 => x100_out_19,
   I2 => x100_out_23,
   I3 => x100_out_2,
   I4 => x102_out_16,
   O => W_43_19_i_13_n_0
);
W_43_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x102_out_16,
   I1 => x80_out_16,
   I2 => x100_out_2,
   I3 => x100_out_23,
   I4 => x100_out_19,
   O => W_43_19_i_14_n_0
);
W_43_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x80_out_15,
   I1 => x100_out_18,
   I2 => x100_out_22,
   I3 => x100_out_1,
   I4 => x102_out_15,
   O => W_43_19_i_15_n_0
);
W_43_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x102_out_15,
   I1 => x80_out_15,
   I2 => x100_out_1,
   I3 => x100_out_22,
   I4 => x100_out_18,
   O => W_43_19_i_16_n_0
);
W_43_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x80_out_14,
   I1 => x100_out_17,
   I2 => x100_out_21,
   I3 => x100_out_0,
   I4 => x102_out_14,
   O => W_43_19_i_17_n_0
);
W_43_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x65_out_28,
   I1 => x65_out_3,
   I2 => x65_out_5,
   I3 => W_43_19_i_10_n_0,
   I4 => W_43_19_i_11_n_0,
   O => W_43_19_i_2_n_0
);
W_43_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x65_out_27,
   I1 => x65_out_2,
   I2 => x65_out_4,
   I3 => W_43_19_i_12_n_0,
   I4 => W_43_19_i_13_n_0,
   O => W_43_19_i_3_n_0
);
W_43_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x65_out_26,
   I1 => x65_out_1,
   I2 => x65_out_3,
   I3 => W_43_19_i_14_n_0,
   I4 => W_43_19_i_15_n_0,
   O => W_43_19_i_4_n_0
);
W_43_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x65_out_25,
   I1 => x65_out_0,
   I2 => x65_out_2,
   I3 => W_43_19_i_16_n_0,
   I4 => W_43_19_i_17_n_0,
   O => W_43_19_i_5_n_0
);
W_43_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_43_19_i_2_n_0,
   I1 => W_43_23_i_16_n_0,
   I2 => x65_out_29,
   I3 => x65_out_4,
   I4 => x65_out_6,
   I5 => W_43_23_i_17_n_0,
   O => W_43_19_i_6_n_0
);
W_43_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_43_19_i_3_n_0,
   I1 => W_43_19_i_10_n_0,
   I2 => x65_out_28,
   I3 => x65_out_3,
   I4 => x65_out_5,
   I5 => W_43_19_i_11_n_0,
   O => W_43_19_i_7_n_0
);
W_43_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_43_19_i_4_n_0,
   I1 => W_43_19_i_12_n_0,
   I2 => x65_out_27,
   I3 => x65_out_2,
   I4 => x65_out_4,
   I5 => W_43_19_i_13_n_0,
   O => W_43_19_i_8_n_0
);
W_43_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_43_19_i_5_n_0,
   I1 => W_43_19_i_14_n_0,
   I2 => x65_out_26,
   I3 => x65_out_1,
   I4 => x65_out_3,
   I5 => W_43_19_i_15_n_0,
   O => W_43_19_i_9_n_0
);
W_43_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x102_out_22,
   I1 => x80_out_22,
   I2 => x100_out_8,
   I3 => x100_out_29,
   I4 => x100_out_25,
   O => W_43_23_i_10_n_0
);
W_43_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x80_out_21,
   I1 => x100_out_24,
   I2 => x100_out_28,
   I3 => x100_out_7,
   I4 => x102_out_21,
   O => W_43_23_i_11_n_0
);
W_43_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x102_out_21,
   I1 => x80_out_21,
   I2 => x100_out_7,
   I3 => x100_out_28,
   I4 => x100_out_24,
   O => W_43_23_i_12_n_0
);
W_43_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x80_out_20,
   I1 => x100_out_23,
   I2 => x100_out_27,
   I3 => x100_out_6,
   I4 => x102_out_20,
   O => W_43_23_i_13_n_0
);
W_43_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x102_out_20,
   I1 => x80_out_20,
   I2 => x100_out_6,
   I3 => x100_out_27,
   I4 => x100_out_23,
   O => W_43_23_i_14_n_0
);
W_43_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x80_out_19,
   I1 => x100_out_22,
   I2 => x100_out_26,
   I3 => x100_out_5,
   I4 => x102_out_19,
   O => W_43_23_i_15_n_0
);
W_43_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x102_out_19,
   I1 => x80_out_19,
   I2 => x100_out_5,
   I3 => x100_out_26,
   I4 => x100_out_22,
   O => W_43_23_i_16_n_0
);
W_43_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x80_out_18,
   I1 => x100_out_21,
   I2 => x100_out_25,
   I3 => x100_out_4,
   I4 => x102_out_18,
   O => W_43_23_i_17_n_0
);
W_43_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x65_out_7,
   I1 => x65_out_9,
   I2 => W_43_23_i_10_n_0,
   I3 => W_43_23_i_11_n_0,
   O => W_43_23_i_2_n_0
);
W_43_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x65_out_31,
   I1 => x65_out_6,
   I2 => x65_out_8,
   I3 => W_43_23_i_12_n_0,
   I4 => W_43_23_i_13_n_0,
   O => W_43_23_i_3_n_0
);
W_43_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x65_out_30,
   I1 => x65_out_5,
   I2 => x65_out_7,
   I3 => W_43_23_i_14_n_0,
   I4 => W_43_23_i_15_n_0,
   O => W_43_23_i_4_n_0
);
W_43_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x65_out_29,
   I1 => x65_out_4,
   I2 => x65_out_6,
   I3 => W_43_23_i_16_n_0,
   I4 => W_43_23_i_17_n_0,
   O => W_43_23_i_5_n_0
);
W_43_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x65_out_8,
   I1 => x65_out_10,
   I2 => W_43_27_i_16_n_0,
   I3 => W_43_27_i_17_n_0,
   I4 => W_43_23_i_2_n_0,
   O => W_43_23_i_6_n_0
);
W_43_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x65_out_7,
   I1 => x65_out_9,
   I2 => W_43_23_i_10_n_0,
   I3 => W_43_23_i_11_n_0,
   I4 => W_43_23_i_3_n_0,
   O => W_43_23_i_7_n_0
);
W_43_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_43_23_i_4_n_0,
   I1 => W_43_23_i_12_n_0,
   I2 => x65_out_31,
   I3 => x65_out_6,
   I4 => x65_out_8,
   I5 => W_43_23_i_13_n_0,
   O => W_43_23_i_8_n_0
);
W_43_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_43_23_i_5_n_0,
   I1 => W_43_23_i_14_n_0,
   I2 => x65_out_30,
   I3 => x65_out_5,
   I4 => x65_out_7,
   I5 => W_43_23_i_15_n_0,
   O => W_43_23_i_9_n_0
);
W_43_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x102_out_26,
   I1 => x80_out_26,
   I2 => x100_out_12,
   I3 => x100_out_1,
   I4 => x100_out_29,
   O => W_43_27_i_10_n_0
);
W_43_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x80_out_25,
   I1 => x100_out_28,
   I2 => x100_out_0,
   I3 => x100_out_11,
   I4 => x102_out_25,
   O => W_43_27_i_11_n_0
);
W_43_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x102_out_25,
   I1 => x80_out_25,
   I2 => x100_out_11,
   I3 => x100_out_0,
   I4 => x100_out_28,
   O => W_43_27_i_12_n_0
);
W_43_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x80_out_24,
   I1 => x100_out_27,
   I2 => x100_out_31,
   I3 => x100_out_10,
   I4 => x102_out_24,
   O => W_43_27_i_13_n_0
);
W_43_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x102_out_24,
   I1 => x80_out_24,
   I2 => x100_out_10,
   I3 => x100_out_31,
   I4 => x100_out_27,
   O => W_43_27_i_14_n_0
);
W_43_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x80_out_23,
   I1 => x100_out_26,
   I2 => x100_out_30,
   I3 => x100_out_9,
   I4 => x102_out_23,
   O => W_43_27_i_15_n_0
);
W_43_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x102_out_23,
   I1 => x80_out_23,
   I2 => x100_out_9,
   I3 => x100_out_30,
   I4 => x100_out_26,
   O => W_43_27_i_16_n_0
);
W_43_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x80_out_22,
   I1 => x100_out_25,
   I2 => x100_out_29,
   I3 => x100_out_8,
   I4 => x102_out_22,
   O => W_43_27_i_17_n_0
);
W_43_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x65_out_11,
   I1 => x65_out_13,
   I2 => W_43_27_i_10_n_0,
   I3 => W_43_27_i_11_n_0,
   O => W_43_27_i_2_n_0
);
W_43_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x65_out_10,
   I1 => x65_out_12,
   I2 => W_43_27_i_12_n_0,
   I3 => W_43_27_i_13_n_0,
   O => W_43_27_i_3_n_0
);
W_43_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x65_out_9,
   I1 => x65_out_11,
   I2 => W_43_27_i_14_n_0,
   I3 => W_43_27_i_15_n_0,
   O => W_43_27_i_4_n_0
);
W_43_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x65_out_8,
   I1 => x65_out_10,
   I2 => W_43_27_i_16_n_0,
   I3 => W_43_27_i_17_n_0,
   O => W_43_27_i_5_n_0
);
W_43_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x65_out_12,
   I1 => x65_out_14,
   I2 => W_43_31_i_13_n_0,
   I3 => W_43_31_i_14_n_0,
   I4 => W_43_27_i_2_n_0,
   O => W_43_27_i_6_n_0
);
W_43_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x65_out_11,
   I1 => x65_out_13,
   I2 => W_43_27_i_10_n_0,
   I3 => W_43_27_i_11_n_0,
   I4 => W_43_27_i_3_n_0,
   O => W_43_27_i_7_n_0
);
W_43_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x65_out_10,
   I1 => x65_out_12,
   I2 => W_43_27_i_12_n_0,
   I3 => W_43_27_i_13_n_0,
   I4 => W_43_27_i_4_n_0,
   O => W_43_27_i_8_n_0
);
W_43_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x65_out_9,
   I1 => x65_out_11,
   I2 => W_43_27_i_14_n_0,
   I3 => W_43_27_i_15_n_0,
   I4 => W_43_27_i_5_n_0,
   O => W_43_27_i_9_n_0
);
W_43_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x80_out_28,
   I1 => x100_out_31,
   I2 => x100_out_3,
   I3 => x100_out_14,
   I4 => x102_out_28,
   O => W_43_31_i_10_n_0
);
W_43_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x102_out_28,
   I1 => x80_out_28,
   I2 => x100_out_14,
   I3 => x100_out_3,
   I4 => x100_out_31,
   O => W_43_31_i_11_n_0
);
W_43_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x80_out_27,
   I1 => x100_out_30,
   I2 => x100_out_2,
   I3 => x100_out_13,
   I4 => x102_out_27,
   O => W_43_31_i_12_n_0
);
W_43_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x102_out_27,
   I1 => x80_out_27,
   I2 => x100_out_13,
   I3 => x100_out_2,
   I4 => x100_out_30,
   O => W_43_31_i_13_n_0
);
W_43_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x80_out_26,
   I1 => x100_out_29,
   I2 => x100_out_1,
   I3 => x100_out_12,
   I4 => x102_out_26,
   O => W_43_31_i_14_n_0
);
W_43_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x80_out_29,
   I1 => x100_out_4,
   I2 => x100_out_15,
   I3 => x102_out_29,
   O => W_43_31_i_15_n_0
);
W_43_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x65_out_17,
   I1 => x65_out_15,
   O => SIGMA_LCASE_1171_out_0_30
);
W_43_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => x100_out_6,
   I1 => x100_out_17,
   I2 => x80_out_31,
   I3 => x102_out_31,
   I4 => x65_out_16,
   I5 => x65_out_18,
   O => W_43_31_i_17_n_0
);
W_43_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x100_out_16,
   I1 => x100_out_5,
   O => SIGMA_LCASE_0167_out_30
);
W_43_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x102_out_30,
   I1 => x80_out_30,
   I2 => x100_out_16,
   I3 => x100_out_5,
   O => W_43_31_i_19_n_0
);
W_43_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x65_out_14,
   I1 => x65_out_16,
   I2 => W_43_31_i_9_n_0,
   I3 => W_43_31_i_10_n_0,
   O => W_43_31_i_2_n_0
);
W_43_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x65_out_13,
   I1 => x65_out_15,
   I2 => W_43_31_i_11_n_0,
   I3 => W_43_31_i_12_n_0,
   O => W_43_31_i_3_n_0
);
W_43_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x65_out_12,
   I1 => x65_out_14,
   I2 => W_43_31_i_13_n_0,
   I3 => W_43_31_i_14_n_0,
   O => W_43_31_i_4_n_0
);
W_43_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_43_31_i_15_n_0,
   I1 => SIGMA_LCASE_1171_out_0_30,
   I2 => W_43_31_i_17_n_0,
   I3 => x80_out_30,
   I4 => SIGMA_LCASE_0167_out_30,
   I5 => x102_out_30,
   O => W_43_31_i_5_n_0
);
W_43_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_43_31_i_2_n_0,
   I1 => W_43_31_i_19_n_0,
   I2 => x65_out_15,
   I3 => x65_out_17,
   I4 => W_43_31_i_15_n_0,
   O => W_43_31_i_6_n_0
);
W_43_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x65_out_14,
   I1 => x65_out_16,
   I2 => W_43_31_i_9_n_0,
   I3 => W_43_31_i_10_n_0,
   I4 => W_43_31_i_3_n_0,
   O => W_43_31_i_7_n_0
);
W_43_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x65_out_13,
   I1 => x65_out_15,
   I2 => W_43_31_i_11_n_0,
   I3 => W_43_31_i_12_n_0,
   I4 => W_43_31_i_4_n_0,
   O => W_43_31_i_8_n_0
);
W_43_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x102_out_29,
   I1 => x80_out_29,
   I2 => x100_out_15,
   I3 => x100_out_4,
   O => W_43_31_i_9_n_0
);
W_43_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x102_out_2,
   I1 => x80_out_2,
   I2 => x100_out_20,
   I3 => x100_out_9,
   I4 => x100_out_5,
   O => W_43_3_i_10_n_0
);
W_43_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x80_out_1,
   I1 => x100_out_4,
   I2 => x100_out_8,
   I3 => x100_out_19,
   I4 => x102_out_1,
   O => W_43_3_i_11_n_0
);
W_43_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x100_out_19,
   I1 => x100_out_8,
   I2 => x100_out_4,
   O => SIGMA_LCASE_0167_out_1
);
W_43_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x65_out_21,
   I1 => x65_out_19,
   I2 => x65_out_12,
   O => SIGMA_LCASE_1171_out_0_2
);
W_43_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x65_out_20,
   I1 => x65_out_18,
   I2 => x65_out_11,
   O => SIGMA_LCASE_1171_out_1
);
W_43_3_i_15 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x102_out_1,
   I1 => x80_out_1,
   I2 => x100_out_19,
   I3 => x100_out_8,
   I4 => x100_out_4,
   O => W_43_3_i_15_n_0
);
W_43_3_i_16 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x100_out_18,
   I1 => x100_out_7,
   I2 => x100_out_3,
   O => SIGMA_LCASE_0167_out_0
);
W_43_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x65_out_12,
   I1 => x65_out_19,
   I2 => x65_out_21,
   I3 => W_43_3_i_10_n_0,
   I4 => W_43_3_i_11_n_0,
   O => W_43_3_i_2_n_0
);
W_43_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_43_3_i_11_n_0,
   I1 => x65_out_21,
   I2 => x65_out_19,
   I3 => x65_out_12,
   I4 => W_43_3_i_10_n_0,
   O => W_43_3_i_3_n_0
);
W_43_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_0167_out_1,
   I1 => x80_out_1,
   I2 => x102_out_1,
   I3 => x65_out_11,
   I4 => x65_out_18,
   I5 => x65_out_20,
   O => W_43_3_i_4_n_0
);
W_43_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x102_out_0,
   I1 => x80_out_0,
   I2 => x100_out_18,
   I3 => x100_out_7,
   I4 => x100_out_3,
   O => W_43_3_i_5_n_0
);
W_43_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_43_3_i_2_n_0,
   I1 => W_43_7_i_16_n_0,
   I2 => x65_out_13,
   I3 => x65_out_20,
   I4 => x65_out_22,
   I5 => W_43_7_i_17_n_0,
   O => W_43_3_i_6_n_0
);
W_43_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_43_3_i_10_n_0,
   I1 => SIGMA_LCASE_1171_out_0_2,
   I2 => x102_out_1,
   I3 => x80_out_1,
   I4 => SIGMA_LCASE_0167_out_1,
   I5 => SIGMA_LCASE_1171_out_1,
   O => W_43_3_i_7_n_0
);
W_43_3_i_8 : LUT5
  generic map(
   INIT => X"99969666"
  )
 port map (
   I0 => SIGMA_LCASE_1171_out_1,
   I1 => W_43_3_i_15_n_0,
   I2 => x102_out_0,
   I3 => SIGMA_LCASE_0167_out_0,
   I4 => x80_out_0,
   O => W_43_3_i_8_n_0
);
W_43_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_43_3_i_5_n_0,
   I1 => x65_out_10,
   I2 => x65_out_17,
   I3 => x65_out_19,
   O => W_43_3_i_9_n_0
);
W_43_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x102_out_6,
   I1 => x80_out_6,
   I2 => x100_out_24,
   I3 => x100_out_13,
   I4 => x100_out_9,
   O => W_43_7_i_10_n_0
);
W_43_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x80_out_5,
   I1 => x100_out_8,
   I2 => x100_out_12,
   I3 => x100_out_23,
   I4 => x102_out_5,
   O => W_43_7_i_11_n_0
);
W_43_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x102_out_5,
   I1 => x80_out_5,
   I2 => x100_out_23,
   I3 => x100_out_12,
   I4 => x100_out_8,
   O => W_43_7_i_12_n_0
);
W_43_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x80_out_4,
   I1 => x100_out_7,
   I2 => x100_out_11,
   I3 => x100_out_22,
   I4 => x102_out_4,
   O => W_43_7_i_13_n_0
);
W_43_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x102_out_4,
   I1 => x80_out_4,
   I2 => x100_out_22,
   I3 => x100_out_11,
   I4 => x100_out_7,
   O => W_43_7_i_14_n_0
);
W_43_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x80_out_3,
   I1 => x100_out_6,
   I2 => x100_out_10,
   I3 => x100_out_21,
   I4 => x102_out_3,
   O => W_43_7_i_15_n_0
);
W_43_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x102_out_3,
   I1 => x80_out_3,
   I2 => x100_out_21,
   I3 => x100_out_10,
   I4 => x100_out_6,
   O => W_43_7_i_16_n_0
);
W_43_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x80_out_2,
   I1 => x100_out_5,
   I2 => x100_out_9,
   I3 => x100_out_20,
   I4 => x102_out_2,
   O => W_43_7_i_17_n_0
);
W_43_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x65_out_16,
   I1 => x65_out_23,
   I2 => x65_out_25,
   I3 => W_43_7_i_10_n_0,
   I4 => W_43_7_i_11_n_0,
   O => W_43_7_i_2_n_0
);
W_43_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x65_out_15,
   I1 => x65_out_22,
   I2 => x65_out_24,
   I3 => W_43_7_i_12_n_0,
   I4 => W_43_7_i_13_n_0,
   O => W_43_7_i_3_n_0
);
W_43_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x65_out_14,
   I1 => x65_out_21,
   I2 => x65_out_23,
   I3 => W_43_7_i_14_n_0,
   I4 => W_43_7_i_15_n_0,
   O => W_43_7_i_4_n_0
);
W_43_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x65_out_13,
   I1 => x65_out_20,
   I2 => x65_out_22,
   I3 => W_43_7_i_16_n_0,
   I4 => W_43_7_i_17_n_0,
   O => W_43_7_i_5_n_0
);
W_43_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_43_7_i_2_n_0,
   I1 => W_43_11_i_16_n_0,
   I2 => x65_out_17,
   I3 => x65_out_24,
   I4 => x65_out_26,
   I5 => W_43_11_i_17_n_0,
   O => W_43_7_i_6_n_0
);
W_43_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_43_7_i_3_n_0,
   I1 => W_43_7_i_10_n_0,
   I2 => x65_out_16,
   I3 => x65_out_23,
   I4 => x65_out_25,
   I5 => W_43_7_i_11_n_0,
   O => W_43_7_i_7_n_0
);
W_43_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_43_7_i_4_n_0,
   I1 => W_43_7_i_12_n_0,
   I2 => x65_out_15,
   I3 => x65_out_22,
   I4 => x65_out_24,
   I5 => W_43_7_i_13_n_0,
   O => W_43_7_i_8_n_0
);
W_43_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_43_7_i_5_n_0,
   I1 => W_43_7_i_14_n_0,
   I2 => x65_out_14,
   I3 => x65_out_21,
   I4 => x65_out_23,
   I5 => W_43_7_i_15_n_0,
   O => W_43_7_i_9_n_0
);
W_44_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x100_out_10,
   I1 => x77_out_10,
   I2 => x98_out_28,
   I3 => x98_out_17,
   I4 => x98_out_13,
   O => W_44_11_i_10_n_0
);
W_44_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x77_out_9,
   I1 => x98_out_12,
   I2 => x98_out_16,
   I3 => x98_out_27,
   I4 => x100_out_9,
   O => W_44_11_i_11_n_0
);
W_44_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x100_out_9,
   I1 => x77_out_9,
   I2 => x98_out_27,
   I3 => x98_out_16,
   I4 => x98_out_12,
   O => W_44_11_i_12_n_0
);
W_44_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x77_out_8,
   I1 => x98_out_11,
   I2 => x98_out_15,
   I3 => x98_out_26,
   I4 => x100_out_8,
   O => W_44_11_i_13_n_0
);
W_44_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x100_out_8,
   I1 => x77_out_8,
   I2 => x98_out_26,
   I3 => x98_out_15,
   I4 => x98_out_11,
   O => W_44_11_i_14_n_0
);
W_44_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x77_out_7,
   I1 => x98_out_10,
   I2 => x98_out_14,
   I3 => x98_out_25,
   I4 => x100_out_7,
   O => W_44_11_i_15_n_0
);
W_44_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x100_out_7,
   I1 => x77_out_7,
   I2 => x98_out_25,
   I3 => x98_out_14,
   I4 => x98_out_10,
   O => W_44_11_i_16_n_0
);
W_44_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x77_out_6,
   I1 => x98_out_9,
   I2 => x98_out_13,
   I3 => x98_out_24,
   I4 => x100_out_6,
   O => W_44_11_i_17_n_0
);
W_44_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x62_out_20,
   I1 => x62_out_27,
   I2 => x62_out_29,
   I3 => W_44_11_i_10_n_0,
   I4 => W_44_11_i_11_n_0,
   O => W_44_11_i_2_n_0
);
W_44_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x62_out_19,
   I1 => x62_out_26,
   I2 => x62_out_28,
   I3 => W_44_11_i_12_n_0,
   I4 => W_44_11_i_13_n_0,
   O => W_44_11_i_3_n_0
);
W_44_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x62_out_18,
   I1 => x62_out_25,
   I2 => x62_out_27,
   I3 => W_44_11_i_14_n_0,
   I4 => W_44_11_i_15_n_0,
   O => W_44_11_i_4_n_0
);
W_44_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x62_out_17,
   I1 => x62_out_24,
   I2 => x62_out_26,
   I3 => W_44_11_i_16_n_0,
   I4 => W_44_11_i_17_n_0,
   O => W_44_11_i_5_n_0
);
W_44_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_44_11_i_2_n_0,
   I1 => W_44_15_i_16_n_0,
   I2 => x62_out_21,
   I3 => x62_out_28,
   I4 => x62_out_30,
   I5 => W_44_15_i_17_n_0,
   O => W_44_11_i_6_n_0
);
W_44_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_44_11_i_3_n_0,
   I1 => W_44_11_i_10_n_0,
   I2 => x62_out_20,
   I3 => x62_out_27,
   I4 => x62_out_29,
   I5 => W_44_11_i_11_n_0,
   O => W_44_11_i_7_n_0
);
W_44_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_44_11_i_4_n_0,
   I1 => W_44_11_i_12_n_0,
   I2 => x62_out_19,
   I3 => x62_out_26,
   I4 => x62_out_28,
   I5 => W_44_11_i_13_n_0,
   O => W_44_11_i_8_n_0
);
W_44_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_44_11_i_5_n_0,
   I1 => W_44_11_i_14_n_0,
   I2 => x62_out_18,
   I3 => x62_out_25,
   I4 => x62_out_27,
   I5 => W_44_11_i_15_n_0,
   O => W_44_11_i_9_n_0
);
W_44_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x100_out_14,
   I1 => x77_out_14,
   I2 => x98_out_0,
   I3 => x98_out_21,
   I4 => x98_out_17,
   O => W_44_15_i_10_n_0
);
W_44_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x77_out_13,
   I1 => x98_out_16,
   I2 => x98_out_20,
   I3 => x98_out_31,
   I4 => x100_out_13,
   O => W_44_15_i_11_n_0
);
W_44_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x100_out_13,
   I1 => x77_out_13,
   I2 => x98_out_31,
   I3 => x98_out_20,
   I4 => x98_out_16,
   O => W_44_15_i_12_n_0
);
W_44_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x77_out_12,
   I1 => x98_out_15,
   I2 => x98_out_19,
   I3 => x98_out_30,
   I4 => x100_out_12,
   O => W_44_15_i_13_n_0
);
W_44_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x100_out_12,
   I1 => x77_out_12,
   I2 => x98_out_30,
   I3 => x98_out_19,
   I4 => x98_out_15,
   O => W_44_15_i_14_n_0
);
W_44_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x77_out_11,
   I1 => x98_out_14,
   I2 => x98_out_18,
   I3 => x98_out_29,
   I4 => x100_out_11,
   O => W_44_15_i_15_n_0
);
W_44_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x100_out_11,
   I1 => x77_out_11,
   I2 => x98_out_29,
   I3 => x98_out_18,
   I4 => x98_out_14,
   O => W_44_15_i_16_n_0
);
W_44_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x77_out_10,
   I1 => x98_out_13,
   I2 => x98_out_17,
   I3 => x98_out_28,
   I4 => x100_out_10,
   O => W_44_15_i_17_n_0
);
W_44_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x62_out_24,
   I1 => x62_out_31,
   I2 => x62_out_1,
   I3 => W_44_15_i_10_n_0,
   I4 => W_44_15_i_11_n_0,
   O => W_44_15_i_2_n_0
);
W_44_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x62_out_23,
   I1 => x62_out_30,
   I2 => x62_out_0,
   I3 => W_44_15_i_12_n_0,
   I4 => W_44_15_i_13_n_0,
   O => W_44_15_i_3_n_0
);
W_44_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x62_out_22,
   I1 => x62_out_29,
   I2 => x62_out_31,
   I3 => W_44_15_i_14_n_0,
   I4 => W_44_15_i_15_n_0,
   O => W_44_15_i_4_n_0
);
W_44_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x62_out_21,
   I1 => x62_out_28,
   I2 => x62_out_30,
   I3 => W_44_15_i_16_n_0,
   I4 => W_44_15_i_17_n_0,
   O => W_44_15_i_5_n_0
);
W_44_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_44_15_i_2_n_0,
   I1 => W_44_19_i_16_n_0,
   I2 => x62_out_25,
   I3 => x62_out_0,
   I4 => x62_out_2,
   I5 => W_44_19_i_17_n_0,
   O => W_44_15_i_6_n_0
);
W_44_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_44_15_i_3_n_0,
   I1 => W_44_15_i_10_n_0,
   I2 => x62_out_24,
   I3 => x62_out_31,
   I4 => x62_out_1,
   I5 => W_44_15_i_11_n_0,
   O => W_44_15_i_7_n_0
);
W_44_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_44_15_i_4_n_0,
   I1 => W_44_15_i_12_n_0,
   I2 => x62_out_23,
   I3 => x62_out_30,
   I4 => x62_out_0,
   I5 => W_44_15_i_13_n_0,
   O => W_44_15_i_8_n_0
);
W_44_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_44_15_i_5_n_0,
   I1 => W_44_15_i_14_n_0,
   I2 => x62_out_22,
   I3 => x62_out_29,
   I4 => x62_out_31,
   I5 => W_44_15_i_15_n_0,
   O => W_44_15_i_9_n_0
);
W_44_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x100_out_18,
   I1 => x77_out_18,
   I2 => x98_out_4,
   I3 => x98_out_25,
   I4 => x98_out_21,
   O => W_44_19_i_10_n_0
);
W_44_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x77_out_17,
   I1 => x98_out_20,
   I2 => x98_out_24,
   I3 => x98_out_3,
   I4 => x100_out_17,
   O => W_44_19_i_11_n_0
);
W_44_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x100_out_17,
   I1 => x77_out_17,
   I2 => x98_out_3,
   I3 => x98_out_24,
   I4 => x98_out_20,
   O => W_44_19_i_12_n_0
);
W_44_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x77_out_16,
   I1 => x98_out_19,
   I2 => x98_out_23,
   I3 => x98_out_2,
   I4 => x100_out_16,
   O => W_44_19_i_13_n_0
);
W_44_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x100_out_16,
   I1 => x77_out_16,
   I2 => x98_out_2,
   I3 => x98_out_23,
   I4 => x98_out_19,
   O => W_44_19_i_14_n_0
);
W_44_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x77_out_15,
   I1 => x98_out_18,
   I2 => x98_out_22,
   I3 => x98_out_1,
   I4 => x100_out_15,
   O => W_44_19_i_15_n_0
);
W_44_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x100_out_15,
   I1 => x77_out_15,
   I2 => x98_out_1,
   I3 => x98_out_22,
   I4 => x98_out_18,
   O => W_44_19_i_16_n_0
);
W_44_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x77_out_14,
   I1 => x98_out_17,
   I2 => x98_out_21,
   I3 => x98_out_0,
   I4 => x100_out_14,
   O => W_44_19_i_17_n_0
);
W_44_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x62_out_28,
   I1 => x62_out_3,
   I2 => x62_out_5,
   I3 => W_44_19_i_10_n_0,
   I4 => W_44_19_i_11_n_0,
   O => W_44_19_i_2_n_0
);
W_44_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x62_out_27,
   I1 => x62_out_2,
   I2 => x62_out_4,
   I3 => W_44_19_i_12_n_0,
   I4 => W_44_19_i_13_n_0,
   O => W_44_19_i_3_n_0
);
W_44_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x62_out_26,
   I1 => x62_out_1,
   I2 => x62_out_3,
   I3 => W_44_19_i_14_n_0,
   I4 => W_44_19_i_15_n_0,
   O => W_44_19_i_4_n_0
);
W_44_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x62_out_25,
   I1 => x62_out_0,
   I2 => x62_out_2,
   I3 => W_44_19_i_16_n_0,
   I4 => W_44_19_i_17_n_0,
   O => W_44_19_i_5_n_0
);
W_44_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_44_19_i_2_n_0,
   I1 => W_44_23_i_16_n_0,
   I2 => x62_out_29,
   I3 => x62_out_4,
   I4 => x62_out_6,
   I5 => W_44_23_i_17_n_0,
   O => W_44_19_i_6_n_0
);
W_44_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_44_19_i_3_n_0,
   I1 => W_44_19_i_10_n_0,
   I2 => x62_out_28,
   I3 => x62_out_3,
   I4 => x62_out_5,
   I5 => W_44_19_i_11_n_0,
   O => W_44_19_i_7_n_0
);
W_44_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_44_19_i_4_n_0,
   I1 => W_44_19_i_12_n_0,
   I2 => x62_out_27,
   I3 => x62_out_2,
   I4 => x62_out_4,
   I5 => W_44_19_i_13_n_0,
   O => W_44_19_i_8_n_0
);
W_44_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_44_19_i_5_n_0,
   I1 => W_44_19_i_14_n_0,
   I2 => x62_out_26,
   I3 => x62_out_1,
   I4 => x62_out_3,
   I5 => W_44_19_i_15_n_0,
   O => W_44_19_i_9_n_0
);
W_44_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x100_out_22,
   I1 => x77_out_22,
   I2 => x98_out_8,
   I3 => x98_out_29,
   I4 => x98_out_25,
   O => W_44_23_i_10_n_0
);
W_44_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x77_out_21,
   I1 => x98_out_24,
   I2 => x98_out_28,
   I3 => x98_out_7,
   I4 => x100_out_21,
   O => W_44_23_i_11_n_0
);
W_44_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x100_out_21,
   I1 => x77_out_21,
   I2 => x98_out_7,
   I3 => x98_out_28,
   I4 => x98_out_24,
   O => W_44_23_i_12_n_0
);
W_44_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x77_out_20,
   I1 => x98_out_23,
   I2 => x98_out_27,
   I3 => x98_out_6,
   I4 => x100_out_20,
   O => W_44_23_i_13_n_0
);
W_44_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x100_out_20,
   I1 => x77_out_20,
   I2 => x98_out_6,
   I3 => x98_out_27,
   I4 => x98_out_23,
   O => W_44_23_i_14_n_0
);
W_44_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x77_out_19,
   I1 => x98_out_22,
   I2 => x98_out_26,
   I3 => x98_out_5,
   I4 => x100_out_19,
   O => W_44_23_i_15_n_0
);
W_44_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x100_out_19,
   I1 => x77_out_19,
   I2 => x98_out_5,
   I3 => x98_out_26,
   I4 => x98_out_22,
   O => W_44_23_i_16_n_0
);
W_44_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x77_out_18,
   I1 => x98_out_21,
   I2 => x98_out_25,
   I3 => x98_out_4,
   I4 => x100_out_18,
   O => W_44_23_i_17_n_0
);
W_44_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x62_out_7,
   I1 => x62_out_9,
   I2 => W_44_23_i_10_n_0,
   I3 => W_44_23_i_11_n_0,
   O => W_44_23_i_2_n_0
);
W_44_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x62_out_31,
   I1 => x62_out_6,
   I2 => x62_out_8,
   I3 => W_44_23_i_12_n_0,
   I4 => W_44_23_i_13_n_0,
   O => W_44_23_i_3_n_0
);
W_44_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x62_out_30,
   I1 => x62_out_5,
   I2 => x62_out_7,
   I3 => W_44_23_i_14_n_0,
   I4 => W_44_23_i_15_n_0,
   O => W_44_23_i_4_n_0
);
W_44_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x62_out_29,
   I1 => x62_out_4,
   I2 => x62_out_6,
   I3 => W_44_23_i_16_n_0,
   I4 => W_44_23_i_17_n_0,
   O => W_44_23_i_5_n_0
);
W_44_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x62_out_8,
   I1 => x62_out_10,
   I2 => W_44_27_i_16_n_0,
   I3 => W_44_27_i_17_n_0,
   I4 => W_44_23_i_2_n_0,
   O => W_44_23_i_6_n_0
);
W_44_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x62_out_7,
   I1 => x62_out_9,
   I2 => W_44_23_i_10_n_0,
   I3 => W_44_23_i_11_n_0,
   I4 => W_44_23_i_3_n_0,
   O => W_44_23_i_7_n_0
);
W_44_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_44_23_i_4_n_0,
   I1 => W_44_23_i_12_n_0,
   I2 => x62_out_31,
   I3 => x62_out_6,
   I4 => x62_out_8,
   I5 => W_44_23_i_13_n_0,
   O => W_44_23_i_8_n_0
);
W_44_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_44_23_i_5_n_0,
   I1 => W_44_23_i_14_n_0,
   I2 => x62_out_30,
   I3 => x62_out_5,
   I4 => x62_out_7,
   I5 => W_44_23_i_15_n_0,
   O => W_44_23_i_9_n_0
);
W_44_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x100_out_26,
   I1 => x77_out_26,
   I2 => x98_out_12,
   I3 => x98_out_1,
   I4 => x98_out_29,
   O => W_44_27_i_10_n_0
);
W_44_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x77_out_25,
   I1 => x98_out_28,
   I2 => x98_out_0,
   I3 => x98_out_11,
   I4 => x100_out_25,
   O => W_44_27_i_11_n_0
);
W_44_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x100_out_25,
   I1 => x77_out_25,
   I2 => x98_out_11,
   I3 => x98_out_0,
   I4 => x98_out_28,
   O => W_44_27_i_12_n_0
);
W_44_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x77_out_24,
   I1 => x98_out_27,
   I2 => x98_out_31,
   I3 => x98_out_10,
   I4 => x100_out_24,
   O => W_44_27_i_13_n_0
);
W_44_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x100_out_24,
   I1 => x77_out_24,
   I2 => x98_out_10,
   I3 => x98_out_31,
   I4 => x98_out_27,
   O => W_44_27_i_14_n_0
);
W_44_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x77_out_23,
   I1 => x98_out_26,
   I2 => x98_out_30,
   I3 => x98_out_9,
   I4 => x100_out_23,
   O => W_44_27_i_15_n_0
);
W_44_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x100_out_23,
   I1 => x77_out_23,
   I2 => x98_out_9,
   I3 => x98_out_30,
   I4 => x98_out_26,
   O => W_44_27_i_16_n_0
);
W_44_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x77_out_22,
   I1 => x98_out_25,
   I2 => x98_out_29,
   I3 => x98_out_8,
   I4 => x100_out_22,
   O => W_44_27_i_17_n_0
);
W_44_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x62_out_11,
   I1 => x62_out_13,
   I2 => W_44_27_i_10_n_0,
   I3 => W_44_27_i_11_n_0,
   O => W_44_27_i_2_n_0
);
W_44_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x62_out_10,
   I1 => x62_out_12,
   I2 => W_44_27_i_12_n_0,
   I3 => W_44_27_i_13_n_0,
   O => W_44_27_i_3_n_0
);
W_44_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x62_out_9,
   I1 => x62_out_11,
   I2 => W_44_27_i_14_n_0,
   I3 => W_44_27_i_15_n_0,
   O => W_44_27_i_4_n_0
);
W_44_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x62_out_8,
   I1 => x62_out_10,
   I2 => W_44_27_i_16_n_0,
   I3 => W_44_27_i_17_n_0,
   O => W_44_27_i_5_n_0
);
W_44_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x62_out_12,
   I1 => x62_out_14,
   I2 => W_44_31_i_13_n_0,
   I3 => W_44_31_i_14_n_0,
   I4 => W_44_27_i_2_n_0,
   O => W_44_27_i_6_n_0
);
W_44_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x62_out_11,
   I1 => x62_out_13,
   I2 => W_44_27_i_10_n_0,
   I3 => W_44_27_i_11_n_0,
   I4 => W_44_27_i_3_n_0,
   O => W_44_27_i_7_n_0
);
W_44_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x62_out_10,
   I1 => x62_out_12,
   I2 => W_44_27_i_12_n_0,
   I3 => W_44_27_i_13_n_0,
   I4 => W_44_27_i_4_n_0,
   O => W_44_27_i_8_n_0
);
W_44_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x62_out_9,
   I1 => x62_out_11,
   I2 => W_44_27_i_14_n_0,
   I3 => W_44_27_i_15_n_0,
   I4 => W_44_27_i_5_n_0,
   O => W_44_27_i_9_n_0
);
W_44_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x77_out_28,
   I1 => x98_out_31,
   I2 => x98_out_3,
   I3 => x98_out_14,
   I4 => x100_out_28,
   O => W_44_31_i_10_n_0
);
W_44_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x100_out_28,
   I1 => x77_out_28,
   I2 => x98_out_14,
   I3 => x98_out_3,
   I4 => x98_out_31,
   O => W_44_31_i_11_n_0
);
W_44_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x77_out_27,
   I1 => x98_out_30,
   I2 => x98_out_2,
   I3 => x98_out_13,
   I4 => x100_out_27,
   O => W_44_31_i_12_n_0
);
W_44_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x100_out_27,
   I1 => x77_out_27,
   I2 => x98_out_13,
   I3 => x98_out_2,
   I4 => x98_out_30,
   O => W_44_31_i_13_n_0
);
W_44_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x77_out_26,
   I1 => x98_out_29,
   I2 => x98_out_1,
   I3 => x98_out_12,
   I4 => x100_out_26,
   O => W_44_31_i_14_n_0
);
W_44_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x77_out_29,
   I1 => x98_out_4,
   I2 => x98_out_15,
   I3 => x100_out_29,
   O => W_44_31_i_15_n_0
);
W_44_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x62_out_17,
   I1 => x62_out_15,
   O => SIGMA_LCASE_1163_out_0_30
);
W_44_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => x98_out_6,
   I1 => x98_out_17,
   I2 => x77_out_31,
   I3 => x100_out_31,
   I4 => x62_out_16,
   I5 => x62_out_18,
   O => W_44_31_i_17_n_0
);
W_44_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x98_out_16,
   I1 => x98_out_5,
   O => SIGMA_LCASE_0159_out_30
);
W_44_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x100_out_30,
   I1 => x77_out_30,
   I2 => x98_out_16,
   I3 => x98_out_5,
   O => W_44_31_i_19_n_0
);
W_44_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x62_out_14,
   I1 => x62_out_16,
   I2 => W_44_31_i_9_n_0,
   I3 => W_44_31_i_10_n_0,
   O => W_44_31_i_2_n_0
);
W_44_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x62_out_13,
   I1 => x62_out_15,
   I2 => W_44_31_i_11_n_0,
   I3 => W_44_31_i_12_n_0,
   O => W_44_31_i_3_n_0
);
W_44_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x62_out_12,
   I1 => x62_out_14,
   I2 => W_44_31_i_13_n_0,
   I3 => W_44_31_i_14_n_0,
   O => W_44_31_i_4_n_0
);
W_44_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_44_31_i_15_n_0,
   I1 => SIGMA_LCASE_1163_out_0_30,
   I2 => W_44_31_i_17_n_0,
   I3 => x77_out_30,
   I4 => SIGMA_LCASE_0159_out_30,
   I5 => x100_out_30,
   O => W_44_31_i_5_n_0
);
W_44_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_44_31_i_2_n_0,
   I1 => W_44_31_i_19_n_0,
   I2 => x62_out_15,
   I3 => x62_out_17,
   I4 => W_44_31_i_15_n_0,
   O => W_44_31_i_6_n_0
);
W_44_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x62_out_14,
   I1 => x62_out_16,
   I2 => W_44_31_i_9_n_0,
   I3 => W_44_31_i_10_n_0,
   I4 => W_44_31_i_3_n_0,
   O => W_44_31_i_7_n_0
);
W_44_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x62_out_13,
   I1 => x62_out_15,
   I2 => W_44_31_i_11_n_0,
   I3 => W_44_31_i_12_n_0,
   I4 => W_44_31_i_4_n_0,
   O => W_44_31_i_8_n_0
);
W_44_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x100_out_29,
   I1 => x77_out_29,
   I2 => x98_out_15,
   I3 => x98_out_4,
   O => W_44_31_i_9_n_0
);
W_44_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x100_out_2,
   I1 => x77_out_2,
   I2 => x98_out_20,
   I3 => x98_out_9,
   I4 => x98_out_5,
   O => W_44_3_i_10_n_0
);
W_44_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x77_out_1,
   I1 => x98_out_4,
   I2 => x98_out_8,
   I3 => x98_out_19,
   I4 => x100_out_1,
   O => W_44_3_i_11_n_0
);
W_44_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x98_out_19,
   I1 => x98_out_8,
   I2 => x98_out_4,
   O => SIGMA_LCASE_0159_out_1
);
W_44_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x62_out_21,
   I1 => x62_out_19,
   I2 => x62_out_12,
   O => SIGMA_LCASE_1163_out_0_2
);
W_44_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x62_out_20,
   I1 => x62_out_18,
   I2 => x62_out_11,
   O => SIGMA_LCASE_1163_out_1
);
W_44_3_i_15 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x100_out_1,
   I1 => x77_out_1,
   I2 => x98_out_19,
   I3 => x98_out_8,
   I4 => x98_out_4,
   O => W_44_3_i_15_n_0
);
W_44_3_i_16 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x98_out_18,
   I1 => x98_out_7,
   I2 => x98_out_3,
   O => SIGMA_LCASE_0159_out_0
);
W_44_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x62_out_12,
   I1 => x62_out_19,
   I2 => x62_out_21,
   I3 => W_44_3_i_10_n_0,
   I4 => W_44_3_i_11_n_0,
   O => W_44_3_i_2_n_0
);
W_44_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_44_3_i_11_n_0,
   I1 => x62_out_21,
   I2 => x62_out_19,
   I3 => x62_out_12,
   I4 => W_44_3_i_10_n_0,
   O => W_44_3_i_3_n_0
);
W_44_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_0159_out_1,
   I1 => x77_out_1,
   I2 => x100_out_1,
   I3 => x62_out_11,
   I4 => x62_out_18,
   I5 => x62_out_20,
   O => W_44_3_i_4_n_0
);
W_44_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x100_out_0,
   I1 => x77_out_0,
   I2 => x98_out_18,
   I3 => x98_out_7,
   I4 => x98_out_3,
   O => W_44_3_i_5_n_0
);
W_44_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_44_3_i_2_n_0,
   I1 => W_44_7_i_16_n_0,
   I2 => x62_out_13,
   I3 => x62_out_20,
   I4 => x62_out_22,
   I5 => W_44_7_i_17_n_0,
   O => W_44_3_i_6_n_0
);
W_44_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_44_3_i_10_n_0,
   I1 => SIGMA_LCASE_1163_out_0_2,
   I2 => x100_out_1,
   I3 => x77_out_1,
   I4 => SIGMA_LCASE_0159_out_1,
   I5 => SIGMA_LCASE_1163_out_1,
   O => W_44_3_i_7_n_0
);
W_44_3_i_8 : LUT5
  generic map(
   INIT => X"99969666"
  )
 port map (
   I0 => SIGMA_LCASE_1163_out_1,
   I1 => W_44_3_i_15_n_0,
   I2 => x100_out_0,
   I3 => SIGMA_LCASE_0159_out_0,
   I4 => x77_out_0,
   O => W_44_3_i_8_n_0
);
W_44_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_44_3_i_5_n_0,
   I1 => x62_out_10,
   I2 => x62_out_17,
   I3 => x62_out_19,
   O => W_44_3_i_9_n_0
);
W_44_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x100_out_6,
   I1 => x77_out_6,
   I2 => x98_out_24,
   I3 => x98_out_13,
   I4 => x98_out_9,
   O => W_44_7_i_10_n_0
);
W_44_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x77_out_5,
   I1 => x98_out_8,
   I2 => x98_out_12,
   I3 => x98_out_23,
   I4 => x100_out_5,
   O => W_44_7_i_11_n_0
);
W_44_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x100_out_5,
   I1 => x77_out_5,
   I2 => x98_out_23,
   I3 => x98_out_12,
   I4 => x98_out_8,
   O => W_44_7_i_12_n_0
);
W_44_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x77_out_4,
   I1 => x98_out_7,
   I2 => x98_out_11,
   I3 => x98_out_22,
   I4 => x100_out_4,
   O => W_44_7_i_13_n_0
);
W_44_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x100_out_4,
   I1 => x77_out_4,
   I2 => x98_out_22,
   I3 => x98_out_11,
   I4 => x98_out_7,
   O => W_44_7_i_14_n_0
);
W_44_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x77_out_3,
   I1 => x98_out_6,
   I2 => x98_out_10,
   I3 => x98_out_21,
   I4 => x100_out_3,
   O => W_44_7_i_15_n_0
);
W_44_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x100_out_3,
   I1 => x77_out_3,
   I2 => x98_out_21,
   I3 => x98_out_10,
   I4 => x98_out_6,
   O => W_44_7_i_16_n_0
);
W_44_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x77_out_2,
   I1 => x98_out_5,
   I2 => x98_out_9,
   I3 => x98_out_20,
   I4 => x100_out_2,
   O => W_44_7_i_17_n_0
);
W_44_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x62_out_16,
   I1 => x62_out_23,
   I2 => x62_out_25,
   I3 => W_44_7_i_10_n_0,
   I4 => W_44_7_i_11_n_0,
   O => W_44_7_i_2_n_0
);
W_44_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x62_out_15,
   I1 => x62_out_22,
   I2 => x62_out_24,
   I3 => W_44_7_i_12_n_0,
   I4 => W_44_7_i_13_n_0,
   O => W_44_7_i_3_n_0
);
W_44_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x62_out_14,
   I1 => x62_out_21,
   I2 => x62_out_23,
   I3 => W_44_7_i_14_n_0,
   I4 => W_44_7_i_15_n_0,
   O => W_44_7_i_4_n_0
);
W_44_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x62_out_13,
   I1 => x62_out_20,
   I2 => x62_out_22,
   I3 => W_44_7_i_16_n_0,
   I4 => W_44_7_i_17_n_0,
   O => W_44_7_i_5_n_0
);
W_44_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_44_7_i_2_n_0,
   I1 => W_44_11_i_16_n_0,
   I2 => x62_out_17,
   I3 => x62_out_24,
   I4 => x62_out_26,
   I5 => W_44_11_i_17_n_0,
   O => W_44_7_i_6_n_0
);
W_44_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_44_7_i_3_n_0,
   I1 => W_44_7_i_10_n_0,
   I2 => x62_out_16,
   I3 => x62_out_23,
   I4 => x62_out_25,
   I5 => W_44_7_i_11_n_0,
   O => W_44_7_i_7_n_0
);
W_44_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_44_7_i_4_n_0,
   I1 => W_44_7_i_12_n_0,
   I2 => x62_out_15,
   I3 => x62_out_22,
   I4 => x62_out_24,
   I5 => W_44_7_i_13_n_0,
   O => W_44_7_i_8_n_0
);
W_44_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_44_7_i_5_n_0,
   I1 => W_44_7_i_14_n_0,
   I2 => x62_out_14,
   I3 => x62_out_21,
   I4 => x62_out_23,
   I5 => W_44_7_i_15_n_0,
   O => W_44_7_i_9_n_0
);
W_45_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x98_out_10,
   I1 => x74_out_10,
   I2 => x96_out_28,
   I3 => x96_out_17,
   I4 => x96_out_13,
   O => W_45_11_i_10_n_0
);
W_45_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x74_out_9,
   I1 => x96_out_12,
   I2 => x96_out_16,
   I3 => x96_out_27,
   I4 => x98_out_9,
   O => W_45_11_i_11_n_0
);
W_45_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x98_out_9,
   I1 => x74_out_9,
   I2 => x96_out_27,
   I3 => x96_out_16,
   I4 => x96_out_12,
   O => W_45_11_i_12_n_0
);
W_45_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x74_out_8,
   I1 => x96_out_11,
   I2 => x96_out_15,
   I3 => x96_out_26,
   I4 => x98_out_8,
   O => W_45_11_i_13_n_0
);
W_45_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x98_out_8,
   I1 => x74_out_8,
   I2 => x96_out_26,
   I3 => x96_out_15,
   I4 => x96_out_11,
   O => W_45_11_i_14_n_0
);
W_45_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x74_out_7,
   I1 => x96_out_10,
   I2 => x96_out_14,
   I3 => x96_out_25,
   I4 => x98_out_7,
   O => W_45_11_i_15_n_0
);
W_45_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x98_out_7,
   I1 => x74_out_7,
   I2 => x96_out_25,
   I3 => x96_out_14,
   I4 => x96_out_10,
   O => W_45_11_i_16_n_0
);
W_45_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x74_out_6,
   I1 => x96_out_9,
   I2 => x96_out_13,
   I3 => x96_out_24,
   I4 => x98_out_6,
   O => W_45_11_i_17_n_0
);
W_45_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x59_out_20,
   I1 => x59_out_27,
   I2 => x59_out_29,
   I3 => W_45_11_i_10_n_0,
   I4 => W_45_11_i_11_n_0,
   O => W_45_11_i_2_n_0
);
W_45_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x59_out_19,
   I1 => x59_out_26,
   I2 => x59_out_28,
   I3 => W_45_11_i_12_n_0,
   I4 => W_45_11_i_13_n_0,
   O => W_45_11_i_3_n_0
);
W_45_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x59_out_18,
   I1 => x59_out_25,
   I2 => x59_out_27,
   I3 => W_45_11_i_14_n_0,
   I4 => W_45_11_i_15_n_0,
   O => W_45_11_i_4_n_0
);
W_45_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x59_out_17,
   I1 => x59_out_24,
   I2 => x59_out_26,
   I3 => W_45_11_i_16_n_0,
   I4 => W_45_11_i_17_n_0,
   O => W_45_11_i_5_n_0
);
W_45_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_45_11_i_2_n_0,
   I1 => W_45_15_i_16_n_0,
   I2 => x59_out_21,
   I3 => x59_out_28,
   I4 => x59_out_30,
   I5 => W_45_15_i_17_n_0,
   O => W_45_11_i_6_n_0
);
W_45_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_45_11_i_3_n_0,
   I1 => W_45_11_i_10_n_0,
   I2 => x59_out_20,
   I3 => x59_out_27,
   I4 => x59_out_29,
   I5 => W_45_11_i_11_n_0,
   O => W_45_11_i_7_n_0
);
W_45_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_45_11_i_4_n_0,
   I1 => W_45_11_i_12_n_0,
   I2 => x59_out_19,
   I3 => x59_out_26,
   I4 => x59_out_28,
   I5 => W_45_11_i_13_n_0,
   O => W_45_11_i_8_n_0
);
W_45_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_45_11_i_5_n_0,
   I1 => W_45_11_i_14_n_0,
   I2 => x59_out_18,
   I3 => x59_out_25,
   I4 => x59_out_27,
   I5 => W_45_11_i_15_n_0,
   O => W_45_11_i_9_n_0
);
W_45_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x98_out_14,
   I1 => x74_out_14,
   I2 => x96_out_0,
   I3 => x96_out_21,
   I4 => x96_out_17,
   O => W_45_15_i_10_n_0
);
W_45_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x74_out_13,
   I1 => x96_out_16,
   I2 => x96_out_20,
   I3 => x96_out_31,
   I4 => x98_out_13,
   O => W_45_15_i_11_n_0
);
W_45_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x98_out_13,
   I1 => x74_out_13,
   I2 => x96_out_31,
   I3 => x96_out_20,
   I4 => x96_out_16,
   O => W_45_15_i_12_n_0
);
W_45_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x74_out_12,
   I1 => x96_out_15,
   I2 => x96_out_19,
   I3 => x96_out_30,
   I4 => x98_out_12,
   O => W_45_15_i_13_n_0
);
W_45_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x98_out_12,
   I1 => x74_out_12,
   I2 => x96_out_30,
   I3 => x96_out_19,
   I4 => x96_out_15,
   O => W_45_15_i_14_n_0
);
W_45_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x74_out_11,
   I1 => x96_out_14,
   I2 => x96_out_18,
   I3 => x96_out_29,
   I4 => x98_out_11,
   O => W_45_15_i_15_n_0
);
W_45_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x98_out_11,
   I1 => x74_out_11,
   I2 => x96_out_29,
   I3 => x96_out_18,
   I4 => x96_out_14,
   O => W_45_15_i_16_n_0
);
W_45_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x74_out_10,
   I1 => x96_out_13,
   I2 => x96_out_17,
   I3 => x96_out_28,
   I4 => x98_out_10,
   O => W_45_15_i_17_n_0
);
W_45_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x59_out_24,
   I1 => x59_out_31,
   I2 => x59_out_1,
   I3 => W_45_15_i_10_n_0,
   I4 => W_45_15_i_11_n_0,
   O => W_45_15_i_2_n_0
);
W_45_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x59_out_23,
   I1 => x59_out_30,
   I2 => x59_out_0,
   I3 => W_45_15_i_12_n_0,
   I4 => W_45_15_i_13_n_0,
   O => W_45_15_i_3_n_0
);
W_45_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x59_out_22,
   I1 => x59_out_29,
   I2 => x59_out_31,
   I3 => W_45_15_i_14_n_0,
   I4 => W_45_15_i_15_n_0,
   O => W_45_15_i_4_n_0
);
W_45_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x59_out_21,
   I1 => x59_out_28,
   I2 => x59_out_30,
   I3 => W_45_15_i_16_n_0,
   I4 => W_45_15_i_17_n_0,
   O => W_45_15_i_5_n_0
);
W_45_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_45_15_i_2_n_0,
   I1 => W_45_19_i_16_n_0,
   I2 => x59_out_25,
   I3 => x59_out_0,
   I4 => x59_out_2,
   I5 => W_45_19_i_17_n_0,
   O => W_45_15_i_6_n_0
);
W_45_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_45_15_i_3_n_0,
   I1 => W_45_15_i_10_n_0,
   I2 => x59_out_24,
   I3 => x59_out_31,
   I4 => x59_out_1,
   I5 => W_45_15_i_11_n_0,
   O => W_45_15_i_7_n_0
);
W_45_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_45_15_i_4_n_0,
   I1 => W_45_15_i_12_n_0,
   I2 => x59_out_23,
   I3 => x59_out_30,
   I4 => x59_out_0,
   I5 => W_45_15_i_13_n_0,
   O => W_45_15_i_8_n_0
);
W_45_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_45_15_i_5_n_0,
   I1 => W_45_15_i_14_n_0,
   I2 => x59_out_22,
   I3 => x59_out_29,
   I4 => x59_out_31,
   I5 => W_45_15_i_15_n_0,
   O => W_45_15_i_9_n_0
);
W_45_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x98_out_18,
   I1 => x74_out_18,
   I2 => x96_out_4,
   I3 => x96_out_25,
   I4 => x96_out_21,
   O => W_45_19_i_10_n_0
);
W_45_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x74_out_17,
   I1 => x96_out_20,
   I2 => x96_out_24,
   I3 => x96_out_3,
   I4 => x98_out_17,
   O => W_45_19_i_11_n_0
);
W_45_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x98_out_17,
   I1 => x74_out_17,
   I2 => x96_out_3,
   I3 => x96_out_24,
   I4 => x96_out_20,
   O => W_45_19_i_12_n_0
);
W_45_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x74_out_16,
   I1 => x96_out_19,
   I2 => x96_out_23,
   I3 => x96_out_2,
   I4 => x98_out_16,
   O => W_45_19_i_13_n_0
);
W_45_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x98_out_16,
   I1 => x74_out_16,
   I2 => x96_out_2,
   I3 => x96_out_23,
   I4 => x96_out_19,
   O => W_45_19_i_14_n_0
);
W_45_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x74_out_15,
   I1 => x96_out_18,
   I2 => x96_out_22,
   I3 => x96_out_1,
   I4 => x98_out_15,
   O => W_45_19_i_15_n_0
);
W_45_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x98_out_15,
   I1 => x74_out_15,
   I2 => x96_out_1,
   I3 => x96_out_22,
   I4 => x96_out_18,
   O => W_45_19_i_16_n_0
);
W_45_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x74_out_14,
   I1 => x96_out_17,
   I2 => x96_out_21,
   I3 => x96_out_0,
   I4 => x98_out_14,
   O => W_45_19_i_17_n_0
);
W_45_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x59_out_28,
   I1 => x59_out_3,
   I2 => x59_out_5,
   I3 => W_45_19_i_10_n_0,
   I4 => W_45_19_i_11_n_0,
   O => W_45_19_i_2_n_0
);
W_45_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x59_out_27,
   I1 => x59_out_2,
   I2 => x59_out_4,
   I3 => W_45_19_i_12_n_0,
   I4 => W_45_19_i_13_n_0,
   O => W_45_19_i_3_n_0
);
W_45_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x59_out_26,
   I1 => x59_out_1,
   I2 => x59_out_3,
   I3 => W_45_19_i_14_n_0,
   I4 => W_45_19_i_15_n_0,
   O => W_45_19_i_4_n_0
);
W_45_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x59_out_25,
   I1 => x59_out_0,
   I2 => x59_out_2,
   I3 => W_45_19_i_16_n_0,
   I4 => W_45_19_i_17_n_0,
   O => W_45_19_i_5_n_0
);
W_45_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_45_19_i_2_n_0,
   I1 => W_45_23_i_16_n_0,
   I2 => x59_out_29,
   I3 => x59_out_4,
   I4 => x59_out_6,
   I5 => W_45_23_i_17_n_0,
   O => W_45_19_i_6_n_0
);
W_45_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_45_19_i_3_n_0,
   I1 => W_45_19_i_10_n_0,
   I2 => x59_out_28,
   I3 => x59_out_3,
   I4 => x59_out_5,
   I5 => W_45_19_i_11_n_0,
   O => W_45_19_i_7_n_0
);
W_45_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_45_19_i_4_n_0,
   I1 => W_45_19_i_12_n_0,
   I2 => x59_out_27,
   I3 => x59_out_2,
   I4 => x59_out_4,
   I5 => W_45_19_i_13_n_0,
   O => W_45_19_i_8_n_0
);
W_45_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_45_19_i_5_n_0,
   I1 => W_45_19_i_14_n_0,
   I2 => x59_out_26,
   I3 => x59_out_1,
   I4 => x59_out_3,
   I5 => W_45_19_i_15_n_0,
   O => W_45_19_i_9_n_0
);
W_45_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x98_out_22,
   I1 => x74_out_22,
   I2 => x96_out_8,
   I3 => x96_out_29,
   I4 => x96_out_25,
   O => W_45_23_i_10_n_0
);
W_45_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x74_out_21,
   I1 => x96_out_24,
   I2 => x96_out_28,
   I3 => x96_out_7,
   I4 => x98_out_21,
   O => W_45_23_i_11_n_0
);
W_45_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x98_out_21,
   I1 => x74_out_21,
   I2 => x96_out_7,
   I3 => x96_out_28,
   I4 => x96_out_24,
   O => W_45_23_i_12_n_0
);
W_45_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x74_out_20,
   I1 => x96_out_23,
   I2 => x96_out_27,
   I3 => x96_out_6,
   I4 => x98_out_20,
   O => W_45_23_i_13_n_0
);
W_45_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x98_out_20,
   I1 => x74_out_20,
   I2 => x96_out_6,
   I3 => x96_out_27,
   I4 => x96_out_23,
   O => W_45_23_i_14_n_0
);
W_45_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x74_out_19,
   I1 => x96_out_22,
   I2 => x96_out_26,
   I3 => x96_out_5,
   I4 => x98_out_19,
   O => W_45_23_i_15_n_0
);
W_45_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x98_out_19,
   I1 => x74_out_19,
   I2 => x96_out_5,
   I3 => x96_out_26,
   I4 => x96_out_22,
   O => W_45_23_i_16_n_0
);
W_45_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x74_out_18,
   I1 => x96_out_21,
   I2 => x96_out_25,
   I3 => x96_out_4,
   I4 => x98_out_18,
   O => W_45_23_i_17_n_0
);
W_45_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x59_out_7,
   I1 => x59_out_9,
   I2 => W_45_23_i_10_n_0,
   I3 => W_45_23_i_11_n_0,
   O => W_45_23_i_2_n_0
);
W_45_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x59_out_31,
   I1 => x59_out_6,
   I2 => x59_out_8,
   I3 => W_45_23_i_12_n_0,
   I4 => W_45_23_i_13_n_0,
   O => W_45_23_i_3_n_0
);
W_45_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x59_out_30,
   I1 => x59_out_5,
   I2 => x59_out_7,
   I3 => W_45_23_i_14_n_0,
   I4 => W_45_23_i_15_n_0,
   O => W_45_23_i_4_n_0
);
W_45_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x59_out_29,
   I1 => x59_out_4,
   I2 => x59_out_6,
   I3 => W_45_23_i_16_n_0,
   I4 => W_45_23_i_17_n_0,
   O => W_45_23_i_5_n_0
);
W_45_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x59_out_8,
   I1 => x59_out_10,
   I2 => W_45_27_i_16_n_0,
   I3 => W_45_27_i_17_n_0,
   I4 => W_45_23_i_2_n_0,
   O => W_45_23_i_6_n_0
);
W_45_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x59_out_7,
   I1 => x59_out_9,
   I2 => W_45_23_i_10_n_0,
   I3 => W_45_23_i_11_n_0,
   I4 => W_45_23_i_3_n_0,
   O => W_45_23_i_7_n_0
);
W_45_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_45_23_i_4_n_0,
   I1 => W_45_23_i_12_n_0,
   I2 => x59_out_31,
   I3 => x59_out_6,
   I4 => x59_out_8,
   I5 => W_45_23_i_13_n_0,
   O => W_45_23_i_8_n_0
);
W_45_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_45_23_i_5_n_0,
   I1 => W_45_23_i_14_n_0,
   I2 => x59_out_30,
   I3 => x59_out_5,
   I4 => x59_out_7,
   I5 => W_45_23_i_15_n_0,
   O => W_45_23_i_9_n_0
);
W_45_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x98_out_26,
   I1 => x74_out_26,
   I2 => x96_out_12,
   I3 => x96_out_1,
   I4 => x96_out_29,
   O => W_45_27_i_10_n_0
);
W_45_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x74_out_25,
   I1 => x96_out_28,
   I2 => x96_out_0,
   I3 => x96_out_11,
   I4 => x98_out_25,
   O => W_45_27_i_11_n_0
);
W_45_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x98_out_25,
   I1 => x74_out_25,
   I2 => x96_out_11,
   I3 => x96_out_0,
   I4 => x96_out_28,
   O => W_45_27_i_12_n_0
);
W_45_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x74_out_24,
   I1 => x96_out_27,
   I2 => x96_out_31,
   I3 => x96_out_10,
   I4 => x98_out_24,
   O => W_45_27_i_13_n_0
);
W_45_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x98_out_24,
   I1 => x74_out_24,
   I2 => x96_out_10,
   I3 => x96_out_31,
   I4 => x96_out_27,
   O => W_45_27_i_14_n_0
);
W_45_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x74_out_23,
   I1 => x96_out_26,
   I2 => x96_out_30,
   I3 => x96_out_9,
   I4 => x98_out_23,
   O => W_45_27_i_15_n_0
);
W_45_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x98_out_23,
   I1 => x74_out_23,
   I2 => x96_out_9,
   I3 => x96_out_30,
   I4 => x96_out_26,
   O => W_45_27_i_16_n_0
);
W_45_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x74_out_22,
   I1 => x96_out_25,
   I2 => x96_out_29,
   I3 => x96_out_8,
   I4 => x98_out_22,
   O => W_45_27_i_17_n_0
);
W_45_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x59_out_11,
   I1 => x59_out_13,
   I2 => W_45_27_i_10_n_0,
   I3 => W_45_27_i_11_n_0,
   O => W_45_27_i_2_n_0
);
W_45_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x59_out_10,
   I1 => x59_out_12,
   I2 => W_45_27_i_12_n_0,
   I3 => W_45_27_i_13_n_0,
   O => W_45_27_i_3_n_0
);
W_45_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x59_out_9,
   I1 => x59_out_11,
   I2 => W_45_27_i_14_n_0,
   I3 => W_45_27_i_15_n_0,
   O => W_45_27_i_4_n_0
);
W_45_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x59_out_8,
   I1 => x59_out_10,
   I2 => W_45_27_i_16_n_0,
   I3 => W_45_27_i_17_n_0,
   O => W_45_27_i_5_n_0
);
W_45_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x59_out_12,
   I1 => x59_out_14,
   I2 => W_45_31_i_13_n_0,
   I3 => W_45_31_i_14_n_0,
   I4 => W_45_27_i_2_n_0,
   O => W_45_27_i_6_n_0
);
W_45_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x59_out_11,
   I1 => x59_out_13,
   I2 => W_45_27_i_10_n_0,
   I3 => W_45_27_i_11_n_0,
   I4 => W_45_27_i_3_n_0,
   O => W_45_27_i_7_n_0
);
W_45_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x59_out_10,
   I1 => x59_out_12,
   I2 => W_45_27_i_12_n_0,
   I3 => W_45_27_i_13_n_0,
   I4 => W_45_27_i_4_n_0,
   O => W_45_27_i_8_n_0
);
W_45_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x59_out_9,
   I1 => x59_out_11,
   I2 => W_45_27_i_14_n_0,
   I3 => W_45_27_i_15_n_0,
   I4 => W_45_27_i_5_n_0,
   O => W_45_27_i_9_n_0
);
W_45_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x74_out_28,
   I1 => x96_out_31,
   I2 => x96_out_3,
   I3 => x96_out_14,
   I4 => x98_out_28,
   O => W_45_31_i_10_n_0
);
W_45_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x98_out_28,
   I1 => x74_out_28,
   I2 => x96_out_14,
   I3 => x96_out_3,
   I4 => x96_out_31,
   O => W_45_31_i_11_n_0
);
W_45_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x74_out_27,
   I1 => x96_out_30,
   I2 => x96_out_2,
   I3 => x96_out_13,
   I4 => x98_out_27,
   O => W_45_31_i_12_n_0
);
W_45_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x98_out_27,
   I1 => x74_out_27,
   I2 => x96_out_13,
   I3 => x96_out_2,
   I4 => x96_out_30,
   O => W_45_31_i_13_n_0
);
W_45_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x74_out_26,
   I1 => x96_out_29,
   I2 => x96_out_1,
   I3 => x96_out_12,
   I4 => x98_out_26,
   O => W_45_31_i_14_n_0
);
W_45_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x74_out_29,
   I1 => x96_out_4,
   I2 => x96_out_15,
   I3 => x98_out_29,
   O => W_45_31_i_15_n_0
);
W_45_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x59_out_17,
   I1 => x59_out_15,
   O => SIGMA_LCASE_1155_out_0_30
);
W_45_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => x96_out_6,
   I1 => x96_out_17,
   I2 => x74_out_31,
   I3 => x98_out_31,
   I4 => x59_out_16,
   I5 => x59_out_18,
   O => W_45_31_i_17_n_0
);
W_45_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x96_out_16,
   I1 => x96_out_5,
   O => SIGMA_LCASE_0151_out_30
);
W_45_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x98_out_30,
   I1 => x74_out_30,
   I2 => x96_out_16,
   I3 => x96_out_5,
   O => W_45_31_i_19_n_0
);
W_45_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x59_out_14,
   I1 => x59_out_16,
   I2 => W_45_31_i_9_n_0,
   I3 => W_45_31_i_10_n_0,
   O => W_45_31_i_2_n_0
);
W_45_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x59_out_13,
   I1 => x59_out_15,
   I2 => W_45_31_i_11_n_0,
   I3 => W_45_31_i_12_n_0,
   O => W_45_31_i_3_n_0
);
W_45_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x59_out_12,
   I1 => x59_out_14,
   I2 => W_45_31_i_13_n_0,
   I3 => W_45_31_i_14_n_0,
   O => W_45_31_i_4_n_0
);
W_45_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_45_31_i_15_n_0,
   I1 => SIGMA_LCASE_1155_out_0_30,
   I2 => W_45_31_i_17_n_0,
   I3 => x74_out_30,
   I4 => SIGMA_LCASE_0151_out_30,
   I5 => x98_out_30,
   O => W_45_31_i_5_n_0
);
W_45_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_45_31_i_2_n_0,
   I1 => W_45_31_i_19_n_0,
   I2 => x59_out_15,
   I3 => x59_out_17,
   I4 => W_45_31_i_15_n_0,
   O => W_45_31_i_6_n_0
);
W_45_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x59_out_14,
   I1 => x59_out_16,
   I2 => W_45_31_i_9_n_0,
   I3 => W_45_31_i_10_n_0,
   I4 => W_45_31_i_3_n_0,
   O => W_45_31_i_7_n_0
);
W_45_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x59_out_13,
   I1 => x59_out_15,
   I2 => W_45_31_i_11_n_0,
   I3 => W_45_31_i_12_n_0,
   I4 => W_45_31_i_4_n_0,
   O => W_45_31_i_8_n_0
);
W_45_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x98_out_29,
   I1 => x74_out_29,
   I2 => x96_out_15,
   I3 => x96_out_4,
   O => W_45_31_i_9_n_0
);
W_45_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x98_out_2,
   I1 => x74_out_2,
   I2 => x96_out_20,
   I3 => x96_out_9,
   I4 => x96_out_5,
   O => W_45_3_i_10_n_0
);
W_45_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x74_out_1,
   I1 => x96_out_4,
   I2 => x96_out_8,
   I3 => x96_out_19,
   I4 => x98_out_1,
   O => W_45_3_i_11_n_0
);
W_45_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x96_out_19,
   I1 => x96_out_8,
   I2 => x96_out_4,
   O => SIGMA_LCASE_0151_out_1
);
W_45_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x59_out_21,
   I1 => x59_out_19,
   I2 => x59_out_12,
   O => SIGMA_LCASE_1155_out_0_2
);
W_45_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x59_out_20,
   I1 => x59_out_18,
   I2 => x59_out_11,
   O => SIGMA_LCASE_1155_out_1
);
W_45_3_i_15 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x98_out_1,
   I1 => x74_out_1,
   I2 => x96_out_19,
   I3 => x96_out_8,
   I4 => x96_out_4,
   O => W_45_3_i_15_n_0
);
W_45_3_i_16 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x96_out_18,
   I1 => x96_out_7,
   I2 => x96_out_3,
   O => SIGMA_LCASE_0151_out_0
);
W_45_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x59_out_12,
   I1 => x59_out_19,
   I2 => x59_out_21,
   I3 => W_45_3_i_10_n_0,
   I4 => W_45_3_i_11_n_0,
   O => W_45_3_i_2_n_0
);
W_45_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_45_3_i_11_n_0,
   I1 => x59_out_21,
   I2 => x59_out_19,
   I3 => x59_out_12,
   I4 => W_45_3_i_10_n_0,
   O => W_45_3_i_3_n_0
);
W_45_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_0151_out_1,
   I1 => x74_out_1,
   I2 => x98_out_1,
   I3 => x59_out_11,
   I4 => x59_out_18,
   I5 => x59_out_20,
   O => W_45_3_i_4_n_0
);
W_45_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x98_out_0,
   I1 => x74_out_0,
   I2 => x96_out_18,
   I3 => x96_out_7,
   I4 => x96_out_3,
   O => W_45_3_i_5_n_0
);
W_45_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_45_3_i_2_n_0,
   I1 => W_45_7_i_16_n_0,
   I2 => x59_out_13,
   I3 => x59_out_20,
   I4 => x59_out_22,
   I5 => W_45_7_i_17_n_0,
   O => W_45_3_i_6_n_0
);
W_45_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_45_3_i_10_n_0,
   I1 => SIGMA_LCASE_1155_out_0_2,
   I2 => x98_out_1,
   I3 => x74_out_1,
   I4 => SIGMA_LCASE_0151_out_1,
   I5 => SIGMA_LCASE_1155_out_1,
   O => W_45_3_i_7_n_0
);
W_45_3_i_8 : LUT5
  generic map(
   INIT => X"99969666"
  )
 port map (
   I0 => SIGMA_LCASE_1155_out_1,
   I1 => W_45_3_i_15_n_0,
   I2 => x98_out_0,
   I3 => SIGMA_LCASE_0151_out_0,
   I4 => x74_out_0,
   O => W_45_3_i_8_n_0
);
W_45_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_45_3_i_5_n_0,
   I1 => x59_out_10,
   I2 => x59_out_17,
   I3 => x59_out_19,
   O => W_45_3_i_9_n_0
);
W_45_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x98_out_6,
   I1 => x74_out_6,
   I2 => x96_out_24,
   I3 => x96_out_13,
   I4 => x96_out_9,
   O => W_45_7_i_10_n_0
);
W_45_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x74_out_5,
   I1 => x96_out_8,
   I2 => x96_out_12,
   I3 => x96_out_23,
   I4 => x98_out_5,
   O => W_45_7_i_11_n_0
);
W_45_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x98_out_5,
   I1 => x74_out_5,
   I2 => x96_out_23,
   I3 => x96_out_12,
   I4 => x96_out_8,
   O => W_45_7_i_12_n_0
);
W_45_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x74_out_4,
   I1 => x96_out_7,
   I2 => x96_out_11,
   I3 => x96_out_22,
   I4 => x98_out_4,
   O => W_45_7_i_13_n_0
);
W_45_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x98_out_4,
   I1 => x74_out_4,
   I2 => x96_out_22,
   I3 => x96_out_11,
   I4 => x96_out_7,
   O => W_45_7_i_14_n_0
);
W_45_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x74_out_3,
   I1 => x96_out_6,
   I2 => x96_out_10,
   I3 => x96_out_21,
   I4 => x98_out_3,
   O => W_45_7_i_15_n_0
);
W_45_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x98_out_3,
   I1 => x74_out_3,
   I2 => x96_out_21,
   I3 => x96_out_10,
   I4 => x96_out_6,
   O => W_45_7_i_16_n_0
);
W_45_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x74_out_2,
   I1 => x96_out_5,
   I2 => x96_out_9,
   I3 => x96_out_20,
   I4 => x98_out_2,
   O => W_45_7_i_17_n_0
);
W_45_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x59_out_16,
   I1 => x59_out_23,
   I2 => x59_out_25,
   I3 => W_45_7_i_10_n_0,
   I4 => W_45_7_i_11_n_0,
   O => W_45_7_i_2_n_0
);
W_45_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x59_out_15,
   I1 => x59_out_22,
   I2 => x59_out_24,
   I3 => W_45_7_i_12_n_0,
   I4 => W_45_7_i_13_n_0,
   O => W_45_7_i_3_n_0
);
W_45_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x59_out_14,
   I1 => x59_out_21,
   I2 => x59_out_23,
   I3 => W_45_7_i_14_n_0,
   I4 => W_45_7_i_15_n_0,
   O => W_45_7_i_4_n_0
);
W_45_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x59_out_13,
   I1 => x59_out_20,
   I2 => x59_out_22,
   I3 => W_45_7_i_16_n_0,
   I4 => W_45_7_i_17_n_0,
   O => W_45_7_i_5_n_0
);
W_45_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_45_7_i_2_n_0,
   I1 => W_45_11_i_16_n_0,
   I2 => x59_out_17,
   I3 => x59_out_24,
   I4 => x59_out_26,
   I5 => W_45_11_i_17_n_0,
   O => W_45_7_i_6_n_0
);
W_45_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_45_7_i_3_n_0,
   I1 => W_45_7_i_10_n_0,
   I2 => x59_out_16,
   I3 => x59_out_23,
   I4 => x59_out_25,
   I5 => W_45_7_i_11_n_0,
   O => W_45_7_i_7_n_0
);
W_45_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_45_7_i_4_n_0,
   I1 => W_45_7_i_12_n_0,
   I2 => x59_out_15,
   I3 => x59_out_22,
   I4 => x59_out_24,
   I5 => W_45_7_i_13_n_0,
   O => W_45_7_i_8_n_0
);
W_45_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_45_7_i_5_n_0,
   I1 => W_45_7_i_14_n_0,
   I2 => x59_out_14,
   I3 => x59_out_21,
   I4 => x59_out_23,
   I5 => W_45_7_i_15_n_0,
   O => W_45_7_i_9_n_0
);
W_46_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x96_out_10,
   I1 => x71_out_10,
   I2 => x94_out_28,
   I3 => x94_out_17,
   I4 => x94_out_13,
   O => W_46_11_i_10_n_0
);
W_46_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x71_out_9,
   I1 => x94_out_12,
   I2 => x94_out_16,
   I3 => x94_out_27,
   I4 => x96_out_9,
   O => W_46_11_i_11_n_0
);
W_46_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x96_out_9,
   I1 => x71_out_9,
   I2 => x94_out_27,
   I3 => x94_out_16,
   I4 => x94_out_12,
   O => W_46_11_i_12_n_0
);
W_46_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x71_out_8,
   I1 => x94_out_11,
   I2 => x94_out_15,
   I3 => x94_out_26,
   I4 => x96_out_8,
   O => W_46_11_i_13_n_0
);
W_46_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x96_out_8,
   I1 => x71_out_8,
   I2 => x94_out_26,
   I3 => x94_out_15,
   I4 => x94_out_11,
   O => W_46_11_i_14_n_0
);
W_46_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x71_out_7,
   I1 => x94_out_10,
   I2 => x94_out_14,
   I3 => x94_out_25,
   I4 => x96_out_7,
   O => W_46_11_i_15_n_0
);
W_46_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x96_out_7,
   I1 => x71_out_7,
   I2 => x94_out_25,
   I3 => x94_out_14,
   I4 => x94_out_10,
   O => W_46_11_i_16_n_0
);
W_46_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x71_out_6,
   I1 => x94_out_9,
   I2 => x94_out_13,
   I3 => x94_out_24,
   I4 => x96_out_6,
   O => W_46_11_i_17_n_0
);
W_46_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x56_out_20,
   I1 => x56_out_27,
   I2 => x56_out_29,
   I3 => W_46_11_i_10_n_0,
   I4 => W_46_11_i_11_n_0,
   O => W_46_11_i_2_n_0
);
W_46_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x56_out_19,
   I1 => x56_out_26,
   I2 => x56_out_28,
   I3 => W_46_11_i_12_n_0,
   I4 => W_46_11_i_13_n_0,
   O => W_46_11_i_3_n_0
);
W_46_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x56_out_18,
   I1 => x56_out_25,
   I2 => x56_out_27,
   I3 => W_46_11_i_14_n_0,
   I4 => W_46_11_i_15_n_0,
   O => W_46_11_i_4_n_0
);
W_46_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x56_out_17,
   I1 => x56_out_24,
   I2 => x56_out_26,
   I3 => W_46_11_i_16_n_0,
   I4 => W_46_11_i_17_n_0,
   O => W_46_11_i_5_n_0
);
W_46_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_46_11_i_2_n_0,
   I1 => W_46_15_i_16_n_0,
   I2 => x56_out_21,
   I3 => x56_out_28,
   I4 => x56_out_30,
   I5 => W_46_15_i_17_n_0,
   O => W_46_11_i_6_n_0
);
W_46_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_46_11_i_3_n_0,
   I1 => W_46_11_i_10_n_0,
   I2 => x56_out_20,
   I3 => x56_out_27,
   I4 => x56_out_29,
   I5 => W_46_11_i_11_n_0,
   O => W_46_11_i_7_n_0
);
W_46_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_46_11_i_4_n_0,
   I1 => W_46_11_i_12_n_0,
   I2 => x56_out_19,
   I3 => x56_out_26,
   I4 => x56_out_28,
   I5 => W_46_11_i_13_n_0,
   O => W_46_11_i_8_n_0
);
W_46_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_46_11_i_5_n_0,
   I1 => W_46_11_i_14_n_0,
   I2 => x56_out_18,
   I3 => x56_out_25,
   I4 => x56_out_27,
   I5 => W_46_11_i_15_n_0,
   O => W_46_11_i_9_n_0
);
W_46_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x96_out_14,
   I1 => x71_out_14,
   I2 => x94_out_0,
   I3 => x94_out_21,
   I4 => x94_out_17,
   O => W_46_15_i_10_n_0
);
W_46_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x71_out_13,
   I1 => x94_out_16,
   I2 => x94_out_20,
   I3 => x94_out_31,
   I4 => x96_out_13,
   O => W_46_15_i_11_n_0
);
W_46_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x96_out_13,
   I1 => x71_out_13,
   I2 => x94_out_31,
   I3 => x94_out_20,
   I4 => x94_out_16,
   O => W_46_15_i_12_n_0
);
W_46_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x71_out_12,
   I1 => x94_out_15,
   I2 => x94_out_19,
   I3 => x94_out_30,
   I4 => x96_out_12,
   O => W_46_15_i_13_n_0
);
W_46_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x96_out_12,
   I1 => x71_out_12,
   I2 => x94_out_30,
   I3 => x94_out_19,
   I4 => x94_out_15,
   O => W_46_15_i_14_n_0
);
W_46_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x71_out_11,
   I1 => x94_out_14,
   I2 => x94_out_18,
   I3 => x94_out_29,
   I4 => x96_out_11,
   O => W_46_15_i_15_n_0
);
W_46_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x96_out_11,
   I1 => x71_out_11,
   I2 => x94_out_29,
   I3 => x94_out_18,
   I4 => x94_out_14,
   O => W_46_15_i_16_n_0
);
W_46_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x71_out_10,
   I1 => x94_out_13,
   I2 => x94_out_17,
   I3 => x94_out_28,
   I4 => x96_out_10,
   O => W_46_15_i_17_n_0
);
W_46_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x56_out_24,
   I1 => x56_out_31,
   I2 => x56_out_1,
   I3 => W_46_15_i_10_n_0,
   I4 => W_46_15_i_11_n_0,
   O => W_46_15_i_2_n_0
);
W_46_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x56_out_23,
   I1 => x56_out_30,
   I2 => x56_out_0,
   I3 => W_46_15_i_12_n_0,
   I4 => W_46_15_i_13_n_0,
   O => W_46_15_i_3_n_0
);
W_46_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x56_out_22,
   I1 => x56_out_29,
   I2 => x56_out_31,
   I3 => W_46_15_i_14_n_0,
   I4 => W_46_15_i_15_n_0,
   O => W_46_15_i_4_n_0
);
W_46_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x56_out_21,
   I1 => x56_out_28,
   I2 => x56_out_30,
   I3 => W_46_15_i_16_n_0,
   I4 => W_46_15_i_17_n_0,
   O => W_46_15_i_5_n_0
);
W_46_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_46_15_i_2_n_0,
   I1 => W_46_19_i_16_n_0,
   I2 => x56_out_25,
   I3 => x56_out_0,
   I4 => x56_out_2,
   I5 => W_46_19_i_17_n_0,
   O => W_46_15_i_6_n_0
);
W_46_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_46_15_i_3_n_0,
   I1 => W_46_15_i_10_n_0,
   I2 => x56_out_24,
   I3 => x56_out_31,
   I4 => x56_out_1,
   I5 => W_46_15_i_11_n_0,
   O => W_46_15_i_7_n_0
);
W_46_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_46_15_i_4_n_0,
   I1 => W_46_15_i_12_n_0,
   I2 => x56_out_23,
   I3 => x56_out_30,
   I4 => x56_out_0,
   I5 => W_46_15_i_13_n_0,
   O => W_46_15_i_8_n_0
);
W_46_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_46_15_i_5_n_0,
   I1 => W_46_15_i_14_n_0,
   I2 => x56_out_22,
   I3 => x56_out_29,
   I4 => x56_out_31,
   I5 => W_46_15_i_15_n_0,
   O => W_46_15_i_9_n_0
);
W_46_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x96_out_18,
   I1 => x71_out_18,
   I2 => x94_out_4,
   I3 => x94_out_25,
   I4 => x94_out_21,
   O => W_46_19_i_10_n_0
);
W_46_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x71_out_17,
   I1 => x94_out_20,
   I2 => x94_out_24,
   I3 => x94_out_3,
   I4 => x96_out_17,
   O => W_46_19_i_11_n_0
);
W_46_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x96_out_17,
   I1 => x71_out_17,
   I2 => x94_out_3,
   I3 => x94_out_24,
   I4 => x94_out_20,
   O => W_46_19_i_12_n_0
);
W_46_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x71_out_16,
   I1 => x94_out_19,
   I2 => x94_out_23,
   I3 => x94_out_2,
   I4 => x96_out_16,
   O => W_46_19_i_13_n_0
);
W_46_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x96_out_16,
   I1 => x71_out_16,
   I2 => x94_out_2,
   I3 => x94_out_23,
   I4 => x94_out_19,
   O => W_46_19_i_14_n_0
);
W_46_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x71_out_15,
   I1 => x94_out_18,
   I2 => x94_out_22,
   I3 => x94_out_1,
   I4 => x96_out_15,
   O => W_46_19_i_15_n_0
);
W_46_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x96_out_15,
   I1 => x71_out_15,
   I2 => x94_out_1,
   I3 => x94_out_22,
   I4 => x94_out_18,
   O => W_46_19_i_16_n_0
);
W_46_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x71_out_14,
   I1 => x94_out_17,
   I2 => x94_out_21,
   I3 => x94_out_0,
   I4 => x96_out_14,
   O => W_46_19_i_17_n_0
);
W_46_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x56_out_28,
   I1 => x56_out_3,
   I2 => x56_out_5,
   I3 => W_46_19_i_10_n_0,
   I4 => W_46_19_i_11_n_0,
   O => W_46_19_i_2_n_0
);
W_46_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x56_out_27,
   I1 => x56_out_2,
   I2 => x56_out_4,
   I3 => W_46_19_i_12_n_0,
   I4 => W_46_19_i_13_n_0,
   O => W_46_19_i_3_n_0
);
W_46_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x56_out_26,
   I1 => x56_out_1,
   I2 => x56_out_3,
   I3 => W_46_19_i_14_n_0,
   I4 => W_46_19_i_15_n_0,
   O => W_46_19_i_4_n_0
);
W_46_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x56_out_25,
   I1 => x56_out_0,
   I2 => x56_out_2,
   I3 => W_46_19_i_16_n_0,
   I4 => W_46_19_i_17_n_0,
   O => W_46_19_i_5_n_0
);
W_46_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_46_19_i_2_n_0,
   I1 => W_46_23_i_16_n_0,
   I2 => x56_out_29,
   I3 => x56_out_4,
   I4 => x56_out_6,
   I5 => W_46_23_i_17_n_0,
   O => W_46_19_i_6_n_0
);
W_46_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_46_19_i_3_n_0,
   I1 => W_46_19_i_10_n_0,
   I2 => x56_out_28,
   I3 => x56_out_3,
   I4 => x56_out_5,
   I5 => W_46_19_i_11_n_0,
   O => W_46_19_i_7_n_0
);
W_46_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_46_19_i_4_n_0,
   I1 => W_46_19_i_12_n_0,
   I2 => x56_out_27,
   I3 => x56_out_2,
   I4 => x56_out_4,
   I5 => W_46_19_i_13_n_0,
   O => W_46_19_i_8_n_0
);
W_46_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_46_19_i_5_n_0,
   I1 => W_46_19_i_14_n_0,
   I2 => x56_out_26,
   I3 => x56_out_1,
   I4 => x56_out_3,
   I5 => W_46_19_i_15_n_0,
   O => W_46_19_i_9_n_0
);
W_46_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x96_out_22,
   I1 => x71_out_22,
   I2 => x94_out_8,
   I3 => x94_out_29,
   I4 => x94_out_25,
   O => W_46_23_i_10_n_0
);
W_46_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x71_out_21,
   I1 => x94_out_24,
   I2 => x94_out_28,
   I3 => x94_out_7,
   I4 => x96_out_21,
   O => W_46_23_i_11_n_0
);
W_46_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x96_out_21,
   I1 => x71_out_21,
   I2 => x94_out_7,
   I3 => x94_out_28,
   I4 => x94_out_24,
   O => W_46_23_i_12_n_0
);
W_46_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x71_out_20,
   I1 => x94_out_23,
   I2 => x94_out_27,
   I3 => x94_out_6,
   I4 => x96_out_20,
   O => W_46_23_i_13_n_0
);
W_46_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x96_out_20,
   I1 => x71_out_20,
   I2 => x94_out_6,
   I3 => x94_out_27,
   I4 => x94_out_23,
   O => W_46_23_i_14_n_0
);
W_46_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x71_out_19,
   I1 => x94_out_22,
   I2 => x94_out_26,
   I3 => x94_out_5,
   I4 => x96_out_19,
   O => W_46_23_i_15_n_0
);
W_46_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x96_out_19,
   I1 => x71_out_19,
   I2 => x94_out_5,
   I3 => x94_out_26,
   I4 => x94_out_22,
   O => W_46_23_i_16_n_0
);
W_46_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x71_out_18,
   I1 => x94_out_21,
   I2 => x94_out_25,
   I3 => x94_out_4,
   I4 => x96_out_18,
   O => W_46_23_i_17_n_0
);
W_46_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x56_out_7,
   I1 => x56_out_9,
   I2 => W_46_23_i_10_n_0,
   I3 => W_46_23_i_11_n_0,
   O => W_46_23_i_2_n_0
);
W_46_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x56_out_31,
   I1 => x56_out_6,
   I2 => x56_out_8,
   I3 => W_46_23_i_12_n_0,
   I4 => W_46_23_i_13_n_0,
   O => W_46_23_i_3_n_0
);
W_46_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x56_out_30,
   I1 => x56_out_5,
   I2 => x56_out_7,
   I3 => W_46_23_i_14_n_0,
   I4 => W_46_23_i_15_n_0,
   O => W_46_23_i_4_n_0
);
W_46_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x56_out_29,
   I1 => x56_out_4,
   I2 => x56_out_6,
   I3 => W_46_23_i_16_n_0,
   I4 => W_46_23_i_17_n_0,
   O => W_46_23_i_5_n_0
);
W_46_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x56_out_8,
   I1 => x56_out_10,
   I2 => W_46_27_i_16_n_0,
   I3 => W_46_27_i_17_n_0,
   I4 => W_46_23_i_2_n_0,
   O => W_46_23_i_6_n_0
);
W_46_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x56_out_7,
   I1 => x56_out_9,
   I2 => W_46_23_i_10_n_0,
   I3 => W_46_23_i_11_n_0,
   I4 => W_46_23_i_3_n_0,
   O => W_46_23_i_7_n_0
);
W_46_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_46_23_i_4_n_0,
   I1 => W_46_23_i_12_n_0,
   I2 => x56_out_31,
   I3 => x56_out_6,
   I4 => x56_out_8,
   I5 => W_46_23_i_13_n_0,
   O => W_46_23_i_8_n_0
);
W_46_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_46_23_i_5_n_0,
   I1 => W_46_23_i_14_n_0,
   I2 => x56_out_30,
   I3 => x56_out_5,
   I4 => x56_out_7,
   I5 => W_46_23_i_15_n_0,
   O => W_46_23_i_9_n_0
);
W_46_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x96_out_26,
   I1 => x71_out_26,
   I2 => x94_out_12,
   I3 => x94_out_1,
   I4 => x94_out_29,
   O => W_46_27_i_10_n_0
);
W_46_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x71_out_25,
   I1 => x94_out_28,
   I2 => x94_out_0,
   I3 => x94_out_11,
   I4 => x96_out_25,
   O => W_46_27_i_11_n_0
);
W_46_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x96_out_25,
   I1 => x71_out_25,
   I2 => x94_out_11,
   I3 => x94_out_0,
   I4 => x94_out_28,
   O => W_46_27_i_12_n_0
);
W_46_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x71_out_24,
   I1 => x94_out_27,
   I2 => x94_out_31,
   I3 => x94_out_10,
   I4 => x96_out_24,
   O => W_46_27_i_13_n_0
);
W_46_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x96_out_24,
   I1 => x71_out_24,
   I2 => x94_out_10,
   I3 => x94_out_31,
   I4 => x94_out_27,
   O => W_46_27_i_14_n_0
);
W_46_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x71_out_23,
   I1 => x94_out_26,
   I2 => x94_out_30,
   I3 => x94_out_9,
   I4 => x96_out_23,
   O => W_46_27_i_15_n_0
);
W_46_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x96_out_23,
   I1 => x71_out_23,
   I2 => x94_out_9,
   I3 => x94_out_30,
   I4 => x94_out_26,
   O => W_46_27_i_16_n_0
);
W_46_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x71_out_22,
   I1 => x94_out_25,
   I2 => x94_out_29,
   I3 => x94_out_8,
   I4 => x96_out_22,
   O => W_46_27_i_17_n_0
);
W_46_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x56_out_11,
   I1 => x56_out_13,
   I2 => W_46_27_i_10_n_0,
   I3 => W_46_27_i_11_n_0,
   O => W_46_27_i_2_n_0
);
W_46_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x56_out_10,
   I1 => x56_out_12,
   I2 => W_46_27_i_12_n_0,
   I3 => W_46_27_i_13_n_0,
   O => W_46_27_i_3_n_0
);
W_46_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x56_out_9,
   I1 => x56_out_11,
   I2 => W_46_27_i_14_n_0,
   I3 => W_46_27_i_15_n_0,
   O => W_46_27_i_4_n_0
);
W_46_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x56_out_8,
   I1 => x56_out_10,
   I2 => W_46_27_i_16_n_0,
   I3 => W_46_27_i_17_n_0,
   O => W_46_27_i_5_n_0
);
W_46_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x56_out_12,
   I1 => x56_out_14,
   I2 => W_46_31_i_13_n_0,
   I3 => W_46_31_i_14_n_0,
   I4 => W_46_27_i_2_n_0,
   O => W_46_27_i_6_n_0
);
W_46_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x56_out_11,
   I1 => x56_out_13,
   I2 => W_46_27_i_10_n_0,
   I3 => W_46_27_i_11_n_0,
   I4 => W_46_27_i_3_n_0,
   O => W_46_27_i_7_n_0
);
W_46_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x56_out_10,
   I1 => x56_out_12,
   I2 => W_46_27_i_12_n_0,
   I3 => W_46_27_i_13_n_0,
   I4 => W_46_27_i_4_n_0,
   O => W_46_27_i_8_n_0
);
W_46_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x56_out_9,
   I1 => x56_out_11,
   I2 => W_46_27_i_14_n_0,
   I3 => W_46_27_i_15_n_0,
   I4 => W_46_27_i_5_n_0,
   O => W_46_27_i_9_n_0
);
W_46_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x71_out_28,
   I1 => x94_out_31,
   I2 => x94_out_3,
   I3 => x94_out_14,
   I4 => x96_out_28,
   O => W_46_31_i_10_n_0
);
W_46_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x96_out_28,
   I1 => x71_out_28,
   I2 => x94_out_14,
   I3 => x94_out_3,
   I4 => x94_out_31,
   O => W_46_31_i_11_n_0
);
W_46_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x71_out_27,
   I1 => x94_out_30,
   I2 => x94_out_2,
   I3 => x94_out_13,
   I4 => x96_out_27,
   O => W_46_31_i_12_n_0
);
W_46_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x96_out_27,
   I1 => x71_out_27,
   I2 => x94_out_13,
   I3 => x94_out_2,
   I4 => x94_out_30,
   O => W_46_31_i_13_n_0
);
W_46_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x71_out_26,
   I1 => x94_out_29,
   I2 => x94_out_1,
   I3 => x94_out_12,
   I4 => x96_out_26,
   O => W_46_31_i_14_n_0
);
W_46_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x71_out_29,
   I1 => x94_out_4,
   I2 => x94_out_15,
   I3 => x96_out_29,
   O => W_46_31_i_15_n_0
);
W_46_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x56_out_17,
   I1 => x56_out_15,
   O => SIGMA_LCASE_1147_out_0_30
);
W_46_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => x94_out_6,
   I1 => x94_out_17,
   I2 => x71_out_31,
   I3 => x96_out_31,
   I4 => x56_out_16,
   I5 => x56_out_18,
   O => W_46_31_i_17_n_0
);
W_46_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x94_out_16,
   I1 => x94_out_5,
   O => SIGMA_LCASE_0143_out_30
);
W_46_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x96_out_30,
   I1 => x71_out_30,
   I2 => x94_out_16,
   I3 => x94_out_5,
   O => W_46_31_i_19_n_0
);
W_46_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x56_out_14,
   I1 => x56_out_16,
   I2 => W_46_31_i_9_n_0,
   I3 => W_46_31_i_10_n_0,
   O => W_46_31_i_2_n_0
);
W_46_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x56_out_13,
   I1 => x56_out_15,
   I2 => W_46_31_i_11_n_0,
   I3 => W_46_31_i_12_n_0,
   O => W_46_31_i_3_n_0
);
W_46_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x56_out_12,
   I1 => x56_out_14,
   I2 => W_46_31_i_13_n_0,
   I3 => W_46_31_i_14_n_0,
   O => W_46_31_i_4_n_0
);
W_46_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_46_31_i_15_n_0,
   I1 => SIGMA_LCASE_1147_out_0_30,
   I2 => W_46_31_i_17_n_0,
   I3 => x71_out_30,
   I4 => SIGMA_LCASE_0143_out_30,
   I5 => x96_out_30,
   O => W_46_31_i_5_n_0
);
W_46_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_46_31_i_2_n_0,
   I1 => W_46_31_i_19_n_0,
   I2 => x56_out_15,
   I3 => x56_out_17,
   I4 => W_46_31_i_15_n_0,
   O => W_46_31_i_6_n_0
);
W_46_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x56_out_14,
   I1 => x56_out_16,
   I2 => W_46_31_i_9_n_0,
   I3 => W_46_31_i_10_n_0,
   I4 => W_46_31_i_3_n_0,
   O => W_46_31_i_7_n_0
);
W_46_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x56_out_13,
   I1 => x56_out_15,
   I2 => W_46_31_i_11_n_0,
   I3 => W_46_31_i_12_n_0,
   I4 => W_46_31_i_4_n_0,
   O => W_46_31_i_8_n_0
);
W_46_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x96_out_29,
   I1 => x71_out_29,
   I2 => x94_out_15,
   I3 => x94_out_4,
   O => W_46_31_i_9_n_0
);
W_46_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x96_out_2,
   I1 => x71_out_2,
   I2 => x94_out_20,
   I3 => x94_out_9,
   I4 => x94_out_5,
   O => W_46_3_i_10_n_0
);
W_46_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x71_out_1,
   I1 => x94_out_4,
   I2 => x94_out_8,
   I3 => x94_out_19,
   I4 => x96_out_1,
   O => W_46_3_i_11_n_0
);
W_46_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x94_out_19,
   I1 => x94_out_8,
   I2 => x94_out_4,
   O => SIGMA_LCASE_0143_out_1
);
W_46_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x56_out_21,
   I1 => x56_out_19,
   I2 => x56_out_12,
   O => SIGMA_LCASE_1147_out_0_2
);
W_46_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x56_out_20,
   I1 => x56_out_18,
   I2 => x56_out_11,
   O => SIGMA_LCASE_1147_out_1
);
W_46_3_i_15 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x96_out_1,
   I1 => x71_out_1,
   I2 => x94_out_19,
   I3 => x94_out_8,
   I4 => x94_out_4,
   O => W_46_3_i_15_n_0
);
W_46_3_i_16 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x94_out_18,
   I1 => x94_out_7,
   I2 => x94_out_3,
   O => SIGMA_LCASE_0143_out_0
);
W_46_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x56_out_12,
   I1 => x56_out_19,
   I2 => x56_out_21,
   I3 => W_46_3_i_10_n_0,
   I4 => W_46_3_i_11_n_0,
   O => W_46_3_i_2_n_0
);
W_46_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_46_3_i_11_n_0,
   I1 => x56_out_21,
   I2 => x56_out_19,
   I3 => x56_out_12,
   I4 => W_46_3_i_10_n_0,
   O => W_46_3_i_3_n_0
);
W_46_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_0143_out_1,
   I1 => x71_out_1,
   I2 => x96_out_1,
   I3 => x56_out_11,
   I4 => x56_out_18,
   I5 => x56_out_20,
   O => W_46_3_i_4_n_0
);
W_46_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x96_out_0,
   I1 => x71_out_0,
   I2 => x94_out_18,
   I3 => x94_out_7,
   I4 => x94_out_3,
   O => W_46_3_i_5_n_0
);
W_46_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_46_3_i_2_n_0,
   I1 => W_46_7_i_16_n_0,
   I2 => x56_out_13,
   I3 => x56_out_20,
   I4 => x56_out_22,
   I5 => W_46_7_i_17_n_0,
   O => W_46_3_i_6_n_0
);
W_46_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_46_3_i_10_n_0,
   I1 => SIGMA_LCASE_1147_out_0_2,
   I2 => x96_out_1,
   I3 => x71_out_1,
   I4 => SIGMA_LCASE_0143_out_1,
   I5 => SIGMA_LCASE_1147_out_1,
   O => W_46_3_i_7_n_0
);
W_46_3_i_8 : LUT5
  generic map(
   INIT => X"99969666"
  )
 port map (
   I0 => SIGMA_LCASE_1147_out_1,
   I1 => W_46_3_i_15_n_0,
   I2 => x96_out_0,
   I3 => SIGMA_LCASE_0143_out_0,
   I4 => x71_out_0,
   O => W_46_3_i_8_n_0
);
W_46_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_46_3_i_5_n_0,
   I1 => x56_out_10,
   I2 => x56_out_17,
   I3 => x56_out_19,
   O => W_46_3_i_9_n_0
);
W_46_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x96_out_6,
   I1 => x71_out_6,
   I2 => x94_out_24,
   I3 => x94_out_13,
   I4 => x94_out_9,
   O => W_46_7_i_10_n_0
);
W_46_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x71_out_5,
   I1 => x94_out_8,
   I2 => x94_out_12,
   I3 => x94_out_23,
   I4 => x96_out_5,
   O => W_46_7_i_11_n_0
);
W_46_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x96_out_5,
   I1 => x71_out_5,
   I2 => x94_out_23,
   I3 => x94_out_12,
   I4 => x94_out_8,
   O => W_46_7_i_12_n_0
);
W_46_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x71_out_4,
   I1 => x94_out_7,
   I2 => x94_out_11,
   I3 => x94_out_22,
   I4 => x96_out_4,
   O => W_46_7_i_13_n_0
);
W_46_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x96_out_4,
   I1 => x71_out_4,
   I2 => x94_out_22,
   I3 => x94_out_11,
   I4 => x94_out_7,
   O => W_46_7_i_14_n_0
);
W_46_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x71_out_3,
   I1 => x94_out_6,
   I2 => x94_out_10,
   I3 => x94_out_21,
   I4 => x96_out_3,
   O => W_46_7_i_15_n_0
);
W_46_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x96_out_3,
   I1 => x71_out_3,
   I2 => x94_out_21,
   I3 => x94_out_10,
   I4 => x94_out_6,
   O => W_46_7_i_16_n_0
);
W_46_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x71_out_2,
   I1 => x94_out_5,
   I2 => x94_out_9,
   I3 => x94_out_20,
   I4 => x96_out_2,
   O => W_46_7_i_17_n_0
);
W_46_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x56_out_16,
   I1 => x56_out_23,
   I2 => x56_out_25,
   I3 => W_46_7_i_10_n_0,
   I4 => W_46_7_i_11_n_0,
   O => W_46_7_i_2_n_0
);
W_46_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x56_out_15,
   I1 => x56_out_22,
   I2 => x56_out_24,
   I3 => W_46_7_i_12_n_0,
   I4 => W_46_7_i_13_n_0,
   O => W_46_7_i_3_n_0
);
W_46_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x56_out_14,
   I1 => x56_out_21,
   I2 => x56_out_23,
   I3 => W_46_7_i_14_n_0,
   I4 => W_46_7_i_15_n_0,
   O => W_46_7_i_4_n_0
);
W_46_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x56_out_13,
   I1 => x56_out_20,
   I2 => x56_out_22,
   I3 => W_46_7_i_16_n_0,
   I4 => W_46_7_i_17_n_0,
   O => W_46_7_i_5_n_0
);
W_46_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_46_7_i_2_n_0,
   I1 => W_46_11_i_16_n_0,
   I2 => x56_out_17,
   I3 => x56_out_24,
   I4 => x56_out_26,
   I5 => W_46_11_i_17_n_0,
   O => W_46_7_i_6_n_0
);
W_46_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_46_7_i_3_n_0,
   I1 => W_46_7_i_10_n_0,
   I2 => x56_out_16,
   I3 => x56_out_23,
   I4 => x56_out_25,
   I5 => W_46_7_i_11_n_0,
   O => W_46_7_i_7_n_0
);
W_46_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_46_7_i_4_n_0,
   I1 => W_46_7_i_12_n_0,
   I2 => x56_out_15,
   I3 => x56_out_22,
   I4 => x56_out_24,
   I5 => W_46_7_i_13_n_0,
   O => W_46_7_i_8_n_0
);
W_46_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_46_7_i_5_n_0,
   I1 => W_46_7_i_14_n_0,
   I2 => x56_out_14,
   I3 => x56_out_21,
   I4 => x56_out_23,
   I5 => W_46_7_i_15_n_0,
   O => W_46_7_i_9_n_0
);
W_47_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x94_out_10,
   I1 => x68_out_10,
   I2 => x92_out_28,
   I3 => x92_out_17,
   I4 => x92_out_13,
   O => W_47_11_i_10_n_0
);
W_47_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x68_out_9,
   I1 => x92_out_12,
   I2 => x92_out_16,
   I3 => x92_out_27,
   I4 => x94_out_9,
   O => W_47_11_i_11_n_0
);
W_47_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x94_out_9,
   I1 => x68_out_9,
   I2 => x92_out_27,
   I3 => x92_out_16,
   I4 => x92_out_12,
   O => W_47_11_i_12_n_0
);
W_47_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x68_out_8,
   I1 => x92_out_11,
   I2 => x92_out_15,
   I3 => x92_out_26,
   I4 => x94_out_8,
   O => W_47_11_i_13_n_0
);
W_47_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x94_out_8,
   I1 => x68_out_8,
   I2 => x92_out_26,
   I3 => x92_out_15,
   I4 => x92_out_11,
   O => W_47_11_i_14_n_0
);
W_47_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x68_out_7,
   I1 => x92_out_10,
   I2 => x92_out_14,
   I3 => x92_out_25,
   I4 => x94_out_7,
   O => W_47_11_i_15_n_0
);
W_47_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x94_out_7,
   I1 => x68_out_7,
   I2 => x92_out_25,
   I3 => x92_out_14,
   I4 => x92_out_10,
   O => W_47_11_i_16_n_0
);
W_47_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x68_out_6,
   I1 => x92_out_9,
   I2 => x92_out_13,
   I3 => x92_out_24,
   I4 => x94_out_6,
   O => W_47_11_i_17_n_0
);
W_47_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x53_out_20,
   I1 => x53_out_27,
   I2 => x53_out_29,
   I3 => W_47_11_i_10_n_0,
   I4 => W_47_11_i_11_n_0,
   O => W_47_11_i_2_n_0
);
W_47_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x53_out_19,
   I1 => x53_out_26,
   I2 => x53_out_28,
   I3 => W_47_11_i_12_n_0,
   I4 => W_47_11_i_13_n_0,
   O => W_47_11_i_3_n_0
);
W_47_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x53_out_18,
   I1 => x53_out_25,
   I2 => x53_out_27,
   I3 => W_47_11_i_14_n_0,
   I4 => W_47_11_i_15_n_0,
   O => W_47_11_i_4_n_0
);
W_47_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x53_out_17,
   I1 => x53_out_24,
   I2 => x53_out_26,
   I3 => W_47_11_i_16_n_0,
   I4 => W_47_11_i_17_n_0,
   O => W_47_11_i_5_n_0
);
W_47_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_47_11_i_2_n_0,
   I1 => W_47_15_i_16_n_0,
   I2 => x53_out_21,
   I3 => x53_out_28,
   I4 => x53_out_30,
   I5 => W_47_15_i_17_n_0,
   O => W_47_11_i_6_n_0
);
W_47_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_47_11_i_3_n_0,
   I1 => W_47_11_i_10_n_0,
   I2 => x53_out_20,
   I3 => x53_out_27,
   I4 => x53_out_29,
   I5 => W_47_11_i_11_n_0,
   O => W_47_11_i_7_n_0
);
W_47_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_47_11_i_4_n_0,
   I1 => W_47_11_i_12_n_0,
   I2 => x53_out_19,
   I3 => x53_out_26,
   I4 => x53_out_28,
   I5 => W_47_11_i_13_n_0,
   O => W_47_11_i_8_n_0
);
W_47_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_47_11_i_5_n_0,
   I1 => W_47_11_i_14_n_0,
   I2 => x53_out_18,
   I3 => x53_out_25,
   I4 => x53_out_27,
   I5 => W_47_11_i_15_n_0,
   O => W_47_11_i_9_n_0
);
W_47_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x94_out_14,
   I1 => x68_out_14,
   I2 => x92_out_0,
   I3 => x92_out_21,
   I4 => x92_out_17,
   O => W_47_15_i_10_n_0
);
W_47_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x68_out_13,
   I1 => x92_out_16,
   I2 => x92_out_20,
   I3 => x92_out_31,
   I4 => x94_out_13,
   O => W_47_15_i_11_n_0
);
W_47_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x94_out_13,
   I1 => x68_out_13,
   I2 => x92_out_31,
   I3 => x92_out_20,
   I4 => x92_out_16,
   O => W_47_15_i_12_n_0
);
W_47_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x68_out_12,
   I1 => x92_out_15,
   I2 => x92_out_19,
   I3 => x92_out_30,
   I4 => x94_out_12,
   O => W_47_15_i_13_n_0
);
W_47_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x94_out_12,
   I1 => x68_out_12,
   I2 => x92_out_30,
   I3 => x92_out_19,
   I4 => x92_out_15,
   O => W_47_15_i_14_n_0
);
W_47_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x68_out_11,
   I1 => x92_out_14,
   I2 => x92_out_18,
   I3 => x92_out_29,
   I4 => x94_out_11,
   O => W_47_15_i_15_n_0
);
W_47_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x94_out_11,
   I1 => x68_out_11,
   I2 => x92_out_29,
   I3 => x92_out_18,
   I4 => x92_out_14,
   O => W_47_15_i_16_n_0
);
W_47_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x68_out_10,
   I1 => x92_out_13,
   I2 => x92_out_17,
   I3 => x92_out_28,
   I4 => x94_out_10,
   O => W_47_15_i_17_n_0
);
W_47_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x53_out_24,
   I1 => x53_out_31,
   I2 => x53_out_1,
   I3 => W_47_15_i_10_n_0,
   I4 => W_47_15_i_11_n_0,
   O => W_47_15_i_2_n_0
);
W_47_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x53_out_23,
   I1 => x53_out_30,
   I2 => x53_out_0,
   I3 => W_47_15_i_12_n_0,
   I4 => W_47_15_i_13_n_0,
   O => W_47_15_i_3_n_0
);
W_47_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x53_out_22,
   I1 => x53_out_29,
   I2 => x53_out_31,
   I3 => W_47_15_i_14_n_0,
   I4 => W_47_15_i_15_n_0,
   O => W_47_15_i_4_n_0
);
W_47_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x53_out_21,
   I1 => x53_out_28,
   I2 => x53_out_30,
   I3 => W_47_15_i_16_n_0,
   I4 => W_47_15_i_17_n_0,
   O => W_47_15_i_5_n_0
);
W_47_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_47_15_i_2_n_0,
   I1 => W_47_19_i_16_n_0,
   I2 => x53_out_25,
   I3 => x53_out_0,
   I4 => x53_out_2,
   I5 => W_47_19_i_17_n_0,
   O => W_47_15_i_6_n_0
);
W_47_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_47_15_i_3_n_0,
   I1 => W_47_15_i_10_n_0,
   I2 => x53_out_24,
   I3 => x53_out_31,
   I4 => x53_out_1,
   I5 => W_47_15_i_11_n_0,
   O => W_47_15_i_7_n_0
);
W_47_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_47_15_i_4_n_0,
   I1 => W_47_15_i_12_n_0,
   I2 => x53_out_23,
   I3 => x53_out_30,
   I4 => x53_out_0,
   I5 => W_47_15_i_13_n_0,
   O => W_47_15_i_8_n_0
);
W_47_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_47_15_i_5_n_0,
   I1 => W_47_15_i_14_n_0,
   I2 => x53_out_22,
   I3 => x53_out_29,
   I4 => x53_out_31,
   I5 => W_47_15_i_15_n_0,
   O => W_47_15_i_9_n_0
);
W_47_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x94_out_18,
   I1 => x68_out_18,
   I2 => x92_out_4,
   I3 => x92_out_25,
   I4 => x92_out_21,
   O => W_47_19_i_10_n_0
);
W_47_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x68_out_17,
   I1 => x92_out_20,
   I2 => x92_out_24,
   I3 => x92_out_3,
   I4 => x94_out_17,
   O => W_47_19_i_11_n_0
);
W_47_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x94_out_17,
   I1 => x68_out_17,
   I2 => x92_out_3,
   I3 => x92_out_24,
   I4 => x92_out_20,
   O => W_47_19_i_12_n_0
);
W_47_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x68_out_16,
   I1 => x92_out_19,
   I2 => x92_out_23,
   I3 => x92_out_2,
   I4 => x94_out_16,
   O => W_47_19_i_13_n_0
);
W_47_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x94_out_16,
   I1 => x68_out_16,
   I2 => x92_out_2,
   I3 => x92_out_23,
   I4 => x92_out_19,
   O => W_47_19_i_14_n_0
);
W_47_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x68_out_15,
   I1 => x92_out_18,
   I2 => x92_out_22,
   I3 => x92_out_1,
   I4 => x94_out_15,
   O => W_47_19_i_15_n_0
);
W_47_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x94_out_15,
   I1 => x68_out_15,
   I2 => x92_out_1,
   I3 => x92_out_22,
   I4 => x92_out_18,
   O => W_47_19_i_16_n_0
);
W_47_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x68_out_14,
   I1 => x92_out_17,
   I2 => x92_out_21,
   I3 => x92_out_0,
   I4 => x94_out_14,
   O => W_47_19_i_17_n_0
);
W_47_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x53_out_28,
   I1 => x53_out_3,
   I2 => x53_out_5,
   I3 => W_47_19_i_10_n_0,
   I4 => W_47_19_i_11_n_0,
   O => W_47_19_i_2_n_0
);
W_47_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x53_out_27,
   I1 => x53_out_2,
   I2 => x53_out_4,
   I3 => W_47_19_i_12_n_0,
   I4 => W_47_19_i_13_n_0,
   O => W_47_19_i_3_n_0
);
W_47_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x53_out_26,
   I1 => x53_out_1,
   I2 => x53_out_3,
   I3 => W_47_19_i_14_n_0,
   I4 => W_47_19_i_15_n_0,
   O => W_47_19_i_4_n_0
);
W_47_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x53_out_25,
   I1 => x53_out_0,
   I2 => x53_out_2,
   I3 => W_47_19_i_16_n_0,
   I4 => W_47_19_i_17_n_0,
   O => W_47_19_i_5_n_0
);
W_47_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_47_19_i_2_n_0,
   I1 => W_47_23_i_16_n_0,
   I2 => x53_out_29,
   I3 => x53_out_4,
   I4 => x53_out_6,
   I5 => W_47_23_i_17_n_0,
   O => W_47_19_i_6_n_0
);
W_47_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_47_19_i_3_n_0,
   I1 => W_47_19_i_10_n_0,
   I2 => x53_out_28,
   I3 => x53_out_3,
   I4 => x53_out_5,
   I5 => W_47_19_i_11_n_0,
   O => W_47_19_i_7_n_0
);
W_47_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_47_19_i_4_n_0,
   I1 => W_47_19_i_12_n_0,
   I2 => x53_out_27,
   I3 => x53_out_2,
   I4 => x53_out_4,
   I5 => W_47_19_i_13_n_0,
   O => W_47_19_i_8_n_0
);
W_47_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_47_19_i_5_n_0,
   I1 => W_47_19_i_14_n_0,
   I2 => x53_out_26,
   I3 => x53_out_1,
   I4 => x53_out_3,
   I5 => W_47_19_i_15_n_0,
   O => W_47_19_i_9_n_0
);
W_47_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x94_out_22,
   I1 => x68_out_22,
   I2 => x92_out_8,
   I3 => x92_out_29,
   I4 => x92_out_25,
   O => W_47_23_i_10_n_0
);
W_47_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x68_out_21,
   I1 => x92_out_24,
   I2 => x92_out_28,
   I3 => x92_out_7,
   I4 => x94_out_21,
   O => W_47_23_i_11_n_0
);
W_47_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x94_out_21,
   I1 => x68_out_21,
   I2 => x92_out_7,
   I3 => x92_out_28,
   I4 => x92_out_24,
   O => W_47_23_i_12_n_0
);
W_47_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x68_out_20,
   I1 => x92_out_23,
   I2 => x92_out_27,
   I3 => x92_out_6,
   I4 => x94_out_20,
   O => W_47_23_i_13_n_0
);
W_47_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x94_out_20,
   I1 => x68_out_20,
   I2 => x92_out_6,
   I3 => x92_out_27,
   I4 => x92_out_23,
   O => W_47_23_i_14_n_0
);
W_47_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x68_out_19,
   I1 => x92_out_22,
   I2 => x92_out_26,
   I3 => x92_out_5,
   I4 => x94_out_19,
   O => W_47_23_i_15_n_0
);
W_47_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x94_out_19,
   I1 => x68_out_19,
   I2 => x92_out_5,
   I3 => x92_out_26,
   I4 => x92_out_22,
   O => W_47_23_i_16_n_0
);
W_47_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x68_out_18,
   I1 => x92_out_21,
   I2 => x92_out_25,
   I3 => x92_out_4,
   I4 => x94_out_18,
   O => W_47_23_i_17_n_0
);
W_47_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x53_out_7,
   I1 => x53_out_9,
   I2 => W_47_23_i_10_n_0,
   I3 => W_47_23_i_11_n_0,
   O => W_47_23_i_2_n_0
);
W_47_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x53_out_31,
   I1 => x53_out_6,
   I2 => x53_out_8,
   I3 => W_47_23_i_12_n_0,
   I4 => W_47_23_i_13_n_0,
   O => W_47_23_i_3_n_0
);
W_47_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x53_out_30,
   I1 => x53_out_5,
   I2 => x53_out_7,
   I3 => W_47_23_i_14_n_0,
   I4 => W_47_23_i_15_n_0,
   O => W_47_23_i_4_n_0
);
W_47_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x53_out_29,
   I1 => x53_out_4,
   I2 => x53_out_6,
   I3 => W_47_23_i_16_n_0,
   I4 => W_47_23_i_17_n_0,
   O => W_47_23_i_5_n_0
);
W_47_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x53_out_8,
   I1 => x53_out_10,
   I2 => W_47_27_i_16_n_0,
   I3 => W_47_27_i_17_n_0,
   I4 => W_47_23_i_2_n_0,
   O => W_47_23_i_6_n_0
);
W_47_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x53_out_7,
   I1 => x53_out_9,
   I2 => W_47_23_i_10_n_0,
   I3 => W_47_23_i_11_n_0,
   I4 => W_47_23_i_3_n_0,
   O => W_47_23_i_7_n_0
);
W_47_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_47_23_i_4_n_0,
   I1 => W_47_23_i_12_n_0,
   I2 => x53_out_31,
   I3 => x53_out_6,
   I4 => x53_out_8,
   I5 => W_47_23_i_13_n_0,
   O => W_47_23_i_8_n_0
);
W_47_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_47_23_i_5_n_0,
   I1 => W_47_23_i_14_n_0,
   I2 => x53_out_30,
   I3 => x53_out_5,
   I4 => x53_out_7,
   I5 => W_47_23_i_15_n_0,
   O => W_47_23_i_9_n_0
);
W_47_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x94_out_26,
   I1 => x68_out_26,
   I2 => x92_out_12,
   I3 => x92_out_1,
   I4 => x92_out_29,
   O => W_47_27_i_10_n_0
);
W_47_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x68_out_25,
   I1 => x92_out_28,
   I2 => x92_out_0,
   I3 => x92_out_11,
   I4 => x94_out_25,
   O => W_47_27_i_11_n_0
);
W_47_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x94_out_25,
   I1 => x68_out_25,
   I2 => x92_out_11,
   I3 => x92_out_0,
   I4 => x92_out_28,
   O => W_47_27_i_12_n_0
);
W_47_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x68_out_24,
   I1 => x92_out_27,
   I2 => x92_out_31,
   I3 => x92_out_10,
   I4 => x94_out_24,
   O => W_47_27_i_13_n_0
);
W_47_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x94_out_24,
   I1 => x68_out_24,
   I2 => x92_out_10,
   I3 => x92_out_31,
   I4 => x92_out_27,
   O => W_47_27_i_14_n_0
);
W_47_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x68_out_23,
   I1 => x92_out_26,
   I2 => x92_out_30,
   I3 => x92_out_9,
   I4 => x94_out_23,
   O => W_47_27_i_15_n_0
);
W_47_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x94_out_23,
   I1 => x68_out_23,
   I2 => x92_out_9,
   I3 => x92_out_30,
   I4 => x92_out_26,
   O => W_47_27_i_16_n_0
);
W_47_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x68_out_22,
   I1 => x92_out_25,
   I2 => x92_out_29,
   I3 => x92_out_8,
   I4 => x94_out_22,
   O => W_47_27_i_17_n_0
);
W_47_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x53_out_11,
   I1 => x53_out_13,
   I2 => W_47_27_i_10_n_0,
   I3 => W_47_27_i_11_n_0,
   O => W_47_27_i_2_n_0
);
W_47_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x53_out_10,
   I1 => x53_out_12,
   I2 => W_47_27_i_12_n_0,
   I3 => W_47_27_i_13_n_0,
   O => W_47_27_i_3_n_0
);
W_47_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x53_out_9,
   I1 => x53_out_11,
   I2 => W_47_27_i_14_n_0,
   I3 => W_47_27_i_15_n_0,
   O => W_47_27_i_4_n_0
);
W_47_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x53_out_8,
   I1 => x53_out_10,
   I2 => W_47_27_i_16_n_0,
   I3 => W_47_27_i_17_n_0,
   O => W_47_27_i_5_n_0
);
W_47_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x53_out_12,
   I1 => x53_out_14,
   I2 => W_47_31_i_13_n_0,
   I3 => W_47_31_i_14_n_0,
   I4 => W_47_27_i_2_n_0,
   O => W_47_27_i_6_n_0
);
W_47_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x53_out_11,
   I1 => x53_out_13,
   I2 => W_47_27_i_10_n_0,
   I3 => W_47_27_i_11_n_0,
   I4 => W_47_27_i_3_n_0,
   O => W_47_27_i_7_n_0
);
W_47_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x53_out_10,
   I1 => x53_out_12,
   I2 => W_47_27_i_12_n_0,
   I3 => W_47_27_i_13_n_0,
   I4 => W_47_27_i_4_n_0,
   O => W_47_27_i_8_n_0
);
W_47_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x53_out_9,
   I1 => x53_out_11,
   I2 => W_47_27_i_14_n_0,
   I3 => W_47_27_i_15_n_0,
   I4 => W_47_27_i_5_n_0,
   O => W_47_27_i_9_n_0
);
W_47_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x68_out_28,
   I1 => x92_out_31,
   I2 => x92_out_3,
   I3 => x92_out_14,
   I4 => x94_out_28,
   O => W_47_31_i_10_n_0
);
W_47_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x94_out_28,
   I1 => x68_out_28,
   I2 => x92_out_14,
   I3 => x92_out_3,
   I4 => x92_out_31,
   O => W_47_31_i_11_n_0
);
W_47_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x68_out_27,
   I1 => x92_out_30,
   I2 => x92_out_2,
   I3 => x92_out_13,
   I4 => x94_out_27,
   O => W_47_31_i_12_n_0
);
W_47_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x94_out_27,
   I1 => x68_out_27,
   I2 => x92_out_13,
   I3 => x92_out_2,
   I4 => x92_out_30,
   O => W_47_31_i_13_n_0
);
W_47_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x68_out_26,
   I1 => x92_out_29,
   I2 => x92_out_1,
   I3 => x92_out_12,
   I4 => x94_out_26,
   O => W_47_31_i_14_n_0
);
W_47_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x68_out_29,
   I1 => x92_out_4,
   I2 => x92_out_15,
   I3 => x94_out_29,
   O => W_47_31_i_15_n_0
);
W_47_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x53_out_17,
   I1 => x53_out_15,
   O => SIGMA_LCASE_1139_out_0_30
);
W_47_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => x92_out_6,
   I1 => x92_out_17,
   I2 => x68_out_31,
   I3 => x94_out_31,
   I4 => x53_out_16,
   I5 => x53_out_18,
   O => W_47_31_i_17_n_0
);
W_47_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x92_out_16,
   I1 => x92_out_5,
   O => SIGMA_LCASE_0135_out_30
);
W_47_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x94_out_30,
   I1 => x68_out_30,
   I2 => x92_out_16,
   I3 => x92_out_5,
   O => W_47_31_i_19_n_0
);
W_47_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x53_out_14,
   I1 => x53_out_16,
   I2 => W_47_31_i_9_n_0,
   I3 => W_47_31_i_10_n_0,
   O => W_47_31_i_2_n_0
);
W_47_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x53_out_13,
   I1 => x53_out_15,
   I2 => W_47_31_i_11_n_0,
   I3 => W_47_31_i_12_n_0,
   O => W_47_31_i_3_n_0
);
W_47_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x53_out_12,
   I1 => x53_out_14,
   I2 => W_47_31_i_13_n_0,
   I3 => W_47_31_i_14_n_0,
   O => W_47_31_i_4_n_0
);
W_47_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_47_31_i_15_n_0,
   I1 => SIGMA_LCASE_1139_out_0_30,
   I2 => W_47_31_i_17_n_0,
   I3 => x68_out_30,
   I4 => SIGMA_LCASE_0135_out_30,
   I5 => x94_out_30,
   O => W_47_31_i_5_n_0
);
W_47_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_47_31_i_2_n_0,
   I1 => W_47_31_i_19_n_0,
   I2 => x53_out_15,
   I3 => x53_out_17,
   I4 => W_47_31_i_15_n_0,
   O => W_47_31_i_6_n_0
);
W_47_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x53_out_14,
   I1 => x53_out_16,
   I2 => W_47_31_i_9_n_0,
   I3 => W_47_31_i_10_n_0,
   I4 => W_47_31_i_3_n_0,
   O => W_47_31_i_7_n_0
);
W_47_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x53_out_13,
   I1 => x53_out_15,
   I2 => W_47_31_i_11_n_0,
   I3 => W_47_31_i_12_n_0,
   I4 => W_47_31_i_4_n_0,
   O => W_47_31_i_8_n_0
);
W_47_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x94_out_29,
   I1 => x68_out_29,
   I2 => x92_out_15,
   I3 => x92_out_4,
   O => W_47_31_i_9_n_0
);
W_47_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x94_out_2,
   I1 => x68_out_2,
   I2 => x92_out_20,
   I3 => x92_out_9,
   I4 => x92_out_5,
   O => W_47_3_i_10_n_0
);
W_47_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x68_out_1,
   I1 => x92_out_4,
   I2 => x92_out_8,
   I3 => x92_out_19,
   I4 => x94_out_1,
   O => W_47_3_i_11_n_0
);
W_47_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x92_out_19,
   I1 => x92_out_8,
   I2 => x92_out_4,
   O => SIGMA_LCASE_0135_out_1
);
W_47_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x53_out_21,
   I1 => x53_out_19,
   I2 => x53_out_12,
   O => SIGMA_LCASE_1139_out_0_2
);
W_47_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x53_out_20,
   I1 => x53_out_18,
   I2 => x53_out_11,
   O => SIGMA_LCASE_1139_out_1
);
W_47_3_i_15 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x94_out_1,
   I1 => x68_out_1,
   I2 => x92_out_19,
   I3 => x92_out_8,
   I4 => x92_out_4,
   O => W_47_3_i_15_n_0
);
W_47_3_i_16 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x92_out_18,
   I1 => x92_out_7,
   I2 => x92_out_3,
   O => SIGMA_LCASE_0135_out_0
);
W_47_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x53_out_12,
   I1 => x53_out_19,
   I2 => x53_out_21,
   I3 => W_47_3_i_10_n_0,
   I4 => W_47_3_i_11_n_0,
   O => W_47_3_i_2_n_0
);
W_47_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_47_3_i_11_n_0,
   I1 => x53_out_21,
   I2 => x53_out_19,
   I3 => x53_out_12,
   I4 => W_47_3_i_10_n_0,
   O => W_47_3_i_3_n_0
);
W_47_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_0135_out_1,
   I1 => x68_out_1,
   I2 => x94_out_1,
   I3 => x53_out_11,
   I4 => x53_out_18,
   I5 => x53_out_20,
   O => W_47_3_i_4_n_0
);
W_47_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x94_out_0,
   I1 => x68_out_0,
   I2 => x92_out_18,
   I3 => x92_out_7,
   I4 => x92_out_3,
   O => W_47_3_i_5_n_0
);
W_47_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_47_3_i_2_n_0,
   I1 => W_47_7_i_16_n_0,
   I2 => x53_out_13,
   I3 => x53_out_20,
   I4 => x53_out_22,
   I5 => W_47_7_i_17_n_0,
   O => W_47_3_i_6_n_0
);
W_47_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_47_3_i_10_n_0,
   I1 => SIGMA_LCASE_1139_out_0_2,
   I2 => x94_out_1,
   I3 => x68_out_1,
   I4 => SIGMA_LCASE_0135_out_1,
   I5 => SIGMA_LCASE_1139_out_1,
   O => W_47_3_i_7_n_0
);
W_47_3_i_8 : LUT5
  generic map(
   INIT => X"99969666"
  )
 port map (
   I0 => SIGMA_LCASE_1139_out_1,
   I1 => W_47_3_i_15_n_0,
   I2 => x94_out_0,
   I3 => SIGMA_LCASE_0135_out_0,
   I4 => x68_out_0,
   O => W_47_3_i_8_n_0
);
W_47_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_47_3_i_5_n_0,
   I1 => x53_out_10,
   I2 => x53_out_17,
   I3 => x53_out_19,
   O => W_47_3_i_9_n_0
);
W_47_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x94_out_6,
   I1 => x68_out_6,
   I2 => x92_out_24,
   I3 => x92_out_13,
   I4 => x92_out_9,
   O => W_47_7_i_10_n_0
);
W_47_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x68_out_5,
   I1 => x92_out_8,
   I2 => x92_out_12,
   I3 => x92_out_23,
   I4 => x94_out_5,
   O => W_47_7_i_11_n_0
);
W_47_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x94_out_5,
   I1 => x68_out_5,
   I2 => x92_out_23,
   I3 => x92_out_12,
   I4 => x92_out_8,
   O => W_47_7_i_12_n_0
);
W_47_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x68_out_4,
   I1 => x92_out_7,
   I2 => x92_out_11,
   I3 => x92_out_22,
   I4 => x94_out_4,
   O => W_47_7_i_13_n_0
);
W_47_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x94_out_4,
   I1 => x68_out_4,
   I2 => x92_out_22,
   I3 => x92_out_11,
   I4 => x92_out_7,
   O => W_47_7_i_14_n_0
);
W_47_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x68_out_3,
   I1 => x92_out_6,
   I2 => x92_out_10,
   I3 => x92_out_21,
   I4 => x94_out_3,
   O => W_47_7_i_15_n_0
);
W_47_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x94_out_3,
   I1 => x68_out_3,
   I2 => x92_out_21,
   I3 => x92_out_10,
   I4 => x92_out_6,
   O => W_47_7_i_16_n_0
);
W_47_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x68_out_2,
   I1 => x92_out_5,
   I2 => x92_out_9,
   I3 => x92_out_20,
   I4 => x94_out_2,
   O => W_47_7_i_17_n_0
);
W_47_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x53_out_16,
   I1 => x53_out_23,
   I2 => x53_out_25,
   I3 => W_47_7_i_10_n_0,
   I4 => W_47_7_i_11_n_0,
   O => W_47_7_i_2_n_0
);
W_47_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x53_out_15,
   I1 => x53_out_22,
   I2 => x53_out_24,
   I3 => W_47_7_i_12_n_0,
   I4 => W_47_7_i_13_n_0,
   O => W_47_7_i_3_n_0
);
W_47_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x53_out_14,
   I1 => x53_out_21,
   I2 => x53_out_23,
   I3 => W_47_7_i_14_n_0,
   I4 => W_47_7_i_15_n_0,
   O => W_47_7_i_4_n_0
);
W_47_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x53_out_13,
   I1 => x53_out_20,
   I2 => x53_out_22,
   I3 => W_47_7_i_16_n_0,
   I4 => W_47_7_i_17_n_0,
   O => W_47_7_i_5_n_0
);
W_47_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_47_7_i_2_n_0,
   I1 => W_47_11_i_16_n_0,
   I2 => x53_out_17,
   I3 => x53_out_24,
   I4 => x53_out_26,
   I5 => W_47_11_i_17_n_0,
   O => W_47_7_i_6_n_0
);
W_47_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_47_7_i_3_n_0,
   I1 => W_47_7_i_10_n_0,
   I2 => x53_out_16,
   I3 => x53_out_23,
   I4 => x53_out_25,
   I5 => W_47_7_i_11_n_0,
   O => W_47_7_i_7_n_0
);
W_47_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_47_7_i_4_n_0,
   I1 => W_47_7_i_12_n_0,
   I2 => x53_out_15,
   I3 => x53_out_22,
   I4 => x53_out_24,
   I5 => W_47_7_i_13_n_0,
   O => W_47_7_i_8_n_0
);
W_47_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_47_7_i_5_n_0,
   I1 => W_47_7_i_14_n_0,
   I2 => x53_out_14,
   I3 => x53_out_21,
   I4 => x53_out_23,
   I5 => W_47_7_i_15_n_0,
   O => W_47_7_i_9_n_0
);
W_48_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x92_out_10,
   I1 => x65_out_10,
   I2 => x89_out_28,
   I3 => x89_out_17,
   I4 => x89_out_13,
   O => W_48_11_i_10_n_0
);
W_48_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x65_out_9,
   I1 => x89_out_12,
   I2 => x89_out_16,
   I3 => x89_out_27,
   I4 => x92_out_9,
   O => W_48_11_i_11_n_0
);
W_48_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x92_out_9,
   I1 => x65_out_9,
   I2 => x89_out_27,
   I3 => x89_out_16,
   I4 => x89_out_12,
   O => W_48_11_i_12_n_0
);
W_48_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x65_out_8,
   I1 => x89_out_11,
   I2 => x89_out_15,
   I3 => x89_out_26,
   I4 => x92_out_8,
   O => W_48_11_i_13_n_0
);
W_48_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x92_out_8,
   I1 => x65_out_8,
   I2 => x89_out_26,
   I3 => x89_out_15,
   I4 => x89_out_11,
   O => W_48_11_i_14_n_0
);
W_48_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x65_out_7,
   I1 => x89_out_10,
   I2 => x89_out_14,
   I3 => x89_out_25,
   I4 => x92_out_7,
   O => W_48_11_i_15_n_0
);
W_48_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x92_out_7,
   I1 => x65_out_7,
   I2 => x89_out_25,
   I3 => x89_out_14,
   I4 => x89_out_10,
   O => W_48_11_i_16_n_0
);
W_48_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x65_out_6,
   I1 => x89_out_9,
   I2 => x89_out_13,
   I3 => x89_out_24,
   I4 => x92_out_6,
   O => W_48_11_i_17_n_0
);
W_48_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x50_out_20,
   I1 => x50_out_27,
   I2 => x50_out_29,
   I3 => W_48_11_i_10_n_0,
   I4 => W_48_11_i_11_n_0,
   O => W_48_11_i_2_n_0
);
W_48_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x50_out_19,
   I1 => x50_out_26,
   I2 => x50_out_28,
   I3 => W_48_11_i_12_n_0,
   I4 => W_48_11_i_13_n_0,
   O => W_48_11_i_3_n_0
);
W_48_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x50_out_18,
   I1 => x50_out_25,
   I2 => x50_out_27,
   I3 => W_48_11_i_14_n_0,
   I4 => W_48_11_i_15_n_0,
   O => W_48_11_i_4_n_0
);
W_48_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x50_out_17,
   I1 => x50_out_24,
   I2 => x50_out_26,
   I3 => W_48_11_i_16_n_0,
   I4 => W_48_11_i_17_n_0,
   O => W_48_11_i_5_n_0
);
W_48_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_48_11_i_2_n_0,
   I1 => W_48_15_i_16_n_0,
   I2 => x50_out_21,
   I3 => x50_out_28,
   I4 => x50_out_30,
   I5 => W_48_15_i_17_n_0,
   O => W_48_11_i_6_n_0
);
W_48_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_48_11_i_3_n_0,
   I1 => W_48_11_i_10_n_0,
   I2 => x50_out_20,
   I3 => x50_out_27,
   I4 => x50_out_29,
   I5 => W_48_11_i_11_n_0,
   O => W_48_11_i_7_n_0
);
W_48_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_48_11_i_4_n_0,
   I1 => W_48_11_i_12_n_0,
   I2 => x50_out_19,
   I3 => x50_out_26,
   I4 => x50_out_28,
   I5 => W_48_11_i_13_n_0,
   O => W_48_11_i_8_n_0
);
W_48_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_48_11_i_5_n_0,
   I1 => W_48_11_i_14_n_0,
   I2 => x50_out_18,
   I3 => x50_out_25,
   I4 => x50_out_27,
   I5 => W_48_11_i_15_n_0,
   O => W_48_11_i_9_n_0
);
W_48_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x92_out_14,
   I1 => x65_out_14,
   I2 => x89_out_0,
   I3 => x89_out_21,
   I4 => x89_out_17,
   O => W_48_15_i_10_n_0
);
W_48_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x65_out_13,
   I1 => x89_out_16,
   I2 => x89_out_20,
   I3 => x89_out_31,
   I4 => x92_out_13,
   O => W_48_15_i_11_n_0
);
W_48_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x92_out_13,
   I1 => x65_out_13,
   I2 => x89_out_31,
   I3 => x89_out_20,
   I4 => x89_out_16,
   O => W_48_15_i_12_n_0
);
W_48_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x65_out_12,
   I1 => x89_out_15,
   I2 => x89_out_19,
   I3 => x89_out_30,
   I4 => x92_out_12,
   O => W_48_15_i_13_n_0
);
W_48_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x92_out_12,
   I1 => x65_out_12,
   I2 => x89_out_30,
   I3 => x89_out_19,
   I4 => x89_out_15,
   O => W_48_15_i_14_n_0
);
W_48_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x65_out_11,
   I1 => x89_out_14,
   I2 => x89_out_18,
   I3 => x89_out_29,
   I4 => x92_out_11,
   O => W_48_15_i_15_n_0
);
W_48_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x92_out_11,
   I1 => x65_out_11,
   I2 => x89_out_29,
   I3 => x89_out_18,
   I4 => x89_out_14,
   O => W_48_15_i_16_n_0
);
W_48_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x65_out_10,
   I1 => x89_out_13,
   I2 => x89_out_17,
   I3 => x89_out_28,
   I4 => x92_out_10,
   O => W_48_15_i_17_n_0
);
W_48_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x50_out_24,
   I1 => x50_out_31,
   I2 => x50_out_1,
   I3 => W_48_15_i_10_n_0,
   I4 => W_48_15_i_11_n_0,
   O => W_48_15_i_2_n_0
);
W_48_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x50_out_23,
   I1 => x50_out_30,
   I2 => x50_out_0,
   I3 => W_48_15_i_12_n_0,
   I4 => W_48_15_i_13_n_0,
   O => W_48_15_i_3_n_0
);
W_48_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x50_out_22,
   I1 => x50_out_29,
   I2 => x50_out_31,
   I3 => W_48_15_i_14_n_0,
   I4 => W_48_15_i_15_n_0,
   O => W_48_15_i_4_n_0
);
W_48_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x50_out_21,
   I1 => x50_out_28,
   I2 => x50_out_30,
   I3 => W_48_15_i_16_n_0,
   I4 => W_48_15_i_17_n_0,
   O => W_48_15_i_5_n_0
);
W_48_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_48_15_i_2_n_0,
   I1 => W_48_19_i_16_n_0,
   I2 => x50_out_25,
   I3 => x50_out_0,
   I4 => x50_out_2,
   I5 => W_48_19_i_17_n_0,
   O => W_48_15_i_6_n_0
);
W_48_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_48_15_i_3_n_0,
   I1 => W_48_15_i_10_n_0,
   I2 => x50_out_24,
   I3 => x50_out_31,
   I4 => x50_out_1,
   I5 => W_48_15_i_11_n_0,
   O => W_48_15_i_7_n_0
);
W_48_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_48_15_i_4_n_0,
   I1 => W_48_15_i_12_n_0,
   I2 => x50_out_23,
   I3 => x50_out_30,
   I4 => x50_out_0,
   I5 => W_48_15_i_13_n_0,
   O => W_48_15_i_8_n_0
);
W_48_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_48_15_i_5_n_0,
   I1 => W_48_15_i_14_n_0,
   I2 => x50_out_22,
   I3 => x50_out_29,
   I4 => x50_out_31,
   I5 => W_48_15_i_15_n_0,
   O => W_48_15_i_9_n_0
);
W_48_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x92_out_18,
   I1 => x65_out_18,
   I2 => x89_out_4,
   I3 => x89_out_25,
   I4 => x89_out_21,
   O => W_48_19_i_10_n_0
);
W_48_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x65_out_17,
   I1 => x89_out_20,
   I2 => x89_out_24,
   I3 => x89_out_3,
   I4 => x92_out_17,
   O => W_48_19_i_11_n_0
);
W_48_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x92_out_17,
   I1 => x65_out_17,
   I2 => x89_out_3,
   I3 => x89_out_24,
   I4 => x89_out_20,
   O => W_48_19_i_12_n_0
);
W_48_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x65_out_16,
   I1 => x89_out_19,
   I2 => x89_out_23,
   I3 => x89_out_2,
   I4 => x92_out_16,
   O => W_48_19_i_13_n_0
);
W_48_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x92_out_16,
   I1 => x65_out_16,
   I2 => x89_out_2,
   I3 => x89_out_23,
   I4 => x89_out_19,
   O => W_48_19_i_14_n_0
);
W_48_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x65_out_15,
   I1 => x89_out_18,
   I2 => x89_out_22,
   I3 => x89_out_1,
   I4 => x92_out_15,
   O => W_48_19_i_15_n_0
);
W_48_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x92_out_15,
   I1 => x65_out_15,
   I2 => x89_out_1,
   I3 => x89_out_22,
   I4 => x89_out_18,
   O => W_48_19_i_16_n_0
);
W_48_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x65_out_14,
   I1 => x89_out_17,
   I2 => x89_out_21,
   I3 => x89_out_0,
   I4 => x92_out_14,
   O => W_48_19_i_17_n_0
);
W_48_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x50_out_28,
   I1 => x50_out_3,
   I2 => x50_out_5,
   I3 => W_48_19_i_10_n_0,
   I4 => W_48_19_i_11_n_0,
   O => W_48_19_i_2_n_0
);
W_48_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x50_out_27,
   I1 => x50_out_2,
   I2 => x50_out_4,
   I3 => W_48_19_i_12_n_0,
   I4 => W_48_19_i_13_n_0,
   O => W_48_19_i_3_n_0
);
W_48_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x50_out_26,
   I1 => x50_out_1,
   I2 => x50_out_3,
   I3 => W_48_19_i_14_n_0,
   I4 => W_48_19_i_15_n_0,
   O => W_48_19_i_4_n_0
);
W_48_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x50_out_25,
   I1 => x50_out_0,
   I2 => x50_out_2,
   I3 => W_48_19_i_16_n_0,
   I4 => W_48_19_i_17_n_0,
   O => W_48_19_i_5_n_0
);
W_48_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_48_19_i_2_n_0,
   I1 => W_48_23_i_16_n_0,
   I2 => x50_out_29,
   I3 => x50_out_4,
   I4 => x50_out_6,
   I5 => W_48_23_i_17_n_0,
   O => W_48_19_i_6_n_0
);
W_48_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_48_19_i_3_n_0,
   I1 => W_48_19_i_10_n_0,
   I2 => x50_out_28,
   I3 => x50_out_3,
   I4 => x50_out_5,
   I5 => W_48_19_i_11_n_0,
   O => W_48_19_i_7_n_0
);
W_48_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_48_19_i_4_n_0,
   I1 => W_48_19_i_12_n_0,
   I2 => x50_out_27,
   I3 => x50_out_2,
   I4 => x50_out_4,
   I5 => W_48_19_i_13_n_0,
   O => W_48_19_i_8_n_0
);
W_48_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_48_19_i_5_n_0,
   I1 => W_48_19_i_14_n_0,
   I2 => x50_out_26,
   I3 => x50_out_1,
   I4 => x50_out_3,
   I5 => W_48_19_i_15_n_0,
   O => W_48_19_i_9_n_0
);
W_48_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x92_out_22,
   I1 => x65_out_22,
   I2 => x89_out_8,
   I3 => x89_out_29,
   I4 => x89_out_25,
   O => W_48_23_i_10_n_0
);
W_48_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x65_out_21,
   I1 => x89_out_24,
   I2 => x89_out_28,
   I3 => x89_out_7,
   I4 => x92_out_21,
   O => W_48_23_i_11_n_0
);
W_48_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x92_out_21,
   I1 => x65_out_21,
   I2 => x89_out_7,
   I3 => x89_out_28,
   I4 => x89_out_24,
   O => W_48_23_i_12_n_0
);
W_48_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x65_out_20,
   I1 => x89_out_23,
   I2 => x89_out_27,
   I3 => x89_out_6,
   I4 => x92_out_20,
   O => W_48_23_i_13_n_0
);
W_48_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x92_out_20,
   I1 => x65_out_20,
   I2 => x89_out_6,
   I3 => x89_out_27,
   I4 => x89_out_23,
   O => W_48_23_i_14_n_0
);
W_48_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x65_out_19,
   I1 => x89_out_22,
   I2 => x89_out_26,
   I3 => x89_out_5,
   I4 => x92_out_19,
   O => W_48_23_i_15_n_0
);
W_48_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x92_out_19,
   I1 => x65_out_19,
   I2 => x89_out_5,
   I3 => x89_out_26,
   I4 => x89_out_22,
   O => W_48_23_i_16_n_0
);
W_48_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x65_out_18,
   I1 => x89_out_21,
   I2 => x89_out_25,
   I3 => x89_out_4,
   I4 => x92_out_18,
   O => W_48_23_i_17_n_0
);
W_48_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x50_out_7,
   I1 => x50_out_9,
   I2 => W_48_23_i_10_n_0,
   I3 => W_48_23_i_11_n_0,
   O => W_48_23_i_2_n_0
);
W_48_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x50_out_31,
   I1 => x50_out_6,
   I2 => x50_out_8,
   I3 => W_48_23_i_12_n_0,
   I4 => W_48_23_i_13_n_0,
   O => W_48_23_i_3_n_0
);
W_48_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x50_out_30,
   I1 => x50_out_5,
   I2 => x50_out_7,
   I3 => W_48_23_i_14_n_0,
   I4 => W_48_23_i_15_n_0,
   O => W_48_23_i_4_n_0
);
W_48_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x50_out_29,
   I1 => x50_out_4,
   I2 => x50_out_6,
   I3 => W_48_23_i_16_n_0,
   I4 => W_48_23_i_17_n_0,
   O => W_48_23_i_5_n_0
);
W_48_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x50_out_8,
   I1 => x50_out_10,
   I2 => W_48_27_i_16_n_0,
   I3 => W_48_27_i_17_n_0,
   I4 => W_48_23_i_2_n_0,
   O => W_48_23_i_6_n_0
);
W_48_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x50_out_7,
   I1 => x50_out_9,
   I2 => W_48_23_i_10_n_0,
   I3 => W_48_23_i_11_n_0,
   I4 => W_48_23_i_3_n_0,
   O => W_48_23_i_7_n_0
);
W_48_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_48_23_i_4_n_0,
   I1 => W_48_23_i_12_n_0,
   I2 => x50_out_31,
   I3 => x50_out_6,
   I4 => x50_out_8,
   I5 => W_48_23_i_13_n_0,
   O => W_48_23_i_8_n_0
);
W_48_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_48_23_i_5_n_0,
   I1 => W_48_23_i_14_n_0,
   I2 => x50_out_30,
   I3 => x50_out_5,
   I4 => x50_out_7,
   I5 => W_48_23_i_15_n_0,
   O => W_48_23_i_9_n_0
);
W_48_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x92_out_26,
   I1 => x65_out_26,
   I2 => x89_out_12,
   I3 => x89_out_1,
   I4 => x89_out_29,
   O => W_48_27_i_10_n_0
);
W_48_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x65_out_25,
   I1 => x89_out_28,
   I2 => x89_out_0,
   I3 => x89_out_11,
   I4 => x92_out_25,
   O => W_48_27_i_11_n_0
);
W_48_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x92_out_25,
   I1 => x65_out_25,
   I2 => x89_out_11,
   I3 => x89_out_0,
   I4 => x89_out_28,
   O => W_48_27_i_12_n_0
);
W_48_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x65_out_24,
   I1 => x89_out_27,
   I2 => x89_out_31,
   I3 => x89_out_10,
   I4 => x92_out_24,
   O => W_48_27_i_13_n_0
);
W_48_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x92_out_24,
   I1 => x65_out_24,
   I2 => x89_out_10,
   I3 => x89_out_31,
   I4 => x89_out_27,
   O => W_48_27_i_14_n_0
);
W_48_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x65_out_23,
   I1 => x89_out_26,
   I2 => x89_out_30,
   I3 => x89_out_9,
   I4 => x92_out_23,
   O => W_48_27_i_15_n_0
);
W_48_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x92_out_23,
   I1 => x65_out_23,
   I2 => x89_out_9,
   I3 => x89_out_30,
   I4 => x89_out_26,
   O => W_48_27_i_16_n_0
);
W_48_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x65_out_22,
   I1 => x89_out_25,
   I2 => x89_out_29,
   I3 => x89_out_8,
   I4 => x92_out_22,
   O => W_48_27_i_17_n_0
);
W_48_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x50_out_11,
   I1 => x50_out_13,
   I2 => W_48_27_i_10_n_0,
   I3 => W_48_27_i_11_n_0,
   O => W_48_27_i_2_n_0
);
W_48_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x50_out_10,
   I1 => x50_out_12,
   I2 => W_48_27_i_12_n_0,
   I3 => W_48_27_i_13_n_0,
   O => W_48_27_i_3_n_0
);
W_48_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x50_out_9,
   I1 => x50_out_11,
   I2 => W_48_27_i_14_n_0,
   I3 => W_48_27_i_15_n_0,
   O => W_48_27_i_4_n_0
);
W_48_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x50_out_8,
   I1 => x50_out_10,
   I2 => W_48_27_i_16_n_0,
   I3 => W_48_27_i_17_n_0,
   O => W_48_27_i_5_n_0
);
W_48_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x50_out_12,
   I1 => x50_out_14,
   I2 => W_48_31_i_14_n_0,
   I3 => W_48_31_i_15_n_0,
   I4 => W_48_27_i_2_n_0,
   O => W_48_27_i_6_n_0
);
W_48_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x50_out_11,
   I1 => x50_out_13,
   I2 => W_48_27_i_10_n_0,
   I3 => W_48_27_i_11_n_0,
   I4 => W_48_27_i_3_n_0,
   O => W_48_27_i_7_n_0
);
W_48_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x50_out_10,
   I1 => x50_out_12,
   I2 => W_48_27_i_12_n_0,
   I3 => W_48_27_i_13_n_0,
   I4 => W_48_27_i_4_n_0,
   O => W_48_27_i_8_n_0
);
W_48_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x50_out_9,
   I1 => x50_out_11,
   I2 => W_48_27_i_14_n_0,
   I3 => W_48_27_i_15_n_0,
   I4 => W_48_27_i_5_n_0,
   O => W_48_27_i_9_n_0
);
W_48_31_i_1 : LUT2
  generic map(
   INIT => X"2"
  )
 port map (
   I0 => W_48,
   I1 => rst_IBUF,
   O => W_reg_48_0
);
W_48_31_i_10 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x92_out_29,
   I1 => x65_out_29,
   I2 => x89_out_15,
   I3 => x89_out_4,
   O => W_48_31_i_10_n_0
);
W_48_31_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x65_out_28,
   I1 => x89_out_31,
   I2 => x89_out_3,
   I3 => x89_out_14,
   I4 => x92_out_28,
   O => W_48_31_i_11_n_0
);
W_48_31_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x92_out_28,
   I1 => x65_out_28,
   I2 => x89_out_14,
   I3 => x89_out_3,
   I4 => x89_out_31,
   O => W_48_31_i_12_n_0
);
W_48_31_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x65_out_27,
   I1 => x89_out_30,
   I2 => x89_out_2,
   I3 => x89_out_13,
   I4 => x92_out_27,
   O => W_48_31_i_13_n_0
);
W_48_31_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x92_out_27,
   I1 => x65_out_27,
   I2 => x89_out_13,
   I3 => x89_out_2,
   I4 => x89_out_30,
   O => W_48_31_i_14_n_0
);
W_48_31_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x65_out_26,
   I1 => x89_out_29,
   I2 => x89_out_1,
   I3 => x89_out_12,
   I4 => x92_out_26,
   O => W_48_31_i_15_n_0
);
W_48_31_i_16 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x65_out_29,
   I1 => x89_out_4,
   I2 => x89_out_15,
   I3 => x92_out_29,
   O => W_48_31_i_16_n_0
);
W_48_31_i_17 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x50_out_17,
   I1 => x50_out_15,
   O => SIGMA_LCASE_1131_out_0_30
);
W_48_31_i_18 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => x89_out_6,
   I1 => x89_out_17,
   I2 => x65_out_31,
   I3 => x92_out_31,
   I4 => x50_out_16,
   I5 => x50_out_18,
   O => W_48_31_i_18_n_0
);
W_48_31_i_19 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x89_out_16,
   I1 => x89_out_5,
   O => SIGMA_LCASE_0127_out_30
);
W_48_31_i_20 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x92_out_30,
   I1 => x65_out_30,
   I2 => x89_out_16,
   I3 => x89_out_5,
   O => W_48_31_i_20_n_0
);
W_48_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x50_out_14,
   I1 => x50_out_16,
   I2 => W_48_31_i_10_n_0,
   I3 => W_48_31_i_11_n_0,
   O => W_48_31_i_3_n_0
);
W_48_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x50_out_13,
   I1 => x50_out_15,
   I2 => W_48_31_i_12_n_0,
   I3 => W_48_31_i_13_n_0,
   O => W_48_31_i_4_n_0
);
W_48_31_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x50_out_12,
   I1 => x50_out_14,
   I2 => W_48_31_i_14_n_0,
   I3 => W_48_31_i_15_n_0,
   O => W_48_31_i_5_n_0
);
W_48_31_i_6 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_48_31_i_16_n_0,
   I1 => SIGMA_LCASE_1131_out_0_30,
   I2 => W_48_31_i_18_n_0,
   I3 => x65_out_30,
   I4 => SIGMA_LCASE_0127_out_30,
   I5 => x92_out_30,
   O => W_48_31_i_6_n_0
);
W_48_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_48_31_i_3_n_0,
   I1 => W_48_31_i_20_n_0,
   I2 => x50_out_15,
   I3 => x50_out_17,
   I4 => W_48_31_i_16_n_0,
   O => W_48_31_i_7_n_0
);
W_48_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x50_out_14,
   I1 => x50_out_16,
   I2 => W_48_31_i_10_n_0,
   I3 => W_48_31_i_11_n_0,
   I4 => W_48_31_i_4_n_0,
   O => W_48_31_i_8_n_0
);
W_48_31_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x50_out_13,
   I1 => x50_out_15,
   I2 => W_48_31_i_12_n_0,
   I3 => W_48_31_i_13_n_0,
   I4 => W_48_31_i_5_n_0,
   O => W_48_31_i_9_n_0
);
W_48_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x92_out_2,
   I1 => x65_out_2,
   I2 => x89_out_20,
   I3 => x89_out_9,
   I4 => x89_out_5,
   O => W_48_3_i_10_n_0
);
W_48_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x65_out_1,
   I1 => x89_out_4,
   I2 => x89_out_8,
   I3 => x89_out_19,
   I4 => x92_out_1,
   O => W_48_3_i_11_n_0
);
W_48_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x89_out_19,
   I1 => x89_out_8,
   I2 => x89_out_4,
   O => SIGMA_LCASE_0127_out_1
);
W_48_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x50_out_21,
   I1 => x50_out_19,
   I2 => x50_out_12,
   O => SIGMA_LCASE_1131_out_0_2
);
W_48_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x50_out_20,
   I1 => x50_out_18,
   I2 => x50_out_11,
   O => SIGMA_LCASE_1131_out_1
);
W_48_3_i_15 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x92_out_1,
   I1 => x65_out_1,
   I2 => x89_out_19,
   I3 => x89_out_8,
   I4 => x89_out_4,
   O => W_48_3_i_15_n_0
);
W_48_3_i_16 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x89_out_18,
   I1 => x89_out_7,
   I2 => x89_out_3,
   O => SIGMA_LCASE_0127_out_0
);
W_48_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x50_out_12,
   I1 => x50_out_19,
   I2 => x50_out_21,
   I3 => W_48_3_i_10_n_0,
   I4 => W_48_3_i_11_n_0,
   O => W_48_3_i_2_n_0
);
W_48_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_48_3_i_11_n_0,
   I1 => x50_out_21,
   I2 => x50_out_19,
   I3 => x50_out_12,
   I4 => W_48_3_i_10_n_0,
   O => W_48_3_i_3_n_0
);
W_48_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_0127_out_1,
   I1 => x65_out_1,
   I2 => x92_out_1,
   I3 => x50_out_11,
   I4 => x50_out_18,
   I5 => x50_out_20,
   O => W_48_3_i_4_n_0
);
W_48_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x92_out_0,
   I1 => x65_out_0,
   I2 => x89_out_18,
   I3 => x89_out_7,
   I4 => x89_out_3,
   O => W_48_3_i_5_n_0
);
W_48_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_48_3_i_2_n_0,
   I1 => W_48_7_i_16_n_0,
   I2 => x50_out_13,
   I3 => x50_out_20,
   I4 => x50_out_22,
   I5 => W_48_7_i_17_n_0,
   O => W_48_3_i_6_n_0
);
W_48_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_48_3_i_10_n_0,
   I1 => SIGMA_LCASE_1131_out_0_2,
   I2 => x92_out_1,
   I3 => x65_out_1,
   I4 => SIGMA_LCASE_0127_out_1,
   I5 => SIGMA_LCASE_1131_out_1,
   O => W_48_3_i_7_n_0
);
W_48_3_i_8 : LUT5
  generic map(
   INIT => X"99969666"
  )
 port map (
   I0 => SIGMA_LCASE_1131_out_1,
   I1 => W_48_3_i_15_n_0,
   I2 => x92_out_0,
   I3 => SIGMA_LCASE_0127_out_0,
   I4 => x65_out_0,
   O => W_48_3_i_8_n_0
);
W_48_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_48_3_i_5_n_0,
   I1 => x50_out_10,
   I2 => x50_out_17,
   I3 => x50_out_19,
   O => W_48_3_i_9_n_0
);
W_48_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x92_out_6,
   I1 => x65_out_6,
   I2 => x89_out_24,
   I3 => x89_out_13,
   I4 => x89_out_9,
   O => W_48_7_i_10_n_0
);
W_48_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x65_out_5,
   I1 => x89_out_8,
   I2 => x89_out_12,
   I3 => x89_out_23,
   I4 => x92_out_5,
   O => W_48_7_i_11_n_0
);
W_48_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x92_out_5,
   I1 => x65_out_5,
   I2 => x89_out_23,
   I3 => x89_out_12,
   I4 => x89_out_8,
   O => W_48_7_i_12_n_0
);
W_48_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x65_out_4,
   I1 => x89_out_7,
   I2 => x89_out_11,
   I3 => x89_out_22,
   I4 => x92_out_4,
   O => W_48_7_i_13_n_0
);
W_48_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x92_out_4,
   I1 => x65_out_4,
   I2 => x89_out_22,
   I3 => x89_out_11,
   I4 => x89_out_7,
   O => W_48_7_i_14_n_0
);
W_48_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x65_out_3,
   I1 => x89_out_6,
   I2 => x89_out_10,
   I3 => x89_out_21,
   I4 => x92_out_3,
   O => W_48_7_i_15_n_0
);
W_48_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x92_out_3,
   I1 => x65_out_3,
   I2 => x89_out_21,
   I3 => x89_out_10,
   I4 => x89_out_6,
   O => W_48_7_i_16_n_0
);
W_48_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x65_out_2,
   I1 => x89_out_5,
   I2 => x89_out_9,
   I3 => x89_out_20,
   I4 => x92_out_2,
   O => W_48_7_i_17_n_0
);
W_48_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x50_out_16,
   I1 => x50_out_23,
   I2 => x50_out_25,
   I3 => W_48_7_i_10_n_0,
   I4 => W_48_7_i_11_n_0,
   O => W_48_7_i_2_n_0
);
W_48_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x50_out_15,
   I1 => x50_out_22,
   I2 => x50_out_24,
   I3 => W_48_7_i_12_n_0,
   I4 => W_48_7_i_13_n_0,
   O => W_48_7_i_3_n_0
);
W_48_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x50_out_14,
   I1 => x50_out_21,
   I2 => x50_out_23,
   I3 => W_48_7_i_14_n_0,
   I4 => W_48_7_i_15_n_0,
   O => W_48_7_i_4_n_0
);
W_48_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x50_out_13,
   I1 => x50_out_20,
   I2 => x50_out_22,
   I3 => W_48_7_i_16_n_0,
   I4 => W_48_7_i_17_n_0,
   O => W_48_7_i_5_n_0
);
W_48_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_48_7_i_2_n_0,
   I1 => W_48_11_i_16_n_0,
   I2 => x50_out_17,
   I3 => x50_out_24,
   I4 => x50_out_26,
   I5 => W_48_11_i_17_n_0,
   O => W_48_7_i_6_n_0
);
W_48_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_48_7_i_3_n_0,
   I1 => W_48_7_i_10_n_0,
   I2 => x50_out_16,
   I3 => x50_out_23,
   I4 => x50_out_25,
   I5 => W_48_7_i_11_n_0,
   O => W_48_7_i_7_n_0
);
W_48_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_48_7_i_4_n_0,
   I1 => W_48_7_i_12_n_0,
   I2 => x50_out_15,
   I3 => x50_out_22,
   I4 => x50_out_24,
   I5 => W_48_7_i_13_n_0,
   O => W_48_7_i_8_n_0
);
W_48_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_48_7_i_5_n_0,
   I1 => W_48_7_i_14_n_0,
   I2 => x50_out_14,
   I3 => x50_out_21,
   I4 => x50_out_23,
   I5 => W_48_7_i_15_n_0,
   O => W_48_7_i_9_n_0
);
W_49_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x89_out_10,
   I1 => x62_out_10,
   I2 => x86_out_28,
   I3 => x86_out_17,
   I4 => x86_out_13,
   O => W_49_11_i_10_n_0
);
W_49_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x62_out_9,
   I1 => x86_out_12,
   I2 => x86_out_16,
   I3 => x86_out_27,
   I4 => x89_out_9,
   O => W_49_11_i_11_n_0
);
W_49_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x89_out_9,
   I1 => x62_out_9,
   I2 => x86_out_27,
   I3 => x86_out_16,
   I4 => x86_out_12,
   O => W_49_11_i_12_n_0
);
W_49_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x62_out_8,
   I1 => x86_out_11,
   I2 => x86_out_15,
   I3 => x86_out_26,
   I4 => x89_out_8,
   O => W_49_11_i_13_n_0
);
W_49_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x89_out_8,
   I1 => x62_out_8,
   I2 => x86_out_26,
   I3 => x86_out_15,
   I4 => x86_out_11,
   O => W_49_11_i_14_n_0
);
W_49_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x62_out_7,
   I1 => x86_out_10,
   I2 => x86_out_14,
   I3 => x86_out_25,
   I4 => x89_out_7,
   O => W_49_11_i_15_n_0
);
W_49_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x89_out_7,
   I1 => x62_out_7,
   I2 => x86_out_25,
   I3 => x86_out_14,
   I4 => x86_out_10,
   O => W_49_11_i_16_n_0
);
W_49_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x62_out_6,
   I1 => x86_out_9,
   I2 => x86_out_13,
   I3 => x86_out_24,
   I4 => x89_out_6,
   O => W_49_11_i_17_n_0
);
W_49_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x47_out_20,
   I1 => x47_out_27,
   I2 => x47_out_29,
   I3 => W_49_11_i_10_n_0,
   I4 => W_49_11_i_11_n_0,
   O => W_49_11_i_2_n_0
);
W_49_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x47_out_19,
   I1 => x47_out_26,
   I2 => x47_out_28,
   I3 => W_49_11_i_12_n_0,
   I4 => W_49_11_i_13_n_0,
   O => W_49_11_i_3_n_0
);
W_49_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x47_out_18,
   I1 => x47_out_25,
   I2 => x47_out_27,
   I3 => W_49_11_i_14_n_0,
   I4 => W_49_11_i_15_n_0,
   O => W_49_11_i_4_n_0
);
W_49_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x47_out_17,
   I1 => x47_out_24,
   I2 => x47_out_26,
   I3 => W_49_11_i_16_n_0,
   I4 => W_49_11_i_17_n_0,
   O => W_49_11_i_5_n_0
);
W_49_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_49_11_i_2_n_0,
   I1 => W_49_15_i_16_n_0,
   I2 => x47_out_21,
   I3 => x47_out_28,
   I4 => x47_out_30,
   I5 => W_49_15_i_17_n_0,
   O => W_49_11_i_6_n_0
);
W_49_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_49_11_i_3_n_0,
   I1 => W_49_11_i_10_n_0,
   I2 => x47_out_20,
   I3 => x47_out_27,
   I4 => x47_out_29,
   I5 => W_49_11_i_11_n_0,
   O => W_49_11_i_7_n_0
);
W_49_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_49_11_i_4_n_0,
   I1 => W_49_11_i_12_n_0,
   I2 => x47_out_19,
   I3 => x47_out_26,
   I4 => x47_out_28,
   I5 => W_49_11_i_13_n_0,
   O => W_49_11_i_8_n_0
);
W_49_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_49_11_i_5_n_0,
   I1 => W_49_11_i_14_n_0,
   I2 => x47_out_18,
   I3 => x47_out_25,
   I4 => x47_out_27,
   I5 => W_49_11_i_15_n_0,
   O => W_49_11_i_9_n_0
);
W_49_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x89_out_14,
   I1 => x62_out_14,
   I2 => x86_out_0,
   I3 => x86_out_21,
   I4 => x86_out_17,
   O => W_49_15_i_10_n_0
);
W_49_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x62_out_13,
   I1 => x86_out_16,
   I2 => x86_out_20,
   I3 => x86_out_31,
   I4 => x89_out_13,
   O => W_49_15_i_11_n_0
);
W_49_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x89_out_13,
   I1 => x62_out_13,
   I2 => x86_out_31,
   I3 => x86_out_20,
   I4 => x86_out_16,
   O => W_49_15_i_12_n_0
);
W_49_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x62_out_12,
   I1 => x86_out_15,
   I2 => x86_out_19,
   I3 => x86_out_30,
   I4 => x89_out_12,
   O => W_49_15_i_13_n_0
);
W_49_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x89_out_12,
   I1 => x62_out_12,
   I2 => x86_out_30,
   I3 => x86_out_19,
   I4 => x86_out_15,
   O => W_49_15_i_14_n_0
);
W_49_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x62_out_11,
   I1 => x86_out_14,
   I2 => x86_out_18,
   I3 => x86_out_29,
   I4 => x89_out_11,
   O => W_49_15_i_15_n_0
);
W_49_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x89_out_11,
   I1 => x62_out_11,
   I2 => x86_out_29,
   I3 => x86_out_18,
   I4 => x86_out_14,
   O => W_49_15_i_16_n_0
);
W_49_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x62_out_10,
   I1 => x86_out_13,
   I2 => x86_out_17,
   I3 => x86_out_28,
   I4 => x89_out_10,
   O => W_49_15_i_17_n_0
);
W_49_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x47_out_24,
   I1 => x47_out_31,
   I2 => x47_out_1,
   I3 => W_49_15_i_10_n_0,
   I4 => W_49_15_i_11_n_0,
   O => W_49_15_i_2_n_0
);
W_49_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x47_out_23,
   I1 => x47_out_30,
   I2 => x47_out_0,
   I3 => W_49_15_i_12_n_0,
   I4 => W_49_15_i_13_n_0,
   O => W_49_15_i_3_n_0
);
W_49_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x47_out_22,
   I1 => x47_out_29,
   I2 => x47_out_31,
   I3 => W_49_15_i_14_n_0,
   I4 => W_49_15_i_15_n_0,
   O => W_49_15_i_4_n_0
);
W_49_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x47_out_21,
   I1 => x47_out_28,
   I2 => x47_out_30,
   I3 => W_49_15_i_16_n_0,
   I4 => W_49_15_i_17_n_0,
   O => W_49_15_i_5_n_0
);
W_49_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_49_15_i_2_n_0,
   I1 => W_49_19_i_16_n_0,
   I2 => x47_out_25,
   I3 => x47_out_0,
   I4 => x47_out_2,
   I5 => W_49_19_i_17_n_0,
   O => W_49_15_i_6_n_0
);
W_49_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_49_15_i_3_n_0,
   I1 => W_49_15_i_10_n_0,
   I2 => x47_out_24,
   I3 => x47_out_31,
   I4 => x47_out_1,
   I5 => W_49_15_i_11_n_0,
   O => W_49_15_i_7_n_0
);
W_49_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_49_15_i_4_n_0,
   I1 => W_49_15_i_12_n_0,
   I2 => x47_out_23,
   I3 => x47_out_30,
   I4 => x47_out_0,
   I5 => W_49_15_i_13_n_0,
   O => W_49_15_i_8_n_0
);
W_49_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_49_15_i_5_n_0,
   I1 => W_49_15_i_14_n_0,
   I2 => x47_out_22,
   I3 => x47_out_29,
   I4 => x47_out_31,
   I5 => W_49_15_i_15_n_0,
   O => W_49_15_i_9_n_0
);
W_49_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x89_out_18,
   I1 => x62_out_18,
   I2 => x86_out_4,
   I3 => x86_out_25,
   I4 => x86_out_21,
   O => W_49_19_i_10_n_0
);
W_49_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x62_out_17,
   I1 => x86_out_20,
   I2 => x86_out_24,
   I3 => x86_out_3,
   I4 => x89_out_17,
   O => W_49_19_i_11_n_0
);
W_49_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x89_out_17,
   I1 => x62_out_17,
   I2 => x86_out_3,
   I3 => x86_out_24,
   I4 => x86_out_20,
   O => W_49_19_i_12_n_0
);
W_49_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x62_out_16,
   I1 => x86_out_19,
   I2 => x86_out_23,
   I3 => x86_out_2,
   I4 => x89_out_16,
   O => W_49_19_i_13_n_0
);
W_49_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x89_out_16,
   I1 => x62_out_16,
   I2 => x86_out_2,
   I3 => x86_out_23,
   I4 => x86_out_19,
   O => W_49_19_i_14_n_0
);
W_49_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x62_out_15,
   I1 => x86_out_18,
   I2 => x86_out_22,
   I3 => x86_out_1,
   I4 => x89_out_15,
   O => W_49_19_i_15_n_0
);
W_49_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x89_out_15,
   I1 => x62_out_15,
   I2 => x86_out_1,
   I3 => x86_out_22,
   I4 => x86_out_18,
   O => W_49_19_i_16_n_0
);
W_49_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x62_out_14,
   I1 => x86_out_17,
   I2 => x86_out_21,
   I3 => x86_out_0,
   I4 => x89_out_14,
   O => W_49_19_i_17_n_0
);
W_49_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x47_out_28,
   I1 => x47_out_3,
   I2 => x47_out_5,
   I3 => W_49_19_i_10_n_0,
   I4 => W_49_19_i_11_n_0,
   O => W_49_19_i_2_n_0
);
W_49_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x47_out_27,
   I1 => x47_out_2,
   I2 => x47_out_4,
   I3 => W_49_19_i_12_n_0,
   I4 => W_49_19_i_13_n_0,
   O => W_49_19_i_3_n_0
);
W_49_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x47_out_26,
   I1 => x47_out_1,
   I2 => x47_out_3,
   I3 => W_49_19_i_14_n_0,
   I4 => W_49_19_i_15_n_0,
   O => W_49_19_i_4_n_0
);
W_49_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x47_out_25,
   I1 => x47_out_0,
   I2 => x47_out_2,
   I3 => W_49_19_i_16_n_0,
   I4 => W_49_19_i_17_n_0,
   O => W_49_19_i_5_n_0
);
W_49_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_49_19_i_2_n_0,
   I1 => W_49_23_i_16_n_0,
   I2 => x47_out_29,
   I3 => x47_out_4,
   I4 => x47_out_6,
   I5 => W_49_23_i_17_n_0,
   O => W_49_19_i_6_n_0
);
W_49_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_49_19_i_3_n_0,
   I1 => W_49_19_i_10_n_0,
   I2 => x47_out_28,
   I3 => x47_out_3,
   I4 => x47_out_5,
   I5 => W_49_19_i_11_n_0,
   O => W_49_19_i_7_n_0
);
W_49_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_49_19_i_4_n_0,
   I1 => W_49_19_i_12_n_0,
   I2 => x47_out_27,
   I3 => x47_out_2,
   I4 => x47_out_4,
   I5 => W_49_19_i_13_n_0,
   O => W_49_19_i_8_n_0
);
W_49_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_49_19_i_5_n_0,
   I1 => W_49_19_i_14_n_0,
   I2 => x47_out_26,
   I3 => x47_out_1,
   I4 => x47_out_3,
   I5 => W_49_19_i_15_n_0,
   O => W_49_19_i_9_n_0
);
W_49_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x89_out_22,
   I1 => x62_out_22,
   I2 => x86_out_8,
   I3 => x86_out_29,
   I4 => x86_out_25,
   O => W_49_23_i_10_n_0
);
W_49_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x62_out_21,
   I1 => x86_out_24,
   I2 => x86_out_28,
   I3 => x86_out_7,
   I4 => x89_out_21,
   O => W_49_23_i_11_n_0
);
W_49_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x89_out_21,
   I1 => x62_out_21,
   I2 => x86_out_7,
   I3 => x86_out_28,
   I4 => x86_out_24,
   O => W_49_23_i_12_n_0
);
W_49_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x62_out_20,
   I1 => x86_out_23,
   I2 => x86_out_27,
   I3 => x86_out_6,
   I4 => x89_out_20,
   O => W_49_23_i_13_n_0
);
W_49_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x89_out_20,
   I1 => x62_out_20,
   I2 => x86_out_6,
   I3 => x86_out_27,
   I4 => x86_out_23,
   O => W_49_23_i_14_n_0
);
W_49_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x62_out_19,
   I1 => x86_out_22,
   I2 => x86_out_26,
   I3 => x86_out_5,
   I4 => x89_out_19,
   O => W_49_23_i_15_n_0
);
W_49_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x89_out_19,
   I1 => x62_out_19,
   I2 => x86_out_5,
   I3 => x86_out_26,
   I4 => x86_out_22,
   O => W_49_23_i_16_n_0
);
W_49_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x62_out_18,
   I1 => x86_out_21,
   I2 => x86_out_25,
   I3 => x86_out_4,
   I4 => x89_out_18,
   O => W_49_23_i_17_n_0
);
W_49_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x47_out_7,
   I1 => x47_out_9,
   I2 => W_49_23_i_10_n_0,
   I3 => W_49_23_i_11_n_0,
   O => W_49_23_i_2_n_0
);
W_49_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x47_out_31,
   I1 => x47_out_6,
   I2 => x47_out_8,
   I3 => W_49_23_i_12_n_0,
   I4 => W_49_23_i_13_n_0,
   O => W_49_23_i_3_n_0
);
W_49_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x47_out_30,
   I1 => x47_out_5,
   I2 => x47_out_7,
   I3 => W_49_23_i_14_n_0,
   I4 => W_49_23_i_15_n_0,
   O => W_49_23_i_4_n_0
);
W_49_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x47_out_29,
   I1 => x47_out_4,
   I2 => x47_out_6,
   I3 => W_49_23_i_16_n_0,
   I4 => W_49_23_i_17_n_0,
   O => W_49_23_i_5_n_0
);
W_49_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x47_out_8,
   I1 => x47_out_10,
   I2 => W_49_27_i_16_n_0,
   I3 => W_49_27_i_17_n_0,
   I4 => W_49_23_i_2_n_0,
   O => W_49_23_i_6_n_0
);
W_49_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x47_out_7,
   I1 => x47_out_9,
   I2 => W_49_23_i_10_n_0,
   I3 => W_49_23_i_11_n_0,
   I4 => W_49_23_i_3_n_0,
   O => W_49_23_i_7_n_0
);
W_49_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_49_23_i_4_n_0,
   I1 => W_49_23_i_12_n_0,
   I2 => x47_out_31,
   I3 => x47_out_6,
   I4 => x47_out_8,
   I5 => W_49_23_i_13_n_0,
   O => W_49_23_i_8_n_0
);
W_49_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_49_23_i_5_n_0,
   I1 => W_49_23_i_14_n_0,
   I2 => x47_out_30,
   I3 => x47_out_5,
   I4 => x47_out_7,
   I5 => W_49_23_i_15_n_0,
   O => W_49_23_i_9_n_0
);
W_49_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x89_out_26,
   I1 => x62_out_26,
   I2 => x86_out_12,
   I3 => x86_out_1,
   I4 => x86_out_29,
   O => W_49_27_i_10_n_0
);
W_49_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x62_out_25,
   I1 => x86_out_28,
   I2 => x86_out_0,
   I3 => x86_out_11,
   I4 => x89_out_25,
   O => W_49_27_i_11_n_0
);
W_49_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x89_out_25,
   I1 => x62_out_25,
   I2 => x86_out_11,
   I3 => x86_out_0,
   I4 => x86_out_28,
   O => W_49_27_i_12_n_0
);
W_49_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x62_out_24,
   I1 => x86_out_27,
   I2 => x86_out_31,
   I3 => x86_out_10,
   I4 => x89_out_24,
   O => W_49_27_i_13_n_0
);
W_49_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x89_out_24,
   I1 => x62_out_24,
   I2 => x86_out_10,
   I3 => x86_out_31,
   I4 => x86_out_27,
   O => W_49_27_i_14_n_0
);
W_49_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x62_out_23,
   I1 => x86_out_26,
   I2 => x86_out_30,
   I3 => x86_out_9,
   I4 => x89_out_23,
   O => W_49_27_i_15_n_0
);
W_49_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x89_out_23,
   I1 => x62_out_23,
   I2 => x86_out_9,
   I3 => x86_out_30,
   I4 => x86_out_26,
   O => W_49_27_i_16_n_0
);
W_49_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x62_out_22,
   I1 => x86_out_25,
   I2 => x86_out_29,
   I3 => x86_out_8,
   I4 => x89_out_22,
   O => W_49_27_i_17_n_0
);
W_49_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x47_out_11,
   I1 => x47_out_13,
   I2 => W_49_27_i_10_n_0,
   I3 => W_49_27_i_11_n_0,
   O => W_49_27_i_2_n_0
);
W_49_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x47_out_10,
   I1 => x47_out_12,
   I2 => W_49_27_i_12_n_0,
   I3 => W_49_27_i_13_n_0,
   O => W_49_27_i_3_n_0
);
W_49_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x47_out_9,
   I1 => x47_out_11,
   I2 => W_49_27_i_14_n_0,
   I3 => W_49_27_i_15_n_0,
   O => W_49_27_i_4_n_0
);
W_49_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x47_out_8,
   I1 => x47_out_10,
   I2 => W_49_27_i_16_n_0,
   I3 => W_49_27_i_17_n_0,
   O => W_49_27_i_5_n_0
);
W_49_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x47_out_12,
   I1 => x47_out_14,
   I2 => W_49_31_i_13_n_0,
   I3 => W_49_31_i_14_n_0,
   I4 => W_49_27_i_2_n_0,
   O => W_49_27_i_6_n_0
);
W_49_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x47_out_11,
   I1 => x47_out_13,
   I2 => W_49_27_i_10_n_0,
   I3 => W_49_27_i_11_n_0,
   I4 => W_49_27_i_3_n_0,
   O => W_49_27_i_7_n_0
);
W_49_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x47_out_10,
   I1 => x47_out_12,
   I2 => W_49_27_i_12_n_0,
   I3 => W_49_27_i_13_n_0,
   I4 => W_49_27_i_4_n_0,
   O => W_49_27_i_8_n_0
);
W_49_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x47_out_9,
   I1 => x47_out_11,
   I2 => W_49_27_i_14_n_0,
   I3 => W_49_27_i_15_n_0,
   I4 => W_49_27_i_5_n_0,
   O => W_49_27_i_9_n_0
);
W_49_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x62_out_28,
   I1 => x86_out_31,
   I2 => x86_out_3,
   I3 => x86_out_14,
   I4 => x89_out_28,
   O => W_49_31_i_10_n_0
);
W_49_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x89_out_28,
   I1 => x62_out_28,
   I2 => x86_out_14,
   I3 => x86_out_3,
   I4 => x86_out_31,
   O => W_49_31_i_11_n_0
);
W_49_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x62_out_27,
   I1 => x86_out_30,
   I2 => x86_out_2,
   I3 => x86_out_13,
   I4 => x89_out_27,
   O => W_49_31_i_12_n_0
);
W_49_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x89_out_27,
   I1 => x62_out_27,
   I2 => x86_out_13,
   I3 => x86_out_2,
   I4 => x86_out_30,
   O => W_49_31_i_13_n_0
);
W_49_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x62_out_26,
   I1 => x86_out_29,
   I2 => x86_out_1,
   I3 => x86_out_12,
   I4 => x89_out_26,
   O => W_49_31_i_14_n_0
);
W_49_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x62_out_29,
   I1 => x86_out_4,
   I2 => x86_out_15,
   I3 => x89_out_29,
   O => W_49_31_i_15_n_0
);
W_49_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x47_out_17,
   I1 => x47_out_15,
   O => SIGMA_LCASE_1123_out_0_30
);
W_49_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => x86_out_6,
   I1 => x86_out_17,
   I2 => x62_out_31,
   I3 => x89_out_31,
   I4 => x47_out_16,
   I5 => x47_out_18,
   O => W_49_31_i_17_n_0
);
W_49_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x86_out_16,
   I1 => x86_out_5,
   O => SIGMA_LCASE_0119_out_30
);
W_49_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x89_out_30,
   I1 => x62_out_30,
   I2 => x86_out_16,
   I3 => x86_out_5,
   O => W_49_31_i_19_n_0
);
W_49_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x47_out_14,
   I1 => x47_out_16,
   I2 => W_49_31_i_9_n_0,
   I3 => W_49_31_i_10_n_0,
   O => W_49_31_i_2_n_0
);
W_49_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x47_out_13,
   I1 => x47_out_15,
   I2 => W_49_31_i_11_n_0,
   I3 => W_49_31_i_12_n_0,
   O => W_49_31_i_3_n_0
);
W_49_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x47_out_12,
   I1 => x47_out_14,
   I2 => W_49_31_i_13_n_0,
   I3 => W_49_31_i_14_n_0,
   O => W_49_31_i_4_n_0
);
W_49_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_49_31_i_15_n_0,
   I1 => SIGMA_LCASE_1123_out_0_30,
   I2 => W_49_31_i_17_n_0,
   I3 => x62_out_30,
   I4 => SIGMA_LCASE_0119_out_30,
   I5 => x89_out_30,
   O => W_49_31_i_5_n_0
);
W_49_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_49_31_i_2_n_0,
   I1 => W_49_31_i_19_n_0,
   I2 => x47_out_15,
   I3 => x47_out_17,
   I4 => W_49_31_i_15_n_0,
   O => W_49_31_i_6_n_0
);
W_49_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x47_out_14,
   I1 => x47_out_16,
   I2 => W_49_31_i_9_n_0,
   I3 => W_49_31_i_10_n_0,
   I4 => W_49_31_i_3_n_0,
   O => W_49_31_i_7_n_0
);
W_49_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x47_out_13,
   I1 => x47_out_15,
   I2 => W_49_31_i_11_n_0,
   I3 => W_49_31_i_12_n_0,
   I4 => W_49_31_i_4_n_0,
   O => W_49_31_i_8_n_0
);
W_49_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x89_out_29,
   I1 => x62_out_29,
   I2 => x86_out_15,
   I3 => x86_out_4,
   O => W_49_31_i_9_n_0
);
W_49_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x89_out_2,
   I1 => x62_out_2,
   I2 => x86_out_20,
   I3 => x86_out_9,
   I4 => x86_out_5,
   O => W_49_3_i_10_n_0
);
W_49_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x62_out_1,
   I1 => x86_out_4,
   I2 => x86_out_8,
   I3 => x86_out_19,
   I4 => x89_out_1,
   O => W_49_3_i_11_n_0
);
W_49_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x86_out_19,
   I1 => x86_out_8,
   I2 => x86_out_4,
   O => SIGMA_LCASE_0119_out_1
);
W_49_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x47_out_21,
   I1 => x47_out_19,
   I2 => x47_out_12,
   O => SIGMA_LCASE_1123_out_0_2
);
W_49_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x47_out_20,
   I1 => x47_out_18,
   I2 => x47_out_11,
   O => SIGMA_LCASE_1123_out_1
);
W_49_3_i_15 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x89_out_1,
   I1 => x62_out_1,
   I2 => x86_out_19,
   I3 => x86_out_8,
   I4 => x86_out_4,
   O => W_49_3_i_15_n_0
);
W_49_3_i_16 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x86_out_18,
   I1 => x86_out_7,
   I2 => x86_out_3,
   O => SIGMA_LCASE_0119_out_0
);
W_49_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x47_out_12,
   I1 => x47_out_19,
   I2 => x47_out_21,
   I3 => W_49_3_i_10_n_0,
   I4 => W_49_3_i_11_n_0,
   O => W_49_3_i_2_n_0
);
W_49_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_49_3_i_11_n_0,
   I1 => x47_out_21,
   I2 => x47_out_19,
   I3 => x47_out_12,
   I4 => W_49_3_i_10_n_0,
   O => W_49_3_i_3_n_0
);
W_49_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_0119_out_1,
   I1 => x62_out_1,
   I2 => x89_out_1,
   I3 => x47_out_11,
   I4 => x47_out_18,
   I5 => x47_out_20,
   O => W_49_3_i_4_n_0
);
W_49_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x89_out_0,
   I1 => x62_out_0,
   I2 => x86_out_18,
   I3 => x86_out_7,
   I4 => x86_out_3,
   O => W_49_3_i_5_n_0
);
W_49_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_49_3_i_2_n_0,
   I1 => W_49_7_i_16_n_0,
   I2 => x47_out_13,
   I3 => x47_out_20,
   I4 => x47_out_22,
   I5 => W_49_7_i_17_n_0,
   O => W_49_3_i_6_n_0
);
W_49_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_49_3_i_10_n_0,
   I1 => SIGMA_LCASE_1123_out_0_2,
   I2 => x89_out_1,
   I3 => x62_out_1,
   I4 => SIGMA_LCASE_0119_out_1,
   I5 => SIGMA_LCASE_1123_out_1,
   O => W_49_3_i_7_n_0
);
W_49_3_i_8 : LUT5
  generic map(
   INIT => X"99969666"
  )
 port map (
   I0 => SIGMA_LCASE_1123_out_1,
   I1 => W_49_3_i_15_n_0,
   I2 => x89_out_0,
   I3 => SIGMA_LCASE_0119_out_0,
   I4 => x62_out_0,
   O => W_49_3_i_8_n_0
);
W_49_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_49_3_i_5_n_0,
   I1 => x47_out_10,
   I2 => x47_out_17,
   I3 => x47_out_19,
   O => W_49_3_i_9_n_0
);
W_49_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x89_out_6,
   I1 => x62_out_6,
   I2 => x86_out_24,
   I3 => x86_out_13,
   I4 => x86_out_9,
   O => W_49_7_i_10_n_0
);
W_49_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x62_out_5,
   I1 => x86_out_8,
   I2 => x86_out_12,
   I3 => x86_out_23,
   I4 => x89_out_5,
   O => W_49_7_i_11_n_0
);
W_49_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x89_out_5,
   I1 => x62_out_5,
   I2 => x86_out_23,
   I3 => x86_out_12,
   I4 => x86_out_8,
   O => W_49_7_i_12_n_0
);
W_49_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x62_out_4,
   I1 => x86_out_7,
   I2 => x86_out_11,
   I3 => x86_out_22,
   I4 => x89_out_4,
   O => W_49_7_i_13_n_0
);
W_49_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x89_out_4,
   I1 => x62_out_4,
   I2 => x86_out_22,
   I3 => x86_out_11,
   I4 => x86_out_7,
   O => W_49_7_i_14_n_0
);
W_49_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x62_out_3,
   I1 => x86_out_6,
   I2 => x86_out_10,
   I3 => x86_out_21,
   I4 => x89_out_3,
   O => W_49_7_i_15_n_0
);
W_49_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x89_out_3,
   I1 => x62_out_3,
   I2 => x86_out_21,
   I3 => x86_out_10,
   I4 => x86_out_6,
   O => W_49_7_i_16_n_0
);
W_49_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x62_out_2,
   I1 => x86_out_5,
   I2 => x86_out_9,
   I3 => x86_out_20,
   I4 => x89_out_2,
   O => W_49_7_i_17_n_0
);
W_49_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x47_out_16,
   I1 => x47_out_23,
   I2 => x47_out_25,
   I3 => W_49_7_i_10_n_0,
   I4 => W_49_7_i_11_n_0,
   O => W_49_7_i_2_n_0
);
W_49_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x47_out_15,
   I1 => x47_out_22,
   I2 => x47_out_24,
   I3 => W_49_7_i_12_n_0,
   I4 => W_49_7_i_13_n_0,
   O => W_49_7_i_3_n_0
);
W_49_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x47_out_14,
   I1 => x47_out_21,
   I2 => x47_out_23,
   I3 => W_49_7_i_14_n_0,
   I4 => W_49_7_i_15_n_0,
   O => W_49_7_i_4_n_0
);
W_49_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x47_out_13,
   I1 => x47_out_20,
   I2 => x47_out_22,
   I3 => W_49_7_i_16_n_0,
   I4 => W_49_7_i_17_n_0,
   O => W_49_7_i_5_n_0
);
W_49_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_49_7_i_2_n_0,
   I1 => W_49_11_i_16_n_0,
   I2 => x47_out_17,
   I3 => x47_out_24,
   I4 => x47_out_26,
   I5 => W_49_11_i_17_n_0,
   O => W_49_7_i_6_n_0
);
W_49_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_49_7_i_3_n_0,
   I1 => W_49_7_i_10_n_0,
   I2 => x47_out_16,
   I3 => x47_out_23,
   I4 => x47_out_25,
   I5 => W_49_7_i_11_n_0,
   O => W_49_7_i_7_n_0
);
W_49_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_49_7_i_4_n_0,
   I1 => W_49_7_i_12_n_0,
   I2 => x47_out_15,
   I3 => x47_out_22,
   I4 => x47_out_24,
   I5 => W_49_7_i_13_n_0,
   O => W_49_7_i_8_n_0
);
W_49_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_49_7_i_5_n_0,
   I1 => W_49_7_i_14_n_0,
   I2 => x47_out_14,
   I3 => x47_out_21,
   I4 => x47_out_23,
   I5 => W_49_7_i_15_n_0,
   O => W_49_7_i_9_n_0
);
W_50_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x86_out_10,
   I1 => x59_out_10,
   I2 => x83_out_28,
   I3 => x83_out_17,
   I4 => x83_out_13,
   O => W_50_11_i_10_n_0
);
W_50_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x59_out_9,
   I1 => x83_out_12,
   I2 => x83_out_16,
   I3 => x83_out_27,
   I4 => x86_out_9,
   O => W_50_11_i_11_n_0
);
W_50_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x86_out_9,
   I1 => x59_out_9,
   I2 => x83_out_27,
   I3 => x83_out_16,
   I4 => x83_out_12,
   O => W_50_11_i_12_n_0
);
W_50_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x59_out_8,
   I1 => x83_out_11,
   I2 => x83_out_15,
   I3 => x83_out_26,
   I4 => x86_out_8,
   O => W_50_11_i_13_n_0
);
W_50_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x86_out_8,
   I1 => x59_out_8,
   I2 => x83_out_26,
   I3 => x83_out_15,
   I4 => x83_out_11,
   O => W_50_11_i_14_n_0
);
W_50_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x59_out_7,
   I1 => x83_out_10,
   I2 => x83_out_14,
   I3 => x83_out_25,
   I4 => x86_out_7,
   O => W_50_11_i_15_n_0
);
W_50_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x86_out_7,
   I1 => x59_out_7,
   I2 => x83_out_25,
   I3 => x83_out_14,
   I4 => x83_out_10,
   O => W_50_11_i_16_n_0
);
W_50_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x59_out_6,
   I1 => x83_out_9,
   I2 => x83_out_13,
   I3 => x83_out_24,
   I4 => x86_out_6,
   O => W_50_11_i_17_n_0
);
W_50_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x44_out_20,
   I1 => x44_out_27,
   I2 => x44_out_29,
   I3 => W_50_11_i_10_n_0,
   I4 => W_50_11_i_11_n_0,
   O => W_50_11_i_2_n_0
);
W_50_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x44_out_19,
   I1 => x44_out_26,
   I2 => x44_out_28,
   I3 => W_50_11_i_12_n_0,
   I4 => W_50_11_i_13_n_0,
   O => W_50_11_i_3_n_0
);
W_50_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x44_out_18,
   I1 => x44_out_25,
   I2 => x44_out_27,
   I3 => W_50_11_i_14_n_0,
   I4 => W_50_11_i_15_n_0,
   O => W_50_11_i_4_n_0
);
W_50_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x44_out_17,
   I1 => x44_out_24,
   I2 => x44_out_26,
   I3 => W_50_11_i_16_n_0,
   I4 => W_50_11_i_17_n_0,
   O => W_50_11_i_5_n_0
);
W_50_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_50_11_i_2_n_0,
   I1 => W_50_15_i_16_n_0,
   I2 => x44_out_21,
   I3 => x44_out_28,
   I4 => x44_out_30,
   I5 => W_50_15_i_17_n_0,
   O => W_50_11_i_6_n_0
);
W_50_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_50_11_i_3_n_0,
   I1 => W_50_11_i_10_n_0,
   I2 => x44_out_20,
   I3 => x44_out_27,
   I4 => x44_out_29,
   I5 => W_50_11_i_11_n_0,
   O => W_50_11_i_7_n_0
);
W_50_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_50_11_i_4_n_0,
   I1 => W_50_11_i_12_n_0,
   I2 => x44_out_19,
   I3 => x44_out_26,
   I4 => x44_out_28,
   I5 => W_50_11_i_13_n_0,
   O => W_50_11_i_8_n_0
);
W_50_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_50_11_i_5_n_0,
   I1 => W_50_11_i_14_n_0,
   I2 => x44_out_18,
   I3 => x44_out_25,
   I4 => x44_out_27,
   I5 => W_50_11_i_15_n_0,
   O => W_50_11_i_9_n_0
);
W_50_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x86_out_14,
   I1 => x59_out_14,
   I2 => x83_out_0,
   I3 => x83_out_21,
   I4 => x83_out_17,
   O => W_50_15_i_10_n_0
);
W_50_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x59_out_13,
   I1 => x83_out_16,
   I2 => x83_out_20,
   I3 => x83_out_31,
   I4 => x86_out_13,
   O => W_50_15_i_11_n_0
);
W_50_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x86_out_13,
   I1 => x59_out_13,
   I2 => x83_out_31,
   I3 => x83_out_20,
   I4 => x83_out_16,
   O => W_50_15_i_12_n_0
);
W_50_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x59_out_12,
   I1 => x83_out_15,
   I2 => x83_out_19,
   I3 => x83_out_30,
   I4 => x86_out_12,
   O => W_50_15_i_13_n_0
);
W_50_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x86_out_12,
   I1 => x59_out_12,
   I2 => x83_out_30,
   I3 => x83_out_19,
   I4 => x83_out_15,
   O => W_50_15_i_14_n_0
);
W_50_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x59_out_11,
   I1 => x83_out_14,
   I2 => x83_out_18,
   I3 => x83_out_29,
   I4 => x86_out_11,
   O => W_50_15_i_15_n_0
);
W_50_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x86_out_11,
   I1 => x59_out_11,
   I2 => x83_out_29,
   I3 => x83_out_18,
   I4 => x83_out_14,
   O => W_50_15_i_16_n_0
);
W_50_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x59_out_10,
   I1 => x83_out_13,
   I2 => x83_out_17,
   I3 => x83_out_28,
   I4 => x86_out_10,
   O => W_50_15_i_17_n_0
);
W_50_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x44_out_24,
   I1 => x44_out_31,
   I2 => x44_out_1,
   I3 => W_50_15_i_10_n_0,
   I4 => W_50_15_i_11_n_0,
   O => W_50_15_i_2_n_0
);
W_50_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x44_out_23,
   I1 => x44_out_30,
   I2 => x44_out_0,
   I3 => W_50_15_i_12_n_0,
   I4 => W_50_15_i_13_n_0,
   O => W_50_15_i_3_n_0
);
W_50_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x44_out_22,
   I1 => x44_out_29,
   I2 => x44_out_31,
   I3 => W_50_15_i_14_n_0,
   I4 => W_50_15_i_15_n_0,
   O => W_50_15_i_4_n_0
);
W_50_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x44_out_21,
   I1 => x44_out_28,
   I2 => x44_out_30,
   I3 => W_50_15_i_16_n_0,
   I4 => W_50_15_i_17_n_0,
   O => W_50_15_i_5_n_0
);
W_50_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_50_15_i_2_n_0,
   I1 => W_50_19_i_16_n_0,
   I2 => x44_out_25,
   I3 => x44_out_0,
   I4 => x44_out_2,
   I5 => W_50_19_i_17_n_0,
   O => W_50_15_i_6_n_0
);
W_50_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_50_15_i_3_n_0,
   I1 => W_50_15_i_10_n_0,
   I2 => x44_out_24,
   I3 => x44_out_31,
   I4 => x44_out_1,
   I5 => W_50_15_i_11_n_0,
   O => W_50_15_i_7_n_0
);
W_50_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_50_15_i_4_n_0,
   I1 => W_50_15_i_12_n_0,
   I2 => x44_out_23,
   I3 => x44_out_30,
   I4 => x44_out_0,
   I5 => W_50_15_i_13_n_0,
   O => W_50_15_i_8_n_0
);
W_50_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_50_15_i_5_n_0,
   I1 => W_50_15_i_14_n_0,
   I2 => x44_out_22,
   I3 => x44_out_29,
   I4 => x44_out_31,
   I5 => W_50_15_i_15_n_0,
   O => W_50_15_i_9_n_0
);
W_50_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x86_out_18,
   I1 => x59_out_18,
   I2 => x83_out_4,
   I3 => x83_out_25,
   I4 => x83_out_21,
   O => W_50_19_i_10_n_0
);
W_50_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x59_out_17,
   I1 => x83_out_20,
   I2 => x83_out_24,
   I3 => x83_out_3,
   I4 => x86_out_17,
   O => W_50_19_i_11_n_0
);
W_50_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x86_out_17,
   I1 => x59_out_17,
   I2 => x83_out_3,
   I3 => x83_out_24,
   I4 => x83_out_20,
   O => W_50_19_i_12_n_0
);
W_50_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x59_out_16,
   I1 => x83_out_19,
   I2 => x83_out_23,
   I3 => x83_out_2,
   I4 => x86_out_16,
   O => W_50_19_i_13_n_0
);
W_50_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x86_out_16,
   I1 => x59_out_16,
   I2 => x83_out_2,
   I3 => x83_out_23,
   I4 => x83_out_19,
   O => W_50_19_i_14_n_0
);
W_50_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x59_out_15,
   I1 => x83_out_18,
   I2 => x83_out_22,
   I3 => x83_out_1,
   I4 => x86_out_15,
   O => W_50_19_i_15_n_0
);
W_50_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x86_out_15,
   I1 => x59_out_15,
   I2 => x83_out_1,
   I3 => x83_out_22,
   I4 => x83_out_18,
   O => W_50_19_i_16_n_0
);
W_50_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x59_out_14,
   I1 => x83_out_17,
   I2 => x83_out_21,
   I3 => x83_out_0,
   I4 => x86_out_14,
   O => W_50_19_i_17_n_0
);
W_50_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x44_out_28,
   I1 => x44_out_3,
   I2 => x44_out_5,
   I3 => W_50_19_i_10_n_0,
   I4 => W_50_19_i_11_n_0,
   O => W_50_19_i_2_n_0
);
W_50_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x44_out_27,
   I1 => x44_out_2,
   I2 => x44_out_4,
   I3 => W_50_19_i_12_n_0,
   I4 => W_50_19_i_13_n_0,
   O => W_50_19_i_3_n_0
);
W_50_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x44_out_26,
   I1 => x44_out_1,
   I2 => x44_out_3,
   I3 => W_50_19_i_14_n_0,
   I4 => W_50_19_i_15_n_0,
   O => W_50_19_i_4_n_0
);
W_50_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x44_out_25,
   I1 => x44_out_0,
   I2 => x44_out_2,
   I3 => W_50_19_i_16_n_0,
   I4 => W_50_19_i_17_n_0,
   O => W_50_19_i_5_n_0
);
W_50_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_50_19_i_2_n_0,
   I1 => W_50_23_i_16_n_0,
   I2 => x44_out_29,
   I3 => x44_out_4,
   I4 => x44_out_6,
   I5 => W_50_23_i_17_n_0,
   O => W_50_19_i_6_n_0
);
W_50_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_50_19_i_3_n_0,
   I1 => W_50_19_i_10_n_0,
   I2 => x44_out_28,
   I3 => x44_out_3,
   I4 => x44_out_5,
   I5 => W_50_19_i_11_n_0,
   O => W_50_19_i_7_n_0
);
W_50_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_50_19_i_4_n_0,
   I1 => W_50_19_i_12_n_0,
   I2 => x44_out_27,
   I3 => x44_out_2,
   I4 => x44_out_4,
   I5 => W_50_19_i_13_n_0,
   O => W_50_19_i_8_n_0
);
W_50_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_50_19_i_5_n_0,
   I1 => W_50_19_i_14_n_0,
   I2 => x44_out_26,
   I3 => x44_out_1,
   I4 => x44_out_3,
   I5 => W_50_19_i_15_n_0,
   O => W_50_19_i_9_n_0
);
W_50_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x86_out_22,
   I1 => x59_out_22,
   I2 => x83_out_8,
   I3 => x83_out_29,
   I4 => x83_out_25,
   O => W_50_23_i_10_n_0
);
W_50_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x59_out_21,
   I1 => x83_out_24,
   I2 => x83_out_28,
   I3 => x83_out_7,
   I4 => x86_out_21,
   O => W_50_23_i_11_n_0
);
W_50_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x86_out_21,
   I1 => x59_out_21,
   I2 => x83_out_7,
   I3 => x83_out_28,
   I4 => x83_out_24,
   O => W_50_23_i_12_n_0
);
W_50_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x59_out_20,
   I1 => x83_out_23,
   I2 => x83_out_27,
   I3 => x83_out_6,
   I4 => x86_out_20,
   O => W_50_23_i_13_n_0
);
W_50_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x86_out_20,
   I1 => x59_out_20,
   I2 => x83_out_6,
   I3 => x83_out_27,
   I4 => x83_out_23,
   O => W_50_23_i_14_n_0
);
W_50_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x59_out_19,
   I1 => x83_out_22,
   I2 => x83_out_26,
   I3 => x83_out_5,
   I4 => x86_out_19,
   O => W_50_23_i_15_n_0
);
W_50_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x86_out_19,
   I1 => x59_out_19,
   I2 => x83_out_5,
   I3 => x83_out_26,
   I4 => x83_out_22,
   O => W_50_23_i_16_n_0
);
W_50_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x59_out_18,
   I1 => x83_out_21,
   I2 => x83_out_25,
   I3 => x83_out_4,
   I4 => x86_out_18,
   O => W_50_23_i_17_n_0
);
W_50_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x44_out_7,
   I1 => x44_out_9,
   I2 => W_50_23_i_10_n_0,
   I3 => W_50_23_i_11_n_0,
   O => W_50_23_i_2_n_0
);
W_50_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x44_out_31,
   I1 => x44_out_6,
   I2 => x44_out_8,
   I3 => W_50_23_i_12_n_0,
   I4 => W_50_23_i_13_n_0,
   O => W_50_23_i_3_n_0
);
W_50_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x44_out_30,
   I1 => x44_out_5,
   I2 => x44_out_7,
   I3 => W_50_23_i_14_n_0,
   I4 => W_50_23_i_15_n_0,
   O => W_50_23_i_4_n_0
);
W_50_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x44_out_29,
   I1 => x44_out_4,
   I2 => x44_out_6,
   I3 => W_50_23_i_16_n_0,
   I4 => W_50_23_i_17_n_0,
   O => W_50_23_i_5_n_0
);
W_50_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x44_out_8,
   I1 => x44_out_10,
   I2 => W_50_27_i_16_n_0,
   I3 => W_50_27_i_17_n_0,
   I4 => W_50_23_i_2_n_0,
   O => W_50_23_i_6_n_0
);
W_50_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x44_out_7,
   I1 => x44_out_9,
   I2 => W_50_23_i_10_n_0,
   I3 => W_50_23_i_11_n_0,
   I4 => W_50_23_i_3_n_0,
   O => W_50_23_i_7_n_0
);
W_50_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_50_23_i_4_n_0,
   I1 => W_50_23_i_12_n_0,
   I2 => x44_out_31,
   I3 => x44_out_6,
   I4 => x44_out_8,
   I5 => W_50_23_i_13_n_0,
   O => W_50_23_i_8_n_0
);
W_50_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_50_23_i_5_n_0,
   I1 => W_50_23_i_14_n_0,
   I2 => x44_out_30,
   I3 => x44_out_5,
   I4 => x44_out_7,
   I5 => W_50_23_i_15_n_0,
   O => W_50_23_i_9_n_0
);
W_50_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x86_out_26,
   I1 => x59_out_26,
   I2 => x83_out_12,
   I3 => x83_out_1,
   I4 => x83_out_29,
   O => W_50_27_i_10_n_0
);
W_50_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x59_out_25,
   I1 => x83_out_28,
   I2 => x83_out_0,
   I3 => x83_out_11,
   I4 => x86_out_25,
   O => W_50_27_i_11_n_0
);
W_50_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x86_out_25,
   I1 => x59_out_25,
   I2 => x83_out_11,
   I3 => x83_out_0,
   I4 => x83_out_28,
   O => W_50_27_i_12_n_0
);
W_50_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x59_out_24,
   I1 => x83_out_27,
   I2 => x83_out_31,
   I3 => x83_out_10,
   I4 => x86_out_24,
   O => W_50_27_i_13_n_0
);
W_50_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x86_out_24,
   I1 => x59_out_24,
   I2 => x83_out_10,
   I3 => x83_out_31,
   I4 => x83_out_27,
   O => W_50_27_i_14_n_0
);
W_50_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x59_out_23,
   I1 => x83_out_26,
   I2 => x83_out_30,
   I3 => x83_out_9,
   I4 => x86_out_23,
   O => W_50_27_i_15_n_0
);
W_50_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x86_out_23,
   I1 => x59_out_23,
   I2 => x83_out_9,
   I3 => x83_out_30,
   I4 => x83_out_26,
   O => W_50_27_i_16_n_0
);
W_50_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x59_out_22,
   I1 => x83_out_25,
   I2 => x83_out_29,
   I3 => x83_out_8,
   I4 => x86_out_22,
   O => W_50_27_i_17_n_0
);
W_50_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x44_out_11,
   I1 => x44_out_13,
   I2 => W_50_27_i_10_n_0,
   I3 => W_50_27_i_11_n_0,
   O => W_50_27_i_2_n_0
);
W_50_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x44_out_10,
   I1 => x44_out_12,
   I2 => W_50_27_i_12_n_0,
   I3 => W_50_27_i_13_n_0,
   O => W_50_27_i_3_n_0
);
W_50_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x44_out_9,
   I1 => x44_out_11,
   I2 => W_50_27_i_14_n_0,
   I3 => W_50_27_i_15_n_0,
   O => W_50_27_i_4_n_0
);
W_50_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x44_out_8,
   I1 => x44_out_10,
   I2 => W_50_27_i_16_n_0,
   I3 => W_50_27_i_17_n_0,
   O => W_50_27_i_5_n_0
);
W_50_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x44_out_12,
   I1 => x44_out_14,
   I2 => W_50_31_i_13_n_0,
   I3 => W_50_31_i_14_n_0,
   I4 => W_50_27_i_2_n_0,
   O => W_50_27_i_6_n_0
);
W_50_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x44_out_11,
   I1 => x44_out_13,
   I2 => W_50_27_i_10_n_0,
   I3 => W_50_27_i_11_n_0,
   I4 => W_50_27_i_3_n_0,
   O => W_50_27_i_7_n_0
);
W_50_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x44_out_10,
   I1 => x44_out_12,
   I2 => W_50_27_i_12_n_0,
   I3 => W_50_27_i_13_n_0,
   I4 => W_50_27_i_4_n_0,
   O => W_50_27_i_8_n_0
);
W_50_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x44_out_9,
   I1 => x44_out_11,
   I2 => W_50_27_i_14_n_0,
   I3 => W_50_27_i_15_n_0,
   I4 => W_50_27_i_5_n_0,
   O => W_50_27_i_9_n_0
);
W_50_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x59_out_28,
   I1 => x83_out_31,
   I2 => x83_out_3,
   I3 => x83_out_14,
   I4 => x86_out_28,
   O => W_50_31_i_10_n_0
);
W_50_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x86_out_28,
   I1 => x59_out_28,
   I2 => x83_out_14,
   I3 => x83_out_3,
   I4 => x83_out_31,
   O => W_50_31_i_11_n_0
);
W_50_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x59_out_27,
   I1 => x83_out_30,
   I2 => x83_out_2,
   I3 => x83_out_13,
   I4 => x86_out_27,
   O => W_50_31_i_12_n_0
);
W_50_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x86_out_27,
   I1 => x59_out_27,
   I2 => x83_out_13,
   I3 => x83_out_2,
   I4 => x83_out_30,
   O => W_50_31_i_13_n_0
);
W_50_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x59_out_26,
   I1 => x83_out_29,
   I2 => x83_out_1,
   I3 => x83_out_12,
   I4 => x86_out_26,
   O => W_50_31_i_14_n_0
);
W_50_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x59_out_29,
   I1 => x83_out_4,
   I2 => x83_out_15,
   I3 => x86_out_29,
   O => W_50_31_i_15_n_0
);
W_50_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x44_out_17,
   I1 => x44_out_15,
   O => SIGMA_LCASE_1115_out_0_30
);
W_50_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => x83_out_6,
   I1 => x83_out_17,
   I2 => x59_out_31,
   I3 => x86_out_31,
   I4 => x44_out_16,
   I5 => x44_out_18,
   O => W_50_31_i_17_n_0
);
W_50_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x83_out_16,
   I1 => x83_out_5,
   O => SIGMA_LCASE_0111_out_30
);
W_50_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x86_out_30,
   I1 => x59_out_30,
   I2 => x83_out_16,
   I3 => x83_out_5,
   O => W_50_31_i_19_n_0
);
W_50_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x44_out_14,
   I1 => x44_out_16,
   I2 => W_50_31_i_9_n_0,
   I3 => W_50_31_i_10_n_0,
   O => W_50_31_i_2_n_0
);
W_50_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x44_out_13,
   I1 => x44_out_15,
   I2 => W_50_31_i_11_n_0,
   I3 => W_50_31_i_12_n_0,
   O => W_50_31_i_3_n_0
);
W_50_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x44_out_12,
   I1 => x44_out_14,
   I2 => W_50_31_i_13_n_0,
   I3 => W_50_31_i_14_n_0,
   O => W_50_31_i_4_n_0
);
W_50_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_50_31_i_15_n_0,
   I1 => SIGMA_LCASE_1115_out_0_30,
   I2 => W_50_31_i_17_n_0,
   I3 => x59_out_30,
   I4 => SIGMA_LCASE_0111_out_30,
   I5 => x86_out_30,
   O => W_50_31_i_5_n_0
);
W_50_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_50_31_i_2_n_0,
   I1 => W_50_31_i_19_n_0,
   I2 => x44_out_15,
   I3 => x44_out_17,
   I4 => W_50_31_i_15_n_0,
   O => W_50_31_i_6_n_0
);
W_50_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x44_out_14,
   I1 => x44_out_16,
   I2 => W_50_31_i_9_n_0,
   I3 => W_50_31_i_10_n_0,
   I4 => W_50_31_i_3_n_0,
   O => W_50_31_i_7_n_0
);
W_50_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x44_out_13,
   I1 => x44_out_15,
   I2 => W_50_31_i_11_n_0,
   I3 => W_50_31_i_12_n_0,
   I4 => W_50_31_i_4_n_0,
   O => W_50_31_i_8_n_0
);
W_50_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x86_out_29,
   I1 => x59_out_29,
   I2 => x83_out_15,
   I3 => x83_out_4,
   O => W_50_31_i_9_n_0
);
W_50_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x86_out_2,
   I1 => x59_out_2,
   I2 => x83_out_20,
   I3 => x83_out_9,
   I4 => x83_out_5,
   O => W_50_3_i_10_n_0
);
W_50_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x59_out_1,
   I1 => x83_out_4,
   I2 => x83_out_8,
   I3 => x83_out_19,
   I4 => x86_out_1,
   O => W_50_3_i_11_n_0
);
W_50_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x83_out_19,
   I1 => x83_out_8,
   I2 => x83_out_4,
   O => SIGMA_LCASE_0111_out_1
);
W_50_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x44_out_21,
   I1 => x44_out_19,
   I2 => x44_out_12,
   O => SIGMA_LCASE_1115_out_0_2
);
W_50_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x44_out_20,
   I1 => x44_out_18,
   I2 => x44_out_11,
   O => SIGMA_LCASE_1115_out_1
);
W_50_3_i_15 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x86_out_1,
   I1 => x59_out_1,
   I2 => x83_out_19,
   I3 => x83_out_8,
   I4 => x83_out_4,
   O => W_50_3_i_15_n_0
);
W_50_3_i_16 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x83_out_18,
   I1 => x83_out_7,
   I2 => x83_out_3,
   O => SIGMA_LCASE_0111_out_0
);
W_50_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x44_out_12,
   I1 => x44_out_19,
   I2 => x44_out_21,
   I3 => W_50_3_i_10_n_0,
   I4 => W_50_3_i_11_n_0,
   O => W_50_3_i_2_n_0
);
W_50_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_50_3_i_11_n_0,
   I1 => x44_out_21,
   I2 => x44_out_19,
   I3 => x44_out_12,
   I4 => W_50_3_i_10_n_0,
   O => W_50_3_i_3_n_0
);
W_50_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_0111_out_1,
   I1 => x59_out_1,
   I2 => x86_out_1,
   I3 => x44_out_11,
   I4 => x44_out_18,
   I5 => x44_out_20,
   O => W_50_3_i_4_n_0
);
W_50_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x86_out_0,
   I1 => x59_out_0,
   I2 => x83_out_18,
   I3 => x83_out_7,
   I4 => x83_out_3,
   O => W_50_3_i_5_n_0
);
W_50_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_50_3_i_2_n_0,
   I1 => W_50_7_i_16_n_0,
   I2 => x44_out_13,
   I3 => x44_out_20,
   I4 => x44_out_22,
   I5 => W_50_7_i_17_n_0,
   O => W_50_3_i_6_n_0
);
W_50_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_50_3_i_10_n_0,
   I1 => SIGMA_LCASE_1115_out_0_2,
   I2 => x86_out_1,
   I3 => x59_out_1,
   I4 => SIGMA_LCASE_0111_out_1,
   I5 => SIGMA_LCASE_1115_out_1,
   O => W_50_3_i_7_n_0
);
W_50_3_i_8 : LUT5
  generic map(
   INIT => X"99969666"
  )
 port map (
   I0 => SIGMA_LCASE_1115_out_1,
   I1 => W_50_3_i_15_n_0,
   I2 => x86_out_0,
   I3 => SIGMA_LCASE_0111_out_0,
   I4 => x59_out_0,
   O => W_50_3_i_8_n_0
);
W_50_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_50_3_i_5_n_0,
   I1 => x44_out_10,
   I2 => x44_out_17,
   I3 => x44_out_19,
   O => W_50_3_i_9_n_0
);
W_50_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x86_out_6,
   I1 => x59_out_6,
   I2 => x83_out_24,
   I3 => x83_out_13,
   I4 => x83_out_9,
   O => W_50_7_i_10_n_0
);
W_50_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x59_out_5,
   I1 => x83_out_8,
   I2 => x83_out_12,
   I3 => x83_out_23,
   I4 => x86_out_5,
   O => W_50_7_i_11_n_0
);
W_50_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x86_out_5,
   I1 => x59_out_5,
   I2 => x83_out_23,
   I3 => x83_out_12,
   I4 => x83_out_8,
   O => W_50_7_i_12_n_0
);
W_50_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x59_out_4,
   I1 => x83_out_7,
   I2 => x83_out_11,
   I3 => x83_out_22,
   I4 => x86_out_4,
   O => W_50_7_i_13_n_0
);
W_50_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x86_out_4,
   I1 => x59_out_4,
   I2 => x83_out_22,
   I3 => x83_out_11,
   I4 => x83_out_7,
   O => W_50_7_i_14_n_0
);
W_50_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x59_out_3,
   I1 => x83_out_6,
   I2 => x83_out_10,
   I3 => x83_out_21,
   I4 => x86_out_3,
   O => W_50_7_i_15_n_0
);
W_50_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x86_out_3,
   I1 => x59_out_3,
   I2 => x83_out_21,
   I3 => x83_out_10,
   I4 => x83_out_6,
   O => W_50_7_i_16_n_0
);
W_50_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x59_out_2,
   I1 => x83_out_5,
   I2 => x83_out_9,
   I3 => x83_out_20,
   I4 => x86_out_2,
   O => W_50_7_i_17_n_0
);
W_50_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x44_out_16,
   I1 => x44_out_23,
   I2 => x44_out_25,
   I3 => W_50_7_i_10_n_0,
   I4 => W_50_7_i_11_n_0,
   O => W_50_7_i_2_n_0
);
W_50_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x44_out_15,
   I1 => x44_out_22,
   I2 => x44_out_24,
   I3 => W_50_7_i_12_n_0,
   I4 => W_50_7_i_13_n_0,
   O => W_50_7_i_3_n_0
);
W_50_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x44_out_14,
   I1 => x44_out_21,
   I2 => x44_out_23,
   I3 => W_50_7_i_14_n_0,
   I4 => W_50_7_i_15_n_0,
   O => W_50_7_i_4_n_0
);
W_50_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x44_out_13,
   I1 => x44_out_20,
   I2 => x44_out_22,
   I3 => W_50_7_i_16_n_0,
   I4 => W_50_7_i_17_n_0,
   O => W_50_7_i_5_n_0
);
W_50_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_50_7_i_2_n_0,
   I1 => W_50_11_i_16_n_0,
   I2 => x44_out_17,
   I3 => x44_out_24,
   I4 => x44_out_26,
   I5 => W_50_11_i_17_n_0,
   O => W_50_7_i_6_n_0
);
W_50_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_50_7_i_3_n_0,
   I1 => W_50_7_i_10_n_0,
   I2 => x44_out_16,
   I3 => x44_out_23,
   I4 => x44_out_25,
   I5 => W_50_7_i_11_n_0,
   O => W_50_7_i_7_n_0
);
W_50_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_50_7_i_4_n_0,
   I1 => W_50_7_i_12_n_0,
   I2 => x44_out_15,
   I3 => x44_out_22,
   I4 => x44_out_24,
   I5 => W_50_7_i_13_n_0,
   O => W_50_7_i_8_n_0
);
W_50_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_50_7_i_5_n_0,
   I1 => W_50_7_i_14_n_0,
   I2 => x44_out_14,
   I3 => x44_out_21,
   I4 => x44_out_23,
   I5 => W_50_7_i_15_n_0,
   O => W_50_7_i_9_n_0
);
W_51_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x83_out_10,
   I1 => x56_out_10,
   I2 => x80_out_28,
   I3 => x80_out_17,
   I4 => x80_out_13,
   O => W_51_11_i_10_n_0
);
W_51_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x56_out_9,
   I1 => x80_out_12,
   I2 => x80_out_16,
   I3 => x80_out_27,
   I4 => x83_out_9,
   O => W_51_11_i_11_n_0
);
W_51_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x83_out_9,
   I1 => x56_out_9,
   I2 => x80_out_27,
   I3 => x80_out_16,
   I4 => x80_out_12,
   O => W_51_11_i_12_n_0
);
W_51_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x56_out_8,
   I1 => x80_out_11,
   I2 => x80_out_15,
   I3 => x80_out_26,
   I4 => x83_out_8,
   O => W_51_11_i_13_n_0
);
W_51_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x83_out_8,
   I1 => x56_out_8,
   I2 => x80_out_26,
   I3 => x80_out_15,
   I4 => x80_out_11,
   O => W_51_11_i_14_n_0
);
W_51_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x56_out_7,
   I1 => x80_out_10,
   I2 => x80_out_14,
   I3 => x80_out_25,
   I4 => x83_out_7,
   O => W_51_11_i_15_n_0
);
W_51_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x83_out_7,
   I1 => x56_out_7,
   I2 => x80_out_25,
   I3 => x80_out_14,
   I4 => x80_out_10,
   O => W_51_11_i_16_n_0
);
W_51_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x56_out_6,
   I1 => x80_out_9,
   I2 => x80_out_13,
   I3 => x80_out_24,
   I4 => x83_out_6,
   O => W_51_11_i_17_n_0
);
W_51_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x41_out_20,
   I1 => x41_out_27,
   I2 => x41_out_29,
   I3 => W_51_11_i_10_n_0,
   I4 => W_51_11_i_11_n_0,
   O => W_51_11_i_2_n_0
);
W_51_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x41_out_19,
   I1 => x41_out_26,
   I2 => x41_out_28,
   I3 => W_51_11_i_12_n_0,
   I4 => W_51_11_i_13_n_0,
   O => W_51_11_i_3_n_0
);
W_51_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x41_out_18,
   I1 => x41_out_25,
   I2 => x41_out_27,
   I3 => W_51_11_i_14_n_0,
   I4 => W_51_11_i_15_n_0,
   O => W_51_11_i_4_n_0
);
W_51_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x41_out_17,
   I1 => x41_out_24,
   I2 => x41_out_26,
   I3 => W_51_11_i_16_n_0,
   I4 => W_51_11_i_17_n_0,
   O => W_51_11_i_5_n_0
);
W_51_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_51_11_i_2_n_0,
   I1 => W_51_15_i_16_n_0,
   I2 => x41_out_21,
   I3 => x41_out_28,
   I4 => x41_out_30,
   I5 => W_51_15_i_17_n_0,
   O => W_51_11_i_6_n_0
);
W_51_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_51_11_i_3_n_0,
   I1 => W_51_11_i_10_n_0,
   I2 => x41_out_20,
   I3 => x41_out_27,
   I4 => x41_out_29,
   I5 => W_51_11_i_11_n_0,
   O => W_51_11_i_7_n_0
);
W_51_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_51_11_i_4_n_0,
   I1 => W_51_11_i_12_n_0,
   I2 => x41_out_19,
   I3 => x41_out_26,
   I4 => x41_out_28,
   I5 => W_51_11_i_13_n_0,
   O => W_51_11_i_8_n_0
);
W_51_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_51_11_i_5_n_0,
   I1 => W_51_11_i_14_n_0,
   I2 => x41_out_18,
   I3 => x41_out_25,
   I4 => x41_out_27,
   I5 => W_51_11_i_15_n_0,
   O => W_51_11_i_9_n_0
);
W_51_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x83_out_14,
   I1 => x56_out_14,
   I2 => x80_out_0,
   I3 => x80_out_21,
   I4 => x80_out_17,
   O => W_51_15_i_10_n_0
);
W_51_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x56_out_13,
   I1 => x80_out_16,
   I2 => x80_out_20,
   I3 => x80_out_31,
   I4 => x83_out_13,
   O => W_51_15_i_11_n_0
);
W_51_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x83_out_13,
   I1 => x56_out_13,
   I2 => x80_out_31,
   I3 => x80_out_20,
   I4 => x80_out_16,
   O => W_51_15_i_12_n_0
);
W_51_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x56_out_12,
   I1 => x80_out_15,
   I2 => x80_out_19,
   I3 => x80_out_30,
   I4 => x83_out_12,
   O => W_51_15_i_13_n_0
);
W_51_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x83_out_12,
   I1 => x56_out_12,
   I2 => x80_out_30,
   I3 => x80_out_19,
   I4 => x80_out_15,
   O => W_51_15_i_14_n_0
);
W_51_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x56_out_11,
   I1 => x80_out_14,
   I2 => x80_out_18,
   I3 => x80_out_29,
   I4 => x83_out_11,
   O => W_51_15_i_15_n_0
);
W_51_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x83_out_11,
   I1 => x56_out_11,
   I2 => x80_out_29,
   I3 => x80_out_18,
   I4 => x80_out_14,
   O => W_51_15_i_16_n_0
);
W_51_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x56_out_10,
   I1 => x80_out_13,
   I2 => x80_out_17,
   I3 => x80_out_28,
   I4 => x83_out_10,
   O => W_51_15_i_17_n_0
);
W_51_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x41_out_24,
   I1 => x41_out_31,
   I2 => x41_out_1,
   I3 => W_51_15_i_10_n_0,
   I4 => W_51_15_i_11_n_0,
   O => W_51_15_i_2_n_0
);
W_51_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x41_out_23,
   I1 => x41_out_30,
   I2 => x41_out_0,
   I3 => W_51_15_i_12_n_0,
   I4 => W_51_15_i_13_n_0,
   O => W_51_15_i_3_n_0
);
W_51_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x41_out_22,
   I1 => x41_out_29,
   I2 => x41_out_31,
   I3 => W_51_15_i_14_n_0,
   I4 => W_51_15_i_15_n_0,
   O => W_51_15_i_4_n_0
);
W_51_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x41_out_21,
   I1 => x41_out_28,
   I2 => x41_out_30,
   I3 => W_51_15_i_16_n_0,
   I4 => W_51_15_i_17_n_0,
   O => W_51_15_i_5_n_0
);
W_51_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_51_15_i_2_n_0,
   I1 => W_51_19_i_16_n_0,
   I2 => x41_out_25,
   I3 => x41_out_0,
   I4 => x41_out_2,
   I5 => W_51_19_i_17_n_0,
   O => W_51_15_i_6_n_0
);
W_51_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_51_15_i_3_n_0,
   I1 => W_51_15_i_10_n_0,
   I2 => x41_out_24,
   I3 => x41_out_31,
   I4 => x41_out_1,
   I5 => W_51_15_i_11_n_0,
   O => W_51_15_i_7_n_0
);
W_51_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_51_15_i_4_n_0,
   I1 => W_51_15_i_12_n_0,
   I2 => x41_out_23,
   I3 => x41_out_30,
   I4 => x41_out_0,
   I5 => W_51_15_i_13_n_0,
   O => W_51_15_i_8_n_0
);
W_51_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_51_15_i_5_n_0,
   I1 => W_51_15_i_14_n_0,
   I2 => x41_out_22,
   I3 => x41_out_29,
   I4 => x41_out_31,
   I5 => W_51_15_i_15_n_0,
   O => W_51_15_i_9_n_0
);
W_51_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x83_out_18,
   I1 => x56_out_18,
   I2 => x80_out_4,
   I3 => x80_out_25,
   I4 => x80_out_21,
   O => W_51_19_i_10_n_0
);
W_51_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x56_out_17,
   I1 => x80_out_20,
   I2 => x80_out_24,
   I3 => x80_out_3,
   I4 => x83_out_17,
   O => W_51_19_i_11_n_0
);
W_51_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x83_out_17,
   I1 => x56_out_17,
   I2 => x80_out_3,
   I3 => x80_out_24,
   I4 => x80_out_20,
   O => W_51_19_i_12_n_0
);
W_51_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x56_out_16,
   I1 => x80_out_19,
   I2 => x80_out_23,
   I3 => x80_out_2,
   I4 => x83_out_16,
   O => W_51_19_i_13_n_0
);
W_51_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x83_out_16,
   I1 => x56_out_16,
   I2 => x80_out_2,
   I3 => x80_out_23,
   I4 => x80_out_19,
   O => W_51_19_i_14_n_0
);
W_51_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x56_out_15,
   I1 => x80_out_18,
   I2 => x80_out_22,
   I3 => x80_out_1,
   I4 => x83_out_15,
   O => W_51_19_i_15_n_0
);
W_51_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x83_out_15,
   I1 => x56_out_15,
   I2 => x80_out_1,
   I3 => x80_out_22,
   I4 => x80_out_18,
   O => W_51_19_i_16_n_0
);
W_51_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x56_out_14,
   I1 => x80_out_17,
   I2 => x80_out_21,
   I3 => x80_out_0,
   I4 => x83_out_14,
   O => W_51_19_i_17_n_0
);
W_51_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x41_out_28,
   I1 => x41_out_3,
   I2 => x41_out_5,
   I3 => W_51_19_i_10_n_0,
   I4 => W_51_19_i_11_n_0,
   O => W_51_19_i_2_n_0
);
W_51_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x41_out_27,
   I1 => x41_out_2,
   I2 => x41_out_4,
   I3 => W_51_19_i_12_n_0,
   I4 => W_51_19_i_13_n_0,
   O => W_51_19_i_3_n_0
);
W_51_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x41_out_26,
   I1 => x41_out_1,
   I2 => x41_out_3,
   I3 => W_51_19_i_14_n_0,
   I4 => W_51_19_i_15_n_0,
   O => W_51_19_i_4_n_0
);
W_51_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x41_out_25,
   I1 => x41_out_0,
   I2 => x41_out_2,
   I3 => W_51_19_i_16_n_0,
   I4 => W_51_19_i_17_n_0,
   O => W_51_19_i_5_n_0
);
W_51_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_51_19_i_2_n_0,
   I1 => W_51_23_i_16_n_0,
   I2 => x41_out_29,
   I3 => x41_out_4,
   I4 => x41_out_6,
   I5 => W_51_23_i_17_n_0,
   O => W_51_19_i_6_n_0
);
W_51_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_51_19_i_3_n_0,
   I1 => W_51_19_i_10_n_0,
   I2 => x41_out_28,
   I3 => x41_out_3,
   I4 => x41_out_5,
   I5 => W_51_19_i_11_n_0,
   O => W_51_19_i_7_n_0
);
W_51_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_51_19_i_4_n_0,
   I1 => W_51_19_i_12_n_0,
   I2 => x41_out_27,
   I3 => x41_out_2,
   I4 => x41_out_4,
   I5 => W_51_19_i_13_n_0,
   O => W_51_19_i_8_n_0
);
W_51_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_51_19_i_5_n_0,
   I1 => W_51_19_i_14_n_0,
   I2 => x41_out_26,
   I3 => x41_out_1,
   I4 => x41_out_3,
   I5 => W_51_19_i_15_n_0,
   O => W_51_19_i_9_n_0
);
W_51_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x83_out_22,
   I1 => x56_out_22,
   I2 => x80_out_8,
   I3 => x80_out_29,
   I4 => x80_out_25,
   O => W_51_23_i_10_n_0
);
W_51_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x56_out_21,
   I1 => x80_out_24,
   I2 => x80_out_28,
   I3 => x80_out_7,
   I4 => x83_out_21,
   O => W_51_23_i_11_n_0
);
W_51_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x83_out_21,
   I1 => x56_out_21,
   I2 => x80_out_7,
   I3 => x80_out_28,
   I4 => x80_out_24,
   O => W_51_23_i_12_n_0
);
W_51_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x56_out_20,
   I1 => x80_out_23,
   I2 => x80_out_27,
   I3 => x80_out_6,
   I4 => x83_out_20,
   O => W_51_23_i_13_n_0
);
W_51_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x83_out_20,
   I1 => x56_out_20,
   I2 => x80_out_6,
   I3 => x80_out_27,
   I4 => x80_out_23,
   O => W_51_23_i_14_n_0
);
W_51_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x56_out_19,
   I1 => x80_out_22,
   I2 => x80_out_26,
   I3 => x80_out_5,
   I4 => x83_out_19,
   O => W_51_23_i_15_n_0
);
W_51_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x83_out_19,
   I1 => x56_out_19,
   I2 => x80_out_5,
   I3 => x80_out_26,
   I4 => x80_out_22,
   O => W_51_23_i_16_n_0
);
W_51_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x56_out_18,
   I1 => x80_out_21,
   I2 => x80_out_25,
   I3 => x80_out_4,
   I4 => x83_out_18,
   O => W_51_23_i_17_n_0
);
W_51_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x41_out_7,
   I1 => x41_out_9,
   I2 => W_51_23_i_10_n_0,
   I3 => W_51_23_i_11_n_0,
   O => W_51_23_i_2_n_0
);
W_51_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x41_out_31,
   I1 => x41_out_6,
   I2 => x41_out_8,
   I3 => W_51_23_i_12_n_0,
   I4 => W_51_23_i_13_n_0,
   O => W_51_23_i_3_n_0
);
W_51_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x41_out_30,
   I1 => x41_out_5,
   I2 => x41_out_7,
   I3 => W_51_23_i_14_n_0,
   I4 => W_51_23_i_15_n_0,
   O => W_51_23_i_4_n_0
);
W_51_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x41_out_29,
   I1 => x41_out_4,
   I2 => x41_out_6,
   I3 => W_51_23_i_16_n_0,
   I4 => W_51_23_i_17_n_0,
   O => W_51_23_i_5_n_0
);
W_51_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x41_out_8,
   I1 => x41_out_10,
   I2 => W_51_27_i_16_n_0,
   I3 => W_51_27_i_17_n_0,
   I4 => W_51_23_i_2_n_0,
   O => W_51_23_i_6_n_0
);
W_51_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x41_out_7,
   I1 => x41_out_9,
   I2 => W_51_23_i_10_n_0,
   I3 => W_51_23_i_11_n_0,
   I4 => W_51_23_i_3_n_0,
   O => W_51_23_i_7_n_0
);
W_51_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_51_23_i_4_n_0,
   I1 => W_51_23_i_12_n_0,
   I2 => x41_out_31,
   I3 => x41_out_6,
   I4 => x41_out_8,
   I5 => W_51_23_i_13_n_0,
   O => W_51_23_i_8_n_0
);
W_51_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_51_23_i_5_n_0,
   I1 => W_51_23_i_14_n_0,
   I2 => x41_out_30,
   I3 => x41_out_5,
   I4 => x41_out_7,
   I5 => W_51_23_i_15_n_0,
   O => W_51_23_i_9_n_0
);
W_51_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x83_out_26,
   I1 => x56_out_26,
   I2 => x80_out_12,
   I3 => x80_out_1,
   I4 => x80_out_29,
   O => W_51_27_i_10_n_0
);
W_51_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x56_out_25,
   I1 => x80_out_28,
   I2 => x80_out_0,
   I3 => x80_out_11,
   I4 => x83_out_25,
   O => W_51_27_i_11_n_0
);
W_51_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x83_out_25,
   I1 => x56_out_25,
   I2 => x80_out_11,
   I3 => x80_out_0,
   I4 => x80_out_28,
   O => W_51_27_i_12_n_0
);
W_51_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x56_out_24,
   I1 => x80_out_27,
   I2 => x80_out_31,
   I3 => x80_out_10,
   I4 => x83_out_24,
   O => W_51_27_i_13_n_0
);
W_51_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x83_out_24,
   I1 => x56_out_24,
   I2 => x80_out_10,
   I3 => x80_out_31,
   I4 => x80_out_27,
   O => W_51_27_i_14_n_0
);
W_51_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x56_out_23,
   I1 => x80_out_26,
   I2 => x80_out_30,
   I3 => x80_out_9,
   I4 => x83_out_23,
   O => W_51_27_i_15_n_0
);
W_51_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x83_out_23,
   I1 => x56_out_23,
   I2 => x80_out_9,
   I3 => x80_out_30,
   I4 => x80_out_26,
   O => W_51_27_i_16_n_0
);
W_51_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x56_out_22,
   I1 => x80_out_25,
   I2 => x80_out_29,
   I3 => x80_out_8,
   I4 => x83_out_22,
   O => W_51_27_i_17_n_0
);
W_51_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x41_out_11,
   I1 => x41_out_13,
   I2 => W_51_27_i_10_n_0,
   I3 => W_51_27_i_11_n_0,
   O => W_51_27_i_2_n_0
);
W_51_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x41_out_10,
   I1 => x41_out_12,
   I2 => W_51_27_i_12_n_0,
   I3 => W_51_27_i_13_n_0,
   O => W_51_27_i_3_n_0
);
W_51_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x41_out_9,
   I1 => x41_out_11,
   I2 => W_51_27_i_14_n_0,
   I3 => W_51_27_i_15_n_0,
   O => W_51_27_i_4_n_0
);
W_51_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x41_out_8,
   I1 => x41_out_10,
   I2 => W_51_27_i_16_n_0,
   I3 => W_51_27_i_17_n_0,
   O => W_51_27_i_5_n_0
);
W_51_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x41_out_12,
   I1 => x41_out_14,
   I2 => W_51_31_i_13_n_0,
   I3 => W_51_31_i_14_n_0,
   I4 => W_51_27_i_2_n_0,
   O => W_51_27_i_6_n_0
);
W_51_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x41_out_11,
   I1 => x41_out_13,
   I2 => W_51_27_i_10_n_0,
   I3 => W_51_27_i_11_n_0,
   I4 => W_51_27_i_3_n_0,
   O => W_51_27_i_7_n_0
);
W_51_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x41_out_10,
   I1 => x41_out_12,
   I2 => W_51_27_i_12_n_0,
   I3 => W_51_27_i_13_n_0,
   I4 => W_51_27_i_4_n_0,
   O => W_51_27_i_8_n_0
);
W_51_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x41_out_9,
   I1 => x41_out_11,
   I2 => W_51_27_i_14_n_0,
   I3 => W_51_27_i_15_n_0,
   I4 => W_51_27_i_5_n_0,
   O => W_51_27_i_9_n_0
);
W_51_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x56_out_28,
   I1 => x80_out_31,
   I2 => x80_out_3,
   I3 => x80_out_14,
   I4 => x83_out_28,
   O => W_51_31_i_10_n_0
);
W_51_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x83_out_28,
   I1 => x56_out_28,
   I2 => x80_out_14,
   I3 => x80_out_3,
   I4 => x80_out_31,
   O => W_51_31_i_11_n_0
);
W_51_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x56_out_27,
   I1 => x80_out_30,
   I2 => x80_out_2,
   I3 => x80_out_13,
   I4 => x83_out_27,
   O => W_51_31_i_12_n_0
);
W_51_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x83_out_27,
   I1 => x56_out_27,
   I2 => x80_out_13,
   I3 => x80_out_2,
   I4 => x80_out_30,
   O => W_51_31_i_13_n_0
);
W_51_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x56_out_26,
   I1 => x80_out_29,
   I2 => x80_out_1,
   I3 => x80_out_12,
   I4 => x83_out_26,
   O => W_51_31_i_14_n_0
);
W_51_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x56_out_29,
   I1 => x80_out_4,
   I2 => x80_out_15,
   I3 => x83_out_29,
   O => W_51_31_i_15_n_0
);
W_51_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x41_out_17,
   I1 => x41_out_15,
   O => SIGMA_LCASE_1107_out_0_30
);
W_51_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => x80_out_6,
   I1 => x80_out_17,
   I2 => x56_out_31,
   I3 => x83_out_31,
   I4 => x41_out_16,
   I5 => x41_out_18,
   O => W_51_31_i_17_n_0
);
W_51_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x80_out_16,
   I1 => x80_out_5,
   O => SIGMA_LCASE_0103_out_30
);
W_51_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x83_out_30,
   I1 => x56_out_30,
   I2 => x80_out_16,
   I3 => x80_out_5,
   O => W_51_31_i_19_n_0
);
W_51_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x41_out_14,
   I1 => x41_out_16,
   I2 => W_51_31_i_9_n_0,
   I3 => W_51_31_i_10_n_0,
   O => W_51_31_i_2_n_0
);
W_51_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x41_out_13,
   I1 => x41_out_15,
   I2 => W_51_31_i_11_n_0,
   I3 => W_51_31_i_12_n_0,
   O => W_51_31_i_3_n_0
);
W_51_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x41_out_12,
   I1 => x41_out_14,
   I2 => W_51_31_i_13_n_0,
   I3 => W_51_31_i_14_n_0,
   O => W_51_31_i_4_n_0
);
W_51_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_51_31_i_15_n_0,
   I1 => SIGMA_LCASE_1107_out_0_30,
   I2 => W_51_31_i_17_n_0,
   I3 => x56_out_30,
   I4 => SIGMA_LCASE_0103_out_30,
   I5 => x83_out_30,
   O => W_51_31_i_5_n_0
);
W_51_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_51_31_i_2_n_0,
   I1 => W_51_31_i_19_n_0,
   I2 => x41_out_15,
   I3 => x41_out_17,
   I4 => W_51_31_i_15_n_0,
   O => W_51_31_i_6_n_0
);
W_51_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x41_out_14,
   I1 => x41_out_16,
   I2 => W_51_31_i_9_n_0,
   I3 => W_51_31_i_10_n_0,
   I4 => W_51_31_i_3_n_0,
   O => W_51_31_i_7_n_0
);
W_51_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x41_out_13,
   I1 => x41_out_15,
   I2 => W_51_31_i_11_n_0,
   I3 => W_51_31_i_12_n_0,
   I4 => W_51_31_i_4_n_0,
   O => W_51_31_i_8_n_0
);
W_51_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x83_out_29,
   I1 => x56_out_29,
   I2 => x80_out_15,
   I3 => x80_out_4,
   O => W_51_31_i_9_n_0
);
W_51_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x83_out_2,
   I1 => x56_out_2,
   I2 => x80_out_20,
   I3 => x80_out_9,
   I4 => x80_out_5,
   O => W_51_3_i_10_n_0
);
W_51_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x56_out_1,
   I1 => x80_out_4,
   I2 => x80_out_8,
   I3 => x80_out_19,
   I4 => x83_out_1,
   O => W_51_3_i_11_n_0
);
W_51_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x80_out_19,
   I1 => x80_out_8,
   I2 => x80_out_4,
   O => SIGMA_LCASE_0103_out_1
);
W_51_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x41_out_21,
   I1 => x41_out_19,
   I2 => x41_out_12,
   O => SIGMA_LCASE_1107_out_0_2
);
W_51_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x41_out_20,
   I1 => x41_out_18,
   I2 => x41_out_11,
   O => SIGMA_LCASE_1107_out_1
);
W_51_3_i_15 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x83_out_1,
   I1 => x56_out_1,
   I2 => x80_out_19,
   I3 => x80_out_8,
   I4 => x80_out_4,
   O => W_51_3_i_15_n_0
);
W_51_3_i_16 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x80_out_18,
   I1 => x80_out_7,
   I2 => x80_out_3,
   O => SIGMA_LCASE_0103_out_0
);
W_51_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x41_out_12,
   I1 => x41_out_19,
   I2 => x41_out_21,
   I3 => W_51_3_i_10_n_0,
   I4 => W_51_3_i_11_n_0,
   O => W_51_3_i_2_n_0
);
W_51_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_51_3_i_11_n_0,
   I1 => x41_out_21,
   I2 => x41_out_19,
   I3 => x41_out_12,
   I4 => W_51_3_i_10_n_0,
   O => W_51_3_i_3_n_0
);
W_51_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_0103_out_1,
   I1 => x56_out_1,
   I2 => x83_out_1,
   I3 => x41_out_11,
   I4 => x41_out_18,
   I5 => x41_out_20,
   O => W_51_3_i_4_n_0
);
W_51_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x83_out_0,
   I1 => x56_out_0,
   I2 => x80_out_18,
   I3 => x80_out_7,
   I4 => x80_out_3,
   O => W_51_3_i_5_n_0
);
W_51_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_51_3_i_2_n_0,
   I1 => W_51_7_i_16_n_0,
   I2 => x41_out_13,
   I3 => x41_out_20,
   I4 => x41_out_22,
   I5 => W_51_7_i_17_n_0,
   O => W_51_3_i_6_n_0
);
W_51_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_51_3_i_10_n_0,
   I1 => SIGMA_LCASE_1107_out_0_2,
   I2 => x83_out_1,
   I3 => x56_out_1,
   I4 => SIGMA_LCASE_0103_out_1,
   I5 => SIGMA_LCASE_1107_out_1,
   O => W_51_3_i_7_n_0
);
W_51_3_i_8 : LUT5
  generic map(
   INIT => X"99969666"
  )
 port map (
   I0 => SIGMA_LCASE_1107_out_1,
   I1 => W_51_3_i_15_n_0,
   I2 => x83_out_0,
   I3 => SIGMA_LCASE_0103_out_0,
   I4 => x56_out_0,
   O => W_51_3_i_8_n_0
);
W_51_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_51_3_i_5_n_0,
   I1 => x41_out_10,
   I2 => x41_out_17,
   I3 => x41_out_19,
   O => W_51_3_i_9_n_0
);
W_51_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x83_out_6,
   I1 => x56_out_6,
   I2 => x80_out_24,
   I3 => x80_out_13,
   I4 => x80_out_9,
   O => W_51_7_i_10_n_0
);
W_51_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x56_out_5,
   I1 => x80_out_8,
   I2 => x80_out_12,
   I3 => x80_out_23,
   I4 => x83_out_5,
   O => W_51_7_i_11_n_0
);
W_51_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x83_out_5,
   I1 => x56_out_5,
   I2 => x80_out_23,
   I3 => x80_out_12,
   I4 => x80_out_8,
   O => W_51_7_i_12_n_0
);
W_51_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x56_out_4,
   I1 => x80_out_7,
   I2 => x80_out_11,
   I3 => x80_out_22,
   I4 => x83_out_4,
   O => W_51_7_i_13_n_0
);
W_51_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x83_out_4,
   I1 => x56_out_4,
   I2 => x80_out_22,
   I3 => x80_out_11,
   I4 => x80_out_7,
   O => W_51_7_i_14_n_0
);
W_51_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x56_out_3,
   I1 => x80_out_6,
   I2 => x80_out_10,
   I3 => x80_out_21,
   I4 => x83_out_3,
   O => W_51_7_i_15_n_0
);
W_51_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x83_out_3,
   I1 => x56_out_3,
   I2 => x80_out_21,
   I3 => x80_out_10,
   I4 => x80_out_6,
   O => W_51_7_i_16_n_0
);
W_51_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x56_out_2,
   I1 => x80_out_5,
   I2 => x80_out_9,
   I3 => x80_out_20,
   I4 => x83_out_2,
   O => W_51_7_i_17_n_0
);
W_51_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x41_out_16,
   I1 => x41_out_23,
   I2 => x41_out_25,
   I3 => W_51_7_i_10_n_0,
   I4 => W_51_7_i_11_n_0,
   O => W_51_7_i_2_n_0
);
W_51_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x41_out_15,
   I1 => x41_out_22,
   I2 => x41_out_24,
   I3 => W_51_7_i_12_n_0,
   I4 => W_51_7_i_13_n_0,
   O => W_51_7_i_3_n_0
);
W_51_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x41_out_14,
   I1 => x41_out_21,
   I2 => x41_out_23,
   I3 => W_51_7_i_14_n_0,
   I4 => W_51_7_i_15_n_0,
   O => W_51_7_i_4_n_0
);
W_51_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x41_out_13,
   I1 => x41_out_20,
   I2 => x41_out_22,
   I3 => W_51_7_i_16_n_0,
   I4 => W_51_7_i_17_n_0,
   O => W_51_7_i_5_n_0
);
W_51_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_51_7_i_2_n_0,
   I1 => W_51_11_i_16_n_0,
   I2 => x41_out_17,
   I3 => x41_out_24,
   I4 => x41_out_26,
   I5 => W_51_11_i_17_n_0,
   O => W_51_7_i_6_n_0
);
W_51_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_51_7_i_3_n_0,
   I1 => W_51_7_i_10_n_0,
   I2 => x41_out_16,
   I3 => x41_out_23,
   I4 => x41_out_25,
   I5 => W_51_7_i_11_n_0,
   O => W_51_7_i_7_n_0
);
W_51_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_51_7_i_4_n_0,
   I1 => W_51_7_i_12_n_0,
   I2 => x41_out_15,
   I3 => x41_out_22,
   I4 => x41_out_24,
   I5 => W_51_7_i_13_n_0,
   O => W_51_7_i_8_n_0
);
W_51_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_51_7_i_5_n_0,
   I1 => W_51_7_i_14_n_0,
   I2 => x41_out_14,
   I3 => x41_out_21,
   I4 => x41_out_23,
   I5 => W_51_7_i_15_n_0,
   O => W_51_7_i_9_n_0
);
W_52_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x80_out_10,
   I1 => x53_out_10,
   I2 => x77_out_28,
   I3 => x77_out_17,
   I4 => x77_out_13,
   O => W_52_11_i_10_n_0
);
W_52_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x53_out_9,
   I1 => x77_out_12,
   I2 => x77_out_16,
   I3 => x77_out_27,
   I4 => x80_out_9,
   O => W_52_11_i_11_n_0
);
W_52_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x80_out_9,
   I1 => x53_out_9,
   I2 => x77_out_27,
   I3 => x77_out_16,
   I4 => x77_out_12,
   O => W_52_11_i_12_n_0
);
W_52_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x53_out_8,
   I1 => x77_out_11,
   I2 => x77_out_15,
   I3 => x77_out_26,
   I4 => x80_out_8,
   O => W_52_11_i_13_n_0
);
W_52_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x80_out_8,
   I1 => x53_out_8,
   I2 => x77_out_26,
   I3 => x77_out_15,
   I4 => x77_out_11,
   O => W_52_11_i_14_n_0
);
W_52_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x53_out_7,
   I1 => x77_out_10,
   I2 => x77_out_14,
   I3 => x77_out_25,
   I4 => x80_out_7,
   O => W_52_11_i_15_n_0
);
W_52_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x80_out_7,
   I1 => x53_out_7,
   I2 => x77_out_25,
   I3 => x77_out_14,
   I4 => x77_out_10,
   O => W_52_11_i_16_n_0
);
W_52_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x53_out_6,
   I1 => x77_out_9,
   I2 => x77_out_13,
   I3 => x77_out_24,
   I4 => x80_out_6,
   O => W_52_11_i_17_n_0
);
W_52_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x38_out_20,
   I1 => x38_out_27,
   I2 => x38_out_29,
   I3 => W_52_11_i_10_n_0,
   I4 => W_52_11_i_11_n_0,
   O => W_52_11_i_2_n_0
);
W_52_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x38_out_19,
   I1 => x38_out_26,
   I2 => x38_out_28,
   I3 => W_52_11_i_12_n_0,
   I4 => W_52_11_i_13_n_0,
   O => W_52_11_i_3_n_0
);
W_52_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x38_out_18,
   I1 => x38_out_25,
   I2 => x38_out_27,
   I3 => W_52_11_i_14_n_0,
   I4 => W_52_11_i_15_n_0,
   O => W_52_11_i_4_n_0
);
W_52_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x38_out_17,
   I1 => x38_out_24,
   I2 => x38_out_26,
   I3 => W_52_11_i_16_n_0,
   I4 => W_52_11_i_17_n_0,
   O => W_52_11_i_5_n_0
);
W_52_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_52_11_i_2_n_0,
   I1 => W_52_15_i_16_n_0,
   I2 => x38_out_21,
   I3 => x38_out_28,
   I4 => x38_out_30,
   I5 => W_52_15_i_17_n_0,
   O => W_52_11_i_6_n_0
);
W_52_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_52_11_i_3_n_0,
   I1 => W_52_11_i_10_n_0,
   I2 => x38_out_20,
   I3 => x38_out_27,
   I4 => x38_out_29,
   I5 => W_52_11_i_11_n_0,
   O => W_52_11_i_7_n_0
);
W_52_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_52_11_i_4_n_0,
   I1 => W_52_11_i_12_n_0,
   I2 => x38_out_19,
   I3 => x38_out_26,
   I4 => x38_out_28,
   I5 => W_52_11_i_13_n_0,
   O => W_52_11_i_8_n_0
);
W_52_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_52_11_i_5_n_0,
   I1 => W_52_11_i_14_n_0,
   I2 => x38_out_18,
   I3 => x38_out_25,
   I4 => x38_out_27,
   I5 => W_52_11_i_15_n_0,
   O => W_52_11_i_9_n_0
);
W_52_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x80_out_14,
   I1 => x53_out_14,
   I2 => x77_out_0,
   I3 => x77_out_21,
   I4 => x77_out_17,
   O => W_52_15_i_10_n_0
);
W_52_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x53_out_13,
   I1 => x77_out_16,
   I2 => x77_out_20,
   I3 => x77_out_31,
   I4 => x80_out_13,
   O => W_52_15_i_11_n_0
);
W_52_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x80_out_13,
   I1 => x53_out_13,
   I2 => x77_out_31,
   I3 => x77_out_20,
   I4 => x77_out_16,
   O => W_52_15_i_12_n_0
);
W_52_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x53_out_12,
   I1 => x77_out_15,
   I2 => x77_out_19,
   I3 => x77_out_30,
   I4 => x80_out_12,
   O => W_52_15_i_13_n_0
);
W_52_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x80_out_12,
   I1 => x53_out_12,
   I2 => x77_out_30,
   I3 => x77_out_19,
   I4 => x77_out_15,
   O => W_52_15_i_14_n_0
);
W_52_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x53_out_11,
   I1 => x77_out_14,
   I2 => x77_out_18,
   I3 => x77_out_29,
   I4 => x80_out_11,
   O => W_52_15_i_15_n_0
);
W_52_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x80_out_11,
   I1 => x53_out_11,
   I2 => x77_out_29,
   I3 => x77_out_18,
   I4 => x77_out_14,
   O => W_52_15_i_16_n_0
);
W_52_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x53_out_10,
   I1 => x77_out_13,
   I2 => x77_out_17,
   I3 => x77_out_28,
   I4 => x80_out_10,
   O => W_52_15_i_17_n_0
);
W_52_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x38_out_24,
   I1 => x38_out_31,
   I2 => x38_out_1,
   I3 => W_52_15_i_10_n_0,
   I4 => W_52_15_i_11_n_0,
   O => W_52_15_i_2_n_0
);
W_52_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x38_out_23,
   I1 => x38_out_30,
   I2 => x38_out_0,
   I3 => W_52_15_i_12_n_0,
   I4 => W_52_15_i_13_n_0,
   O => W_52_15_i_3_n_0
);
W_52_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x38_out_22,
   I1 => x38_out_29,
   I2 => x38_out_31,
   I3 => W_52_15_i_14_n_0,
   I4 => W_52_15_i_15_n_0,
   O => W_52_15_i_4_n_0
);
W_52_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x38_out_21,
   I1 => x38_out_28,
   I2 => x38_out_30,
   I3 => W_52_15_i_16_n_0,
   I4 => W_52_15_i_17_n_0,
   O => W_52_15_i_5_n_0
);
W_52_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_52_15_i_2_n_0,
   I1 => W_52_19_i_16_n_0,
   I2 => x38_out_25,
   I3 => x38_out_0,
   I4 => x38_out_2,
   I5 => W_52_19_i_17_n_0,
   O => W_52_15_i_6_n_0
);
W_52_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_52_15_i_3_n_0,
   I1 => W_52_15_i_10_n_0,
   I2 => x38_out_24,
   I3 => x38_out_31,
   I4 => x38_out_1,
   I5 => W_52_15_i_11_n_0,
   O => W_52_15_i_7_n_0
);
W_52_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_52_15_i_4_n_0,
   I1 => W_52_15_i_12_n_0,
   I2 => x38_out_23,
   I3 => x38_out_30,
   I4 => x38_out_0,
   I5 => W_52_15_i_13_n_0,
   O => W_52_15_i_8_n_0
);
W_52_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_52_15_i_5_n_0,
   I1 => W_52_15_i_14_n_0,
   I2 => x38_out_22,
   I3 => x38_out_29,
   I4 => x38_out_31,
   I5 => W_52_15_i_15_n_0,
   O => W_52_15_i_9_n_0
);
W_52_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x80_out_18,
   I1 => x53_out_18,
   I2 => x77_out_4,
   I3 => x77_out_25,
   I4 => x77_out_21,
   O => W_52_19_i_10_n_0
);
W_52_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x53_out_17,
   I1 => x77_out_20,
   I2 => x77_out_24,
   I3 => x77_out_3,
   I4 => x80_out_17,
   O => W_52_19_i_11_n_0
);
W_52_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x80_out_17,
   I1 => x53_out_17,
   I2 => x77_out_3,
   I3 => x77_out_24,
   I4 => x77_out_20,
   O => W_52_19_i_12_n_0
);
W_52_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x53_out_16,
   I1 => x77_out_19,
   I2 => x77_out_23,
   I3 => x77_out_2,
   I4 => x80_out_16,
   O => W_52_19_i_13_n_0
);
W_52_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x80_out_16,
   I1 => x53_out_16,
   I2 => x77_out_2,
   I3 => x77_out_23,
   I4 => x77_out_19,
   O => W_52_19_i_14_n_0
);
W_52_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x53_out_15,
   I1 => x77_out_18,
   I2 => x77_out_22,
   I3 => x77_out_1,
   I4 => x80_out_15,
   O => W_52_19_i_15_n_0
);
W_52_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x80_out_15,
   I1 => x53_out_15,
   I2 => x77_out_1,
   I3 => x77_out_22,
   I4 => x77_out_18,
   O => W_52_19_i_16_n_0
);
W_52_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x53_out_14,
   I1 => x77_out_17,
   I2 => x77_out_21,
   I3 => x77_out_0,
   I4 => x80_out_14,
   O => W_52_19_i_17_n_0
);
W_52_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x38_out_28,
   I1 => x38_out_3,
   I2 => x38_out_5,
   I3 => W_52_19_i_10_n_0,
   I4 => W_52_19_i_11_n_0,
   O => W_52_19_i_2_n_0
);
W_52_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x38_out_27,
   I1 => x38_out_2,
   I2 => x38_out_4,
   I3 => W_52_19_i_12_n_0,
   I4 => W_52_19_i_13_n_0,
   O => W_52_19_i_3_n_0
);
W_52_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x38_out_26,
   I1 => x38_out_1,
   I2 => x38_out_3,
   I3 => W_52_19_i_14_n_0,
   I4 => W_52_19_i_15_n_0,
   O => W_52_19_i_4_n_0
);
W_52_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x38_out_25,
   I1 => x38_out_0,
   I2 => x38_out_2,
   I3 => W_52_19_i_16_n_0,
   I4 => W_52_19_i_17_n_0,
   O => W_52_19_i_5_n_0
);
W_52_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_52_19_i_2_n_0,
   I1 => W_52_23_i_16_n_0,
   I2 => x38_out_29,
   I3 => x38_out_4,
   I4 => x38_out_6,
   I5 => W_52_23_i_17_n_0,
   O => W_52_19_i_6_n_0
);
W_52_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_52_19_i_3_n_0,
   I1 => W_52_19_i_10_n_0,
   I2 => x38_out_28,
   I3 => x38_out_3,
   I4 => x38_out_5,
   I5 => W_52_19_i_11_n_0,
   O => W_52_19_i_7_n_0
);
W_52_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_52_19_i_4_n_0,
   I1 => W_52_19_i_12_n_0,
   I2 => x38_out_27,
   I3 => x38_out_2,
   I4 => x38_out_4,
   I5 => W_52_19_i_13_n_0,
   O => W_52_19_i_8_n_0
);
W_52_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_52_19_i_5_n_0,
   I1 => W_52_19_i_14_n_0,
   I2 => x38_out_26,
   I3 => x38_out_1,
   I4 => x38_out_3,
   I5 => W_52_19_i_15_n_0,
   O => W_52_19_i_9_n_0
);
W_52_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x80_out_22,
   I1 => x53_out_22,
   I2 => x77_out_8,
   I3 => x77_out_29,
   I4 => x77_out_25,
   O => W_52_23_i_10_n_0
);
W_52_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x53_out_21,
   I1 => x77_out_24,
   I2 => x77_out_28,
   I3 => x77_out_7,
   I4 => x80_out_21,
   O => W_52_23_i_11_n_0
);
W_52_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x80_out_21,
   I1 => x53_out_21,
   I2 => x77_out_7,
   I3 => x77_out_28,
   I4 => x77_out_24,
   O => W_52_23_i_12_n_0
);
W_52_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x53_out_20,
   I1 => x77_out_23,
   I2 => x77_out_27,
   I3 => x77_out_6,
   I4 => x80_out_20,
   O => W_52_23_i_13_n_0
);
W_52_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x80_out_20,
   I1 => x53_out_20,
   I2 => x77_out_6,
   I3 => x77_out_27,
   I4 => x77_out_23,
   O => W_52_23_i_14_n_0
);
W_52_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x53_out_19,
   I1 => x77_out_22,
   I2 => x77_out_26,
   I3 => x77_out_5,
   I4 => x80_out_19,
   O => W_52_23_i_15_n_0
);
W_52_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x80_out_19,
   I1 => x53_out_19,
   I2 => x77_out_5,
   I3 => x77_out_26,
   I4 => x77_out_22,
   O => W_52_23_i_16_n_0
);
W_52_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x53_out_18,
   I1 => x77_out_21,
   I2 => x77_out_25,
   I3 => x77_out_4,
   I4 => x80_out_18,
   O => W_52_23_i_17_n_0
);
W_52_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x38_out_7,
   I1 => x38_out_9,
   I2 => W_52_23_i_10_n_0,
   I3 => W_52_23_i_11_n_0,
   O => W_52_23_i_2_n_0
);
W_52_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x38_out_31,
   I1 => x38_out_6,
   I2 => x38_out_8,
   I3 => W_52_23_i_12_n_0,
   I4 => W_52_23_i_13_n_0,
   O => W_52_23_i_3_n_0
);
W_52_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x38_out_30,
   I1 => x38_out_5,
   I2 => x38_out_7,
   I3 => W_52_23_i_14_n_0,
   I4 => W_52_23_i_15_n_0,
   O => W_52_23_i_4_n_0
);
W_52_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x38_out_29,
   I1 => x38_out_4,
   I2 => x38_out_6,
   I3 => W_52_23_i_16_n_0,
   I4 => W_52_23_i_17_n_0,
   O => W_52_23_i_5_n_0
);
W_52_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x38_out_8,
   I1 => x38_out_10,
   I2 => W_52_27_i_16_n_0,
   I3 => W_52_27_i_17_n_0,
   I4 => W_52_23_i_2_n_0,
   O => W_52_23_i_6_n_0
);
W_52_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x38_out_7,
   I1 => x38_out_9,
   I2 => W_52_23_i_10_n_0,
   I3 => W_52_23_i_11_n_0,
   I4 => W_52_23_i_3_n_0,
   O => W_52_23_i_7_n_0
);
W_52_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_52_23_i_4_n_0,
   I1 => W_52_23_i_12_n_0,
   I2 => x38_out_31,
   I3 => x38_out_6,
   I4 => x38_out_8,
   I5 => W_52_23_i_13_n_0,
   O => W_52_23_i_8_n_0
);
W_52_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_52_23_i_5_n_0,
   I1 => W_52_23_i_14_n_0,
   I2 => x38_out_30,
   I3 => x38_out_5,
   I4 => x38_out_7,
   I5 => W_52_23_i_15_n_0,
   O => W_52_23_i_9_n_0
);
W_52_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x80_out_26,
   I1 => x53_out_26,
   I2 => x77_out_12,
   I3 => x77_out_1,
   I4 => x77_out_29,
   O => W_52_27_i_10_n_0
);
W_52_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x53_out_25,
   I1 => x77_out_28,
   I2 => x77_out_0,
   I3 => x77_out_11,
   I4 => x80_out_25,
   O => W_52_27_i_11_n_0
);
W_52_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x80_out_25,
   I1 => x53_out_25,
   I2 => x77_out_11,
   I3 => x77_out_0,
   I4 => x77_out_28,
   O => W_52_27_i_12_n_0
);
W_52_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x53_out_24,
   I1 => x77_out_27,
   I2 => x77_out_31,
   I3 => x77_out_10,
   I4 => x80_out_24,
   O => W_52_27_i_13_n_0
);
W_52_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x80_out_24,
   I1 => x53_out_24,
   I2 => x77_out_10,
   I3 => x77_out_31,
   I4 => x77_out_27,
   O => W_52_27_i_14_n_0
);
W_52_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x53_out_23,
   I1 => x77_out_26,
   I2 => x77_out_30,
   I3 => x77_out_9,
   I4 => x80_out_23,
   O => W_52_27_i_15_n_0
);
W_52_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x80_out_23,
   I1 => x53_out_23,
   I2 => x77_out_9,
   I3 => x77_out_30,
   I4 => x77_out_26,
   O => W_52_27_i_16_n_0
);
W_52_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x53_out_22,
   I1 => x77_out_25,
   I2 => x77_out_29,
   I3 => x77_out_8,
   I4 => x80_out_22,
   O => W_52_27_i_17_n_0
);
W_52_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x38_out_11,
   I1 => x38_out_13,
   I2 => W_52_27_i_10_n_0,
   I3 => W_52_27_i_11_n_0,
   O => W_52_27_i_2_n_0
);
W_52_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x38_out_10,
   I1 => x38_out_12,
   I2 => W_52_27_i_12_n_0,
   I3 => W_52_27_i_13_n_0,
   O => W_52_27_i_3_n_0
);
W_52_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x38_out_9,
   I1 => x38_out_11,
   I2 => W_52_27_i_14_n_0,
   I3 => W_52_27_i_15_n_0,
   O => W_52_27_i_4_n_0
);
W_52_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x38_out_8,
   I1 => x38_out_10,
   I2 => W_52_27_i_16_n_0,
   I3 => W_52_27_i_17_n_0,
   O => W_52_27_i_5_n_0
);
W_52_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x38_out_12,
   I1 => x38_out_14,
   I2 => W_52_31_i_13_n_0,
   I3 => W_52_31_i_14_n_0,
   I4 => W_52_27_i_2_n_0,
   O => W_52_27_i_6_n_0
);
W_52_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x38_out_11,
   I1 => x38_out_13,
   I2 => W_52_27_i_10_n_0,
   I3 => W_52_27_i_11_n_0,
   I4 => W_52_27_i_3_n_0,
   O => W_52_27_i_7_n_0
);
W_52_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x38_out_10,
   I1 => x38_out_12,
   I2 => W_52_27_i_12_n_0,
   I3 => W_52_27_i_13_n_0,
   I4 => W_52_27_i_4_n_0,
   O => W_52_27_i_8_n_0
);
W_52_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x38_out_9,
   I1 => x38_out_11,
   I2 => W_52_27_i_14_n_0,
   I3 => W_52_27_i_15_n_0,
   I4 => W_52_27_i_5_n_0,
   O => W_52_27_i_9_n_0
);
W_52_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x53_out_28,
   I1 => x77_out_31,
   I2 => x77_out_3,
   I3 => x77_out_14,
   I4 => x80_out_28,
   O => W_52_31_i_10_n_0
);
W_52_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x80_out_28,
   I1 => x53_out_28,
   I2 => x77_out_14,
   I3 => x77_out_3,
   I4 => x77_out_31,
   O => W_52_31_i_11_n_0
);
W_52_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x53_out_27,
   I1 => x77_out_30,
   I2 => x77_out_2,
   I3 => x77_out_13,
   I4 => x80_out_27,
   O => W_52_31_i_12_n_0
);
W_52_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x80_out_27,
   I1 => x53_out_27,
   I2 => x77_out_13,
   I3 => x77_out_2,
   I4 => x77_out_30,
   O => W_52_31_i_13_n_0
);
W_52_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x53_out_26,
   I1 => x77_out_29,
   I2 => x77_out_1,
   I3 => x77_out_12,
   I4 => x80_out_26,
   O => W_52_31_i_14_n_0
);
W_52_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x53_out_29,
   I1 => x77_out_4,
   I2 => x77_out_15,
   I3 => x80_out_29,
   O => W_52_31_i_15_n_0
);
W_52_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x38_out_17,
   I1 => x38_out_15,
   O => SIGMA_LCASE_199_out_0_30
);
W_52_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => x77_out_6,
   I1 => x77_out_17,
   I2 => x53_out_31,
   I3 => x80_out_31,
   I4 => x38_out_16,
   I5 => x38_out_18,
   O => W_52_31_i_17_n_0
);
W_52_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x77_out_16,
   I1 => x77_out_5,
   O => SIGMA_LCASE_095_out_30
);
W_52_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x80_out_30,
   I1 => x53_out_30,
   I2 => x77_out_16,
   I3 => x77_out_5,
   O => W_52_31_i_19_n_0
);
W_52_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x38_out_14,
   I1 => x38_out_16,
   I2 => W_52_31_i_9_n_0,
   I3 => W_52_31_i_10_n_0,
   O => W_52_31_i_2_n_0
);
W_52_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x38_out_13,
   I1 => x38_out_15,
   I2 => W_52_31_i_11_n_0,
   I3 => W_52_31_i_12_n_0,
   O => W_52_31_i_3_n_0
);
W_52_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x38_out_12,
   I1 => x38_out_14,
   I2 => W_52_31_i_13_n_0,
   I3 => W_52_31_i_14_n_0,
   O => W_52_31_i_4_n_0
);
W_52_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_52_31_i_15_n_0,
   I1 => SIGMA_LCASE_199_out_0_30,
   I2 => W_52_31_i_17_n_0,
   I3 => x53_out_30,
   I4 => SIGMA_LCASE_095_out_30,
   I5 => x80_out_30,
   O => W_52_31_i_5_n_0
);
W_52_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_52_31_i_2_n_0,
   I1 => W_52_31_i_19_n_0,
   I2 => x38_out_15,
   I3 => x38_out_17,
   I4 => W_52_31_i_15_n_0,
   O => W_52_31_i_6_n_0
);
W_52_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x38_out_14,
   I1 => x38_out_16,
   I2 => W_52_31_i_9_n_0,
   I3 => W_52_31_i_10_n_0,
   I4 => W_52_31_i_3_n_0,
   O => W_52_31_i_7_n_0
);
W_52_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x38_out_13,
   I1 => x38_out_15,
   I2 => W_52_31_i_11_n_0,
   I3 => W_52_31_i_12_n_0,
   I4 => W_52_31_i_4_n_0,
   O => W_52_31_i_8_n_0
);
W_52_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x80_out_29,
   I1 => x53_out_29,
   I2 => x77_out_15,
   I3 => x77_out_4,
   O => W_52_31_i_9_n_0
);
W_52_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x80_out_2,
   I1 => x53_out_2,
   I2 => x77_out_20,
   I3 => x77_out_9,
   I4 => x77_out_5,
   O => W_52_3_i_10_n_0
);
W_52_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x53_out_1,
   I1 => x77_out_4,
   I2 => x77_out_8,
   I3 => x77_out_19,
   I4 => x80_out_1,
   O => W_52_3_i_11_n_0
);
W_52_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x77_out_19,
   I1 => x77_out_8,
   I2 => x77_out_4,
   O => SIGMA_LCASE_095_out_1
);
W_52_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x38_out_21,
   I1 => x38_out_19,
   I2 => x38_out_12,
   O => SIGMA_LCASE_199_out_0_2
);
W_52_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x38_out_20,
   I1 => x38_out_18,
   I2 => x38_out_11,
   O => SIGMA_LCASE_199_out_1
);
W_52_3_i_15 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x80_out_1,
   I1 => x53_out_1,
   I2 => x77_out_19,
   I3 => x77_out_8,
   I4 => x77_out_4,
   O => W_52_3_i_15_n_0
);
W_52_3_i_16 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x77_out_18,
   I1 => x77_out_7,
   I2 => x77_out_3,
   O => SIGMA_LCASE_095_out_0
);
W_52_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x38_out_12,
   I1 => x38_out_19,
   I2 => x38_out_21,
   I3 => W_52_3_i_10_n_0,
   I4 => W_52_3_i_11_n_0,
   O => W_52_3_i_2_n_0
);
W_52_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_52_3_i_11_n_0,
   I1 => x38_out_21,
   I2 => x38_out_19,
   I3 => x38_out_12,
   I4 => W_52_3_i_10_n_0,
   O => W_52_3_i_3_n_0
);
W_52_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_095_out_1,
   I1 => x53_out_1,
   I2 => x80_out_1,
   I3 => x38_out_11,
   I4 => x38_out_18,
   I5 => x38_out_20,
   O => W_52_3_i_4_n_0
);
W_52_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x80_out_0,
   I1 => x53_out_0,
   I2 => x77_out_18,
   I3 => x77_out_7,
   I4 => x77_out_3,
   O => W_52_3_i_5_n_0
);
W_52_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_52_3_i_2_n_0,
   I1 => W_52_7_i_16_n_0,
   I2 => x38_out_13,
   I3 => x38_out_20,
   I4 => x38_out_22,
   I5 => W_52_7_i_17_n_0,
   O => W_52_3_i_6_n_0
);
W_52_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_52_3_i_10_n_0,
   I1 => SIGMA_LCASE_199_out_0_2,
   I2 => x80_out_1,
   I3 => x53_out_1,
   I4 => SIGMA_LCASE_095_out_1,
   I5 => SIGMA_LCASE_199_out_1,
   O => W_52_3_i_7_n_0
);
W_52_3_i_8 : LUT5
  generic map(
   INIT => X"99969666"
  )
 port map (
   I0 => SIGMA_LCASE_199_out_1,
   I1 => W_52_3_i_15_n_0,
   I2 => x80_out_0,
   I3 => SIGMA_LCASE_095_out_0,
   I4 => x53_out_0,
   O => W_52_3_i_8_n_0
);
W_52_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_52_3_i_5_n_0,
   I1 => x38_out_10,
   I2 => x38_out_17,
   I3 => x38_out_19,
   O => W_52_3_i_9_n_0
);
W_52_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x80_out_6,
   I1 => x53_out_6,
   I2 => x77_out_24,
   I3 => x77_out_13,
   I4 => x77_out_9,
   O => W_52_7_i_10_n_0
);
W_52_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x53_out_5,
   I1 => x77_out_8,
   I2 => x77_out_12,
   I3 => x77_out_23,
   I4 => x80_out_5,
   O => W_52_7_i_11_n_0
);
W_52_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x80_out_5,
   I1 => x53_out_5,
   I2 => x77_out_23,
   I3 => x77_out_12,
   I4 => x77_out_8,
   O => W_52_7_i_12_n_0
);
W_52_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x53_out_4,
   I1 => x77_out_7,
   I2 => x77_out_11,
   I3 => x77_out_22,
   I4 => x80_out_4,
   O => W_52_7_i_13_n_0
);
W_52_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x80_out_4,
   I1 => x53_out_4,
   I2 => x77_out_22,
   I3 => x77_out_11,
   I4 => x77_out_7,
   O => W_52_7_i_14_n_0
);
W_52_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x53_out_3,
   I1 => x77_out_6,
   I2 => x77_out_10,
   I3 => x77_out_21,
   I4 => x80_out_3,
   O => W_52_7_i_15_n_0
);
W_52_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x80_out_3,
   I1 => x53_out_3,
   I2 => x77_out_21,
   I3 => x77_out_10,
   I4 => x77_out_6,
   O => W_52_7_i_16_n_0
);
W_52_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x53_out_2,
   I1 => x77_out_5,
   I2 => x77_out_9,
   I3 => x77_out_20,
   I4 => x80_out_2,
   O => W_52_7_i_17_n_0
);
W_52_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x38_out_16,
   I1 => x38_out_23,
   I2 => x38_out_25,
   I3 => W_52_7_i_10_n_0,
   I4 => W_52_7_i_11_n_0,
   O => W_52_7_i_2_n_0
);
W_52_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x38_out_15,
   I1 => x38_out_22,
   I2 => x38_out_24,
   I3 => W_52_7_i_12_n_0,
   I4 => W_52_7_i_13_n_0,
   O => W_52_7_i_3_n_0
);
W_52_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x38_out_14,
   I1 => x38_out_21,
   I2 => x38_out_23,
   I3 => W_52_7_i_14_n_0,
   I4 => W_52_7_i_15_n_0,
   O => W_52_7_i_4_n_0
);
W_52_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x38_out_13,
   I1 => x38_out_20,
   I2 => x38_out_22,
   I3 => W_52_7_i_16_n_0,
   I4 => W_52_7_i_17_n_0,
   O => W_52_7_i_5_n_0
);
W_52_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_52_7_i_2_n_0,
   I1 => W_52_11_i_16_n_0,
   I2 => x38_out_17,
   I3 => x38_out_24,
   I4 => x38_out_26,
   I5 => W_52_11_i_17_n_0,
   O => W_52_7_i_6_n_0
);
W_52_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_52_7_i_3_n_0,
   I1 => W_52_7_i_10_n_0,
   I2 => x38_out_16,
   I3 => x38_out_23,
   I4 => x38_out_25,
   I5 => W_52_7_i_11_n_0,
   O => W_52_7_i_7_n_0
);
W_52_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_52_7_i_4_n_0,
   I1 => W_52_7_i_12_n_0,
   I2 => x38_out_15,
   I3 => x38_out_22,
   I4 => x38_out_24,
   I5 => W_52_7_i_13_n_0,
   O => W_52_7_i_8_n_0
);
W_52_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_52_7_i_5_n_0,
   I1 => W_52_7_i_14_n_0,
   I2 => x38_out_14,
   I3 => x38_out_21,
   I4 => x38_out_23,
   I5 => W_52_7_i_15_n_0,
   O => W_52_7_i_9_n_0
);
W_53_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x77_out_10,
   I1 => x50_out_10,
   I2 => x74_out_28,
   I3 => x74_out_17,
   I4 => x74_out_13,
   O => W_53_11_i_10_n_0
);
W_53_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x50_out_9,
   I1 => x74_out_12,
   I2 => x74_out_16,
   I3 => x74_out_27,
   I4 => x77_out_9,
   O => W_53_11_i_11_n_0
);
W_53_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x77_out_9,
   I1 => x50_out_9,
   I2 => x74_out_27,
   I3 => x74_out_16,
   I4 => x74_out_12,
   O => W_53_11_i_12_n_0
);
W_53_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x50_out_8,
   I1 => x74_out_11,
   I2 => x74_out_15,
   I3 => x74_out_26,
   I4 => x77_out_8,
   O => W_53_11_i_13_n_0
);
W_53_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x77_out_8,
   I1 => x50_out_8,
   I2 => x74_out_26,
   I3 => x74_out_15,
   I4 => x74_out_11,
   O => W_53_11_i_14_n_0
);
W_53_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x50_out_7,
   I1 => x74_out_10,
   I2 => x74_out_14,
   I3 => x74_out_25,
   I4 => x77_out_7,
   O => W_53_11_i_15_n_0
);
W_53_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x77_out_7,
   I1 => x50_out_7,
   I2 => x74_out_25,
   I3 => x74_out_14,
   I4 => x74_out_10,
   O => W_53_11_i_16_n_0
);
W_53_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x50_out_6,
   I1 => x74_out_9,
   I2 => x74_out_13,
   I3 => x74_out_24,
   I4 => x77_out_6,
   O => W_53_11_i_17_n_0
);
W_53_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x35_out_20,
   I1 => x35_out_27,
   I2 => x35_out_29,
   I3 => W_53_11_i_10_n_0,
   I4 => W_53_11_i_11_n_0,
   O => W_53_11_i_2_n_0
);
W_53_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x35_out_19,
   I1 => x35_out_26,
   I2 => x35_out_28,
   I3 => W_53_11_i_12_n_0,
   I4 => W_53_11_i_13_n_0,
   O => W_53_11_i_3_n_0
);
W_53_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x35_out_18,
   I1 => x35_out_25,
   I2 => x35_out_27,
   I3 => W_53_11_i_14_n_0,
   I4 => W_53_11_i_15_n_0,
   O => W_53_11_i_4_n_0
);
W_53_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x35_out_17,
   I1 => x35_out_24,
   I2 => x35_out_26,
   I3 => W_53_11_i_16_n_0,
   I4 => W_53_11_i_17_n_0,
   O => W_53_11_i_5_n_0
);
W_53_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_53_11_i_2_n_0,
   I1 => W_53_15_i_16_n_0,
   I2 => x35_out_21,
   I3 => x35_out_28,
   I4 => x35_out_30,
   I5 => W_53_15_i_17_n_0,
   O => W_53_11_i_6_n_0
);
W_53_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_53_11_i_3_n_0,
   I1 => W_53_11_i_10_n_0,
   I2 => x35_out_20,
   I3 => x35_out_27,
   I4 => x35_out_29,
   I5 => W_53_11_i_11_n_0,
   O => W_53_11_i_7_n_0
);
W_53_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_53_11_i_4_n_0,
   I1 => W_53_11_i_12_n_0,
   I2 => x35_out_19,
   I3 => x35_out_26,
   I4 => x35_out_28,
   I5 => W_53_11_i_13_n_0,
   O => W_53_11_i_8_n_0
);
W_53_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_53_11_i_5_n_0,
   I1 => W_53_11_i_14_n_0,
   I2 => x35_out_18,
   I3 => x35_out_25,
   I4 => x35_out_27,
   I5 => W_53_11_i_15_n_0,
   O => W_53_11_i_9_n_0
);
W_53_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x77_out_14,
   I1 => x50_out_14,
   I2 => x74_out_0,
   I3 => x74_out_21,
   I4 => x74_out_17,
   O => W_53_15_i_10_n_0
);
W_53_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x50_out_13,
   I1 => x74_out_16,
   I2 => x74_out_20,
   I3 => x74_out_31,
   I4 => x77_out_13,
   O => W_53_15_i_11_n_0
);
W_53_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x77_out_13,
   I1 => x50_out_13,
   I2 => x74_out_31,
   I3 => x74_out_20,
   I4 => x74_out_16,
   O => W_53_15_i_12_n_0
);
W_53_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x50_out_12,
   I1 => x74_out_15,
   I2 => x74_out_19,
   I3 => x74_out_30,
   I4 => x77_out_12,
   O => W_53_15_i_13_n_0
);
W_53_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x77_out_12,
   I1 => x50_out_12,
   I2 => x74_out_30,
   I3 => x74_out_19,
   I4 => x74_out_15,
   O => W_53_15_i_14_n_0
);
W_53_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x50_out_11,
   I1 => x74_out_14,
   I2 => x74_out_18,
   I3 => x74_out_29,
   I4 => x77_out_11,
   O => W_53_15_i_15_n_0
);
W_53_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x77_out_11,
   I1 => x50_out_11,
   I2 => x74_out_29,
   I3 => x74_out_18,
   I4 => x74_out_14,
   O => W_53_15_i_16_n_0
);
W_53_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x50_out_10,
   I1 => x74_out_13,
   I2 => x74_out_17,
   I3 => x74_out_28,
   I4 => x77_out_10,
   O => W_53_15_i_17_n_0
);
W_53_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x35_out_24,
   I1 => x35_out_31,
   I2 => x35_out_1,
   I3 => W_53_15_i_10_n_0,
   I4 => W_53_15_i_11_n_0,
   O => W_53_15_i_2_n_0
);
W_53_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x35_out_23,
   I1 => x35_out_30,
   I2 => x35_out_0,
   I3 => W_53_15_i_12_n_0,
   I4 => W_53_15_i_13_n_0,
   O => W_53_15_i_3_n_0
);
W_53_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x35_out_22,
   I1 => x35_out_29,
   I2 => x35_out_31,
   I3 => W_53_15_i_14_n_0,
   I4 => W_53_15_i_15_n_0,
   O => W_53_15_i_4_n_0
);
W_53_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x35_out_21,
   I1 => x35_out_28,
   I2 => x35_out_30,
   I3 => W_53_15_i_16_n_0,
   I4 => W_53_15_i_17_n_0,
   O => W_53_15_i_5_n_0
);
W_53_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_53_15_i_2_n_0,
   I1 => W_53_19_i_16_n_0,
   I2 => x35_out_25,
   I3 => x35_out_0,
   I4 => x35_out_2,
   I5 => W_53_19_i_17_n_0,
   O => W_53_15_i_6_n_0
);
W_53_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_53_15_i_3_n_0,
   I1 => W_53_15_i_10_n_0,
   I2 => x35_out_24,
   I3 => x35_out_31,
   I4 => x35_out_1,
   I5 => W_53_15_i_11_n_0,
   O => W_53_15_i_7_n_0
);
W_53_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_53_15_i_4_n_0,
   I1 => W_53_15_i_12_n_0,
   I2 => x35_out_23,
   I3 => x35_out_30,
   I4 => x35_out_0,
   I5 => W_53_15_i_13_n_0,
   O => W_53_15_i_8_n_0
);
W_53_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_53_15_i_5_n_0,
   I1 => W_53_15_i_14_n_0,
   I2 => x35_out_22,
   I3 => x35_out_29,
   I4 => x35_out_31,
   I5 => W_53_15_i_15_n_0,
   O => W_53_15_i_9_n_0
);
W_53_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x77_out_18,
   I1 => x50_out_18,
   I2 => x74_out_4,
   I3 => x74_out_25,
   I4 => x74_out_21,
   O => W_53_19_i_10_n_0
);
W_53_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x50_out_17,
   I1 => x74_out_20,
   I2 => x74_out_24,
   I3 => x74_out_3,
   I4 => x77_out_17,
   O => W_53_19_i_11_n_0
);
W_53_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x77_out_17,
   I1 => x50_out_17,
   I2 => x74_out_3,
   I3 => x74_out_24,
   I4 => x74_out_20,
   O => W_53_19_i_12_n_0
);
W_53_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x50_out_16,
   I1 => x74_out_19,
   I2 => x74_out_23,
   I3 => x74_out_2,
   I4 => x77_out_16,
   O => W_53_19_i_13_n_0
);
W_53_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x77_out_16,
   I1 => x50_out_16,
   I2 => x74_out_2,
   I3 => x74_out_23,
   I4 => x74_out_19,
   O => W_53_19_i_14_n_0
);
W_53_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x50_out_15,
   I1 => x74_out_18,
   I2 => x74_out_22,
   I3 => x74_out_1,
   I4 => x77_out_15,
   O => W_53_19_i_15_n_0
);
W_53_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x77_out_15,
   I1 => x50_out_15,
   I2 => x74_out_1,
   I3 => x74_out_22,
   I4 => x74_out_18,
   O => W_53_19_i_16_n_0
);
W_53_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x50_out_14,
   I1 => x74_out_17,
   I2 => x74_out_21,
   I3 => x74_out_0,
   I4 => x77_out_14,
   O => W_53_19_i_17_n_0
);
W_53_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x35_out_28,
   I1 => x35_out_3,
   I2 => x35_out_5,
   I3 => W_53_19_i_10_n_0,
   I4 => W_53_19_i_11_n_0,
   O => W_53_19_i_2_n_0
);
W_53_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x35_out_27,
   I1 => x35_out_2,
   I2 => x35_out_4,
   I3 => W_53_19_i_12_n_0,
   I4 => W_53_19_i_13_n_0,
   O => W_53_19_i_3_n_0
);
W_53_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x35_out_26,
   I1 => x35_out_1,
   I2 => x35_out_3,
   I3 => W_53_19_i_14_n_0,
   I4 => W_53_19_i_15_n_0,
   O => W_53_19_i_4_n_0
);
W_53_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x35_out_25,
   I1 => x35_out_0,
   I2 => x35_out_2,
   I3 => W_53_19_i_16_n_0,
   I4 => W_53_19_i_17_n_0,
   O => W_53_19_i_5_n_0
);
W_53_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_53_19_i_2_n_0,
   I1 => W_53_23_i_16_n_0,
   I2 => x35_out_29,
   I3 => x35_out_4,
   I4 => x35_out_6,
   I5 => W_53_23_i_17_n_0,
   O => W_53_19_i_6_n_0
);
W_53_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_53_19_i_3_n_0,
   I1 => W_53_19_i_10_n_0,
   I2 => x35_out_28,
   I3 => x35_out_3,
   I4 => x35_out_5,
   I5 => W_53_19_i_11_n_0,
   O => W_53_19_i_7_n_0
);
W_53_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_53_19_i_4_n_0,
   I1 => W_53_19_i_12_n_0,
   I2 => x35_out_27,
   I3 => x35_out_2,
   I4 => x35_out_4,
   I5 => W_53_19_i_13_n_0,
   O => W_53_19_i_8_n_0
);
W_53_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_53_19_i_5_n_0,
   I1 => W_53_19_i_14_n_0,
   I2 => x35_out_26,
   I3 => x35_out_1,
   I4 => x35_out_3,
   I5 => W_53_19_i_15_n_0,
   O => W_53_19_i_9_n_0
);
W_53_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x77_out_22,
   I1 => x50_out_22,
   I2 => x74_out_8,
   I3 => x74_out_29,
   I4 => x74_out_25,
   O => W_53_23_i_10_n_0
);
W_53_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x50_out_21,
   I1 => x74_out_24,
   I2 => x74_out_28,
   I3 => x74_out_7,
   I4 => x77_out_21,
   O => W_53_23_i_11_n_0
);
W_53_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x77_out_21,
   I1 => x50_out_21,
   I2 => x74_out_7,
   I3 => x74_out_28,
   I4 => x74_out_24,
   O => W_53_23_i_12_n_0
);
W_53_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x50_out_20,
   I1 => x74_out_23,
   I2 => x74_out_27,
   I3 => x74_out_6,
   I4 => x77_out_20,
   O => W_53_23_i_13_n_0
);
W_53_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x77_out_20,
   I1 => x50_out_20,
   I2 => x74_out_6,
   I3 => x74_out_27,
   I4 => x74_out_23,
   O => W_53_23_i_14_n_0
);
W_53_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x50_out_19,
   I1 => x74_out_22,
   I2 => x74_out_26,
   I3 => x74_out_5,
   I4 => x77_out_19,
   O => W_53_23_i_15_n_0
);
W_53_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x77_out_19,
   I1 => x50_out_19,
   I2 => x74_out_5,
   I3 => x74_out_26,
   I4 => x74_out_22,
   O => W_53_23_i_16_n_0
);
W_53_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x50_out_18,
   I1 => x74_out_21,
   I2 => x74_out_25,
   I3 => x74_out_4,
   I4 => x77_out_18,
   O => W_53_23_i_17_n_0
);
W_53_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x35_out_7,
   I1 => x35_out_9,
   I2 => W_53_23_i_10_n_0,
   I3 => W_53_23_i_11_n_0,
   O => W_53_23_i_2_n_0
);
W_53_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x35_out_31,
   I1 => x35_out_6,
   I2 => x35_out_8,
   I3 => W_53_23_i_12_n_0,
   I4 => W_53_23_i_13_n_0,
   O => W_53_23_i_3_n_0
);
W_53_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x35_out_30,
   I1 => x35_out_5,
   I2 => x35_out_7,
   I3 => W_53_23_i_14_n_0,
   I4 => W_53_23_i_15_n_0,
   O => W_53_23_i_4_n_0
);
W_53_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x35_out_29,
   I1 => x35_out_4,
   I2 => x35_out_6,
   I3 => W_53_23_i_16_n_0,
   I4 => W_53_23_i_17_n_0,
   O => W_53_23_i_5_n_0
);
W_53_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x35_out_8,
   I1 => x35_out_10,
   I2 => W_53_27_i_16_n_0,
   I3 => W_53_27_i_17_n_0,
   I4 => W_53_23_i_2_n_0,
   O => W_53_23_i_6_n_0
);
W_53_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x35_out_7,
   I1 => x35_out_9,
   I2 => W_53_23_i_10_n_0,
   I3 => W_53_23_i_11_n_0,
   I4 => W_53_23_i_3_n_0,
   O => W_53_23_i_7_n_0
);
W_53_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_53_23_i_4_n_0,
   I1 => W_53_23_i_12_n_0,
   I2 => x35_out_31,
   I3 => x35_out_6,
   I4 => x35_out_8,
   I5 => W_53_23_i_13_n_0,
   O => W_53_23_i_8_n_0
);
W_53_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_53_23_i_5_n_0,
   I1 => W_53_23_i_14_n_0,
   I2 => x35_out_30,
   I3 => x35_out_5,
   I4 => x35_out_7,
   I5 => W_53_23_i_15_n_0,
   O => W_53_23_i_9_n_0
);
W_53_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x77_out_26,
   I1 => x50_out_26,
   I2 => x74_out_12,
   I3 => x74_out_1,
   I4 => x74_out_29,
   O => W_53_27_i_10_n_0
);
W_53_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x50_out_25,
   I1 => x74_out_28,
   I2 => x74_out_0,
   I3 => x74_out_11,
   I4 => x77_out_25,
   O => W_53_27_i_11_n_0
);
W_53_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x77_out_25,
   I1 => x50_out_25,
   I2 => x74_out_11,
   I3 => x74_out_0,
   I4 => x74_out_28,
   O => W_53_27_i_12_n_0
);
W_53_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x50_out_24,
   I1 => x74_out_27,
   I2 => x74_out_31,
   I3 => x74_out_10,
   I4 => x77_out_24,
   O => W_53_27_i_13_n_0
);
W_53_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x77_out_24,
   I1 => x50_out_24,
   I2 => x74_out_10,
   I3 => x74_out_31,
   I4 => x74_out_27,
   O => W_53_27_i_14_n_0
);
W_53_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x50_out_23,
   I1 => x74_out_26,
   I2 => x74_out_30,
   I3 => x74_out_9,
   I4 => x77_out_23,
   O => W_53_27_i_15_n_0
);
W_53_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x77_out_23,
   I1 => x50_out_23,
   I2 => x74_out_9,
   I3 => x74_out_30,
   I4 => x74_out_26,
   O => W_53_27_i_16_n_0
);
W_53_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x50_out_22,
   I1 => x74_out_25,
   I2 => x74_out_29,
   I3 => x74_out_8,
   I4 => x77_out_22,
   O => W_53_27_i_17_n_0
);
W_53_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x35_out_11,
   I1 => x35_out_13,
   I2 => W_53_27_i_10_n_0,
   I3 => W_53_27_i_11_n_0,
   O => W_53_27_i_2_n_0
);
W_53_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x35_out_10,
   I1 => x35_out_12,
   I2 => W_53_27_i_12_n_0,
   I3 => W_53_27_i_13_n_0,
   O => W_53_27_i_3_n_0
);
W_53_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x35_out_9,
   I1 => x35_out_11,
   I2 => W_53_27_i_14_n_0,
   I3 => W_53_27_i_15_n_0,
   O => W_53_27_i_4_n_0
);
W_53_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x35_out_8,
   I1 => x35_out_10,
   I2 => W_53_27_i_16_n_0,
   I3 => W_53_27_i_17_n_0,
   O => W_53_27_i_5_n_0
);
W_53_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x35_out_12,
   I1 => x35_out_14,
   I2 => W_53_31_i_13_n_0,
   I3 => W_53_31_i_14_n_0,
   I4 => W_53_27_i_2_n_0,
   O => W_53_27_i_6_n_0
);
W_53_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x35_out_11,
   I1 => x35_out_13,
   I2 => W_53_27_i_10_n_0,
   I3 => W_53_27_i_11_n_0,
   I4 => W_53_27_i_3_n_0,
   O => W_53_27_i_7_n_0
);
W_53_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x35_out_10,
   I1 => x35_out_12,
   I2 => W_53_27_i_12_n_0,
   I3 => W_53_27_i_13_n_0,
   I4 => W_53_27_i_4_n_0,
   O => W_53_27_i_8_n_0
);
W_53_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x35_out_9,
   I1 => x35_out_11,
   I2 => W_53_27_i_14_n_0,
   I3 => W_53_27_i_15_n_0,
   I4 => W_53_27_i_5_n_0,
   O => W_53_27_i_9_n_0
);
W_53_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x50_out_28,
   I1 => x74_out_31,
   I2 => x74_out_3,
   I3 => x74_out_14,
   I4 => x77_out_28,
   O => W_53_31_i_10_n_0
);
W_53_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x77_out_28,
   I1 => x50_out_28,
   I2 => x74_out_14,
   I3 => x74_out_3,
   I4 => x74_out_31,
   O => W_53_31_i_11_n_0
);
W_53_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x50_out_27,
   I1 => x74_out_30,
   I2 => x74_out_2,
   I3 => x74_out_13,
   I4 => x77_out_27,
   O => W_53_31_i_12_n_0
);
W_53_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x77_out_27,
   I1 => x50_out_27,
   I2 => x74_out_13,
   I3 => x74_out_2,
   I4 => x74_out_30,
   O => W_53_31_i_13_n_0
);
W_53_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x50_out_26,
   I1 => x74_out_29,
   I2 => x74_out_1,
   I3 => x74_out_12,
   I4 => x77_out_26,
   O => W_53_31_i_14_n_0
);
W_53_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x50_out_29,
   I1 => x74_out_4,
   I2 => x74_out_15,
   I3 => x77_out_29,
   O => W_53_31_i_15_n_0
);
W_53_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x35_out_17,
   I1 => x35_out_15,
   O => SIGMA_LCASE_191_out_0_30
);
W_53_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => x74_out_6,
   I1 => x74_out_17,
   I2 => x50_out_31,
   I3 => x77_out_31,
   I4 => x35_out_16,
   I5 => x35_out_18,
   O => W_53_31_i_17_n_0
);
W_53_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x74_out_16,
   I1 => x74_out_5,
   O => SIGMA_LCASE_087_out_30
);
W_53_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x77_out_30,
   I1 => x50_out_30,
   I2 => x74_out_16,
   I3 => x74_out_5,
   O => W_53_31_i_19_n_0
);
W_53_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x35_out_14,
   I1 => x35_out_16,
   I2 => W_53_31_i_9_n_0,
   I3 => W_53_31_i_10_n_0,
   O => W_53_31_i_2_n_0
);
W_53_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x35_out_13,
   I1 => x35_out_15,
   I2 => W_53_31_i_11_n_0,
   I3 => W_53_31_i_12_n_0,
   O => W_53_31_i_3_n_0
);
W_53_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x35_out_12,
   I1 => x35_out_14,
   I2 => W_53_31_i_13_n_0,
   I3 => W_53_31_i_14_n_0,
   O => W_53_31_i_4_n_0
);
W_53_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_53_31_i_15_n_0,
   I1 => SIGMA_LCASE_191_out_0_30,
   I2 => W_53_31_i_17_n_0,
   I3 => x50_out_30,
   I4 => SIGMA_LCASE_087_out_30,
   I5 => x77_out_30,
   O => W_53_31_i_5_n_0
);
W_53_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_53_31_i_2_n_0,
   I1 => W_53_31_i_19_n_0,
   I2 => x35_out_15,
   I3 => x35_out_17,
   I4 => W_53_31_i_15_n_0,
   O => W_53_31_i_6_n_0
);
W_53_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x35_out_14,
   I1 => x35_out_16,
   I2 => W_53_31_i_9_n_0,
   I3 => W_53_31_i_10_n_0,
   I4 => W_53_31_i_3_n_0,
   O => W_53_31_i_7_n_0
);
W_53_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x35_out_13,
   I1 => x35_out_15,
   I2 => W_53_31_i_11_n_0,
   I3 => W_53_31_i_12_n_0,
   I4 => W_53_31_i_4_n_0,
   O => W_53_31_i_8_n_0
);
W_53_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x77_out_29,
   I1 => x50_out_29,
   I2 => x74_out_15,
   I3 => x74_out_4,
   O => W_53_31_i_9_n_0
);
W_53_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x77_out_2,
   I1 => x50_out_2,
   I2 => x74_out_20,
   I3 => x74_out_9,
   I4 => x74_out_5,
   O => W_53_3_i_10_n_0
);
W_53_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x50_out_1,
   I1 => x74_out_4,
   I2 => x74_out_8,
   I3 => x74_out_19,
   I4 => x77_out_1,
   O => W_53_3_i_11_n_0
);
W_53_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x74_out_19,
   I1 => x74_out_8,
   I2 => x74_out_4,
   O => SIGMA_LCASE_087_out_1
);
W_53_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x35_out_21,
   I1 => x35_out_19,
   I2 => x35_out_12,
   O => SIGMA_LCASE_191_out_0_2
);
W_53_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x35_out_20,
   I1 => x35_out_18,
   I2 => x35_out_11,
   O => SIGMA_LCASE_191_out_1
);
W_53_3_i_15 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x77_out_1,
   I1 => x50_out_1,
   I2 => x74_out_19,
   I3 => x74_out_8,
   I4 => x74_out_4,
   O => W_53_3_i_15_n_0
);
W_53_3_i_16 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x74_out_18,
   I1 => x74_out_7,
   I2 => x74_out_3,
   O => SIGMA_LCASE_087_out_0
);
W_53_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x35_out_12,
   I1 => x35_out_19,
   I2 => x35_out_21,
   I3 => W_53_3_i_10_n_0,
   I4 => W_53_3_i_11_n_0,
   O => W_53_3_i_2_n_0
);
W_53_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_53_3_i_11_n_0,
   I1 => x35_out_21,
   I2 => x35_out_19,
   I3 => x35_out_12,
   I4 => W_53_3_i_10_n_0,
   O => W_53_3_i_3_n_0
);
W_53_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_087_out_1,
   I1 => x50_out_1,
   I2 => x77_out_1,
   I3 => x35_out_11,
   I4 => x35_out_18,
   I5 => x35_out_20,
   O => W_53_3_i_4_n_0
);
W_53_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x77_out_0,
   I1 => x50_out_0,
   I2 => x74_out_18,
   I3 => x74_out_7,
   I4 => x74_out_3,
   O => W_53_3_i_5_n_0
);
W_53_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_53_3_i_2_n_0,
   I1 => W_53_7_i_16_n_0,
   I2 => x35_out_13,
   I3 => x35_out_20,
   I4 => x35_out_22,
   I5 => W_53_7_i_17_n_0,
   O => W_53_3_i_6_n_0
);
W_53_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_53_3_i_10_n_0,
   I1 => SIGMA_LCASE_191_out_0_2,
   I2 => x77_out_1,
   I3 => x50_out_1,
   I4 => SIGMA_LCASE_087_out_1,
   I5 => SIGMA_LCASE_191_out_1,
   O => W_53_3_i_7_n_0
);
W_53_3_i_8 : LUT5
  generic map(
   INIT => X"99969666"
  )
 port map (
   I0 => SIGMA_LCASE_191_out_1,
   I1 => W_53_3_i_15_n_0,
   I2 => x77_out_0,
   I3 => SIGMA_LCASE_087_out_0,
   I4 => x50_out_0,
   O => W_53_3_i_8_n_0
);
W_53_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_53_3_i_5_n_0,
   I1 => x35_out_10,
   I2 => x35_out_17,
   I3 => x35_out_19,
   O => W_53_3_i_9_n_0
);
W_53_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x77_out_6,
   I1 => x50_out_6,
   I2 => x74_out_24,
   I3 => x74_out_13,
   I4 => x74_out_9,
   O => W_53_7_i_10_n_0
);
W_53_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x50_out_5,
   I1 => x74_out_8,
   I2 => x74_out_12,
   I3 => x74_out_23,
   I4 => x77_out_5,
   O => W_53_7_i_11_n_0
);
W_53_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x77_out_5,
   I1 => x50_out_5,
   I2 => x74_out_23,
   I3 => x74_out_12,
   I4 => x74_out_8,
   O => W_53_7_i_12_n_0
);
W_53_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x50_out_4,
   I1 => x74_out_7,
   I2 => x74_out_11,
   I3 => x74_out_22,
   I4 => x77_out_4,
   O => W_53_7_i_13_n_0
);
W_53_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x77_out_4,
   I1 => x50_out_4,
   I2 => x74_out_22,
   I3 => x74_out_11,
   I4 => x74_out_7,
   O => W_53_7_i_14_n_0
);
W_53_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x50_out_3,
   I1 => x74_out_6,
   I2 => x74_out_10,
   I3 => x74_out_21,
   I4 => x77_out_3,
   O => W_53_7_i_15_n_0
);
W_53_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x77_out_3,
   I1 => x50_out_3,
   I2 => x74_out_21,
   I3 => x74_out_10,
   I4 => x74_out_6,
   O => W_53_7_i_16_n_0
);
W_53_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x50_out_2,
   I1 => x74_out_5,
   I2 => x74_out_9,
   I3 => x74_out_20,
   I4 => x77_out_2,
   O => W_53_7_i_17_n_0
);
W_53_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x35_out_16,
   I1 => x35_out_23,
   I2 => x35_out_25,
   I3 => W_53_7_i_10_n_0,
   I4 => W_53_7_i_11_n_0,
   O => W_53_7_i_2_n_0
);
W_53_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x35_out_15,
   I1 => x35_out_22,
   I2 => x35_out_24,
   I3 => W_53_7_i_12_n_0,
   I4 => W_53_7_i_13_n_0,
   O => W_53_7_i_3_n_0
);
W_53_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x35_out_14,
   I1 => x35_out_21,
   I2 => x35_out_23,
   I3 => W_53_7_i_14_n_0,
   I4 => W_53_7_i_15_n_0,
   O => W_53_7_i_4_n_0
);
W_53_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x35_out_13,
   I1 => x35_out_20,
   I2 => x35_out_22,
   I3 => W_53_7_i_16_n_0,
   I4 => W_53_7_i_17_n_0,
   O => W_53_7_i_5_n_0
);
W_53_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_53_7_i_2_n_0,
   I1 => W_53_11_i_16_n_0,
   I2 => x35_out_17,
   I3 => x35_out_24,
   I4 => x35_out_26,
   I5 => W_53_11_i_17_n_0,
   O => W_53_7_i_6_n_0
);
W_53_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_53_7_i_3_n_0,
   I1 => W_53_7_i_10_n_0,
   I2 => x35_out_16,
   I3 => x35_out_23,
   I4 => x35_out_25,
   I5 => W_53_7_i_11_n_0,
   O => W_53_7_i_7_n_0
);
W_53_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_53_7_i_4_n_0,
   I1 => W_53_7_i_12_n_0,
   I2 => x35_out_15,
   I3 => x35_out_22,
   I4 => x35_out_24,
   I5 => W_53_7_i_13_n_0,
   O => W_53_7_i_8_n_0
);
W_53_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_53_7_i_5_n_0,
   I1 => W_53_7_i_14_n_0,
   I2 => x35_out_14,
   I3 => x35_out_21,
   I4 => x35_out_23,
   I5 => W_53_7_i_15_n_0,
   O => W_53_7_i_9_n_0
);
W_54_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x74_out_10,
   I1 => x47_out_10,
   I2 => x71_out_28,
   I3 => x71_out_17,
   I4 => x71_out_13,
   O => W_54_11_i_10_n_0
);
W_54_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x47_out_9,
   I1 => x71_out_12,
   I2 => x71_out_16,
   I3 => x71_out_27,
   I4 => x74_out_9,
   O => W_54_11_i_11_n_0
);
W_54_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x74_out_9,
   I1 => x47_out_9,
   I2 => x71_out_27,
   I3 => x71_out_16,
   I4 => x71_out_12,
   O => W_54_11_i_12_n_0
);
W_54_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x47_out_8,
   I1 => x71_out_11,
   I2 => x71_out_15,
   I3 => x71_out_26,
   I4 => x74_out_8,
   O => W_54_11_i_13_n_0
);
W_54_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x74_out_8,
   I1 => x47_out_8,
   I2 => x71_out_26,
   I3 => x71_out_15,
   I4 => x71_out_11,
   O => W_54_11_i_14_n_0
);
W_54_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x47_out_7,
   I1 => x71_out_10,
   I2 => x71_out_14,
   I3 => x71_out_25,
   I4 => x74_out_7,
   O => W_54_11_i_15_n_0
);
W_54_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x74_out_7,
   I1 => x47_out_7,
   I2 => x71_out_25,
   I3 => x71_out_14,
   I4 => x71_out_10,
   O => W_54_11_i_16_n_0
);
W_54_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x47_out_6,
   I1 => x71_out_9,
   I2 => x71_out_13,
   I3 => x71_out_24,
   I4 => x74_out_6,
   O => W_54_11_i_17_n_0
);
W_54_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x32_out_20,
   I1 => x32_out_27,
   I2 => x32_out_29,
   I3 => W_54_11_i_10_n_0,
   I4 => W_54_11_i_11_n_0,
   O => W_54_11_i_2_n_0
);
W_54_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x32_out_19,
   I1 => x32_out_26,
   I2 => x32_out_28,
   I3 => W_54_11_i_12_n_0,
   I4 => W_54_11_i_13_n_0,
   O => W_54_11_i_3_n_0
);
W_54_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x32_out_18,
   I1 => x32_out_25,
   I2 => x32_out_27,
   I3 => W_54_11_i_14_n_0,
   I4 => W_54_11_i_15_n_0,
   O => W_54_11_i_4_n_0
);
W_54_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x32_out_17,
   I1 => x32_out_24,
   I2 => x32_out_26,
   I3 => W_54_11_i_16_n_0,
   I4 => W_54_11_i_17_n_0,
   O => W_54_11_i_5_n_0
);
W_54_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_54_11_i_2_n_0,
   I1 => W_54_15_i_16_n_0,
   I2 => x32_out_21,
   I3 => x32_out_28,
   I4 => x32_out_30,
   I5 => W_54_15_i_17_n_0,
   O => W_54_11_i_6_n_0
);
W_54_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_54_11_i_3_n_0,
   I1 => W_54_11_i_10_n_0,
   I2 => x32_out_20,
   I3 => x32_out_27,
   I4 => x32_out_29,
   I5 => W_54_11_i_11_n_0,
   O => W_54_11_i_7_n_0
);
W_54_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_54_11_i_4_n_0,
   I1 => W_54_11_i_12_n_0,
   I2 => x32_out_19,
   I3 => x32_out_26,
   I4 => x32_out_28,
   I5 => W_54_11_i_13_n_0,
   O => W_54_11_i_8_n_0
);
W_54_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_54_11_i_5_n_0,
   I1 => W_54_11_i_14_n_0,
   I2 => x32_out_18,
   I3 => x32_out_25,
   I4 => x32_out_27,
   I5 => W_54_11_i_15_n_0,
   O => W_54_11_i_9_n_0
);
W_54_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x74_out_14,
   I1 => x47_out_14,
   I2 => x71_out_0,
   I3 => x71_out_21,
   I4 => x71_out_17,
   O => W_54_15_i_10_n_0
);
W_54_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x47_out_13,
   I1 => x71_out_16,
   I2 => x71_out_20,
   I3 => x71_out_31,
   I4 => x74_out_13,
   O => W_54_15_i_11_n_0
);
W_54_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x74_out_13,
   I1 => x47_out_13,
   I2 => x71_out_31,
   I3 => x71_out_20,
   I4 => x71_out_16,
   O => W_54_15_i_12_n_0
);
W_54_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x47_out_12,
   I1 => x71_out_15,
   I2 => x71_out_19,
   I3 => x71_out_30,
   I4 => x74_out_12,
   O => W_54_15_i_13_n_0
);
W_54_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x74_out_12,
   I1 => x47_out_12,
   I2 => x71_out_30,
   I3 => x71_out_19,
   I4 => x71_out_15,
   O => W_54_15_i_14_n_0
);
W_54_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x47_out_11,
   I1 => x71_out_14,
   I2 => x71_out_18,
   I3 => x71_out_29,
   I4 => x74_out_11,
   O => W_54_15_i_15_n_0
);
W_54_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x74_out_11,
   I1 => x47_out_11,
   I2 => x71_out_29,
   I3 => x71_out_18,
   I4 => x71_out_14,
   O => W_54_15_i_16_n_0
);
W_54_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x47_out_10,
   I1 => x71_out_13,
   I2 => x71_out_17,
   I3 => x71_out_28,
   I4 => x74_out_10,
   O => W_54_15_i_17_n_0
);
W_54_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x32_out_24,
   I1 => x32_out_31,
   I2 => x32_out_1,
   I3 => W_54_15_i_10_n_0,
   I4 => W_54_15_i_11_n_0,
   O => W_54_15_i_2_n_0
);
W_54_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x32_out_23,
   I1 => x32_out_30,
   I2 => x32_out_0,
   I3 => W_54_15_i_12_n_0,
   I4 => W_54_15_i_13_n_0,
   O => W_54_15_i_3_n_0
);
W_54_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x32_out_22,
   I1 => x32_out_29,
   I2 => x32_out_31,
   I3 => W_54_15_i_14_n_0,
   I4 => W_54_15_i_15_n_0,
   O => W_54_15_i_4_n_0
);
W_54_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x32_out_21,
   I1 => x32_out_28,
   I2 => x32_out_30,
   I3 => W_54_15_i_16_n_0,
   I4 => W_54_15_i_17_n_0,
   O => W_54_15_i_5_n_0
);
W_54_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_54_15_i_2_n_0,
   I1 => W_54_19_i_16_n_0,
   I2 => x32_out_25,
   I3 => x32_out_0,
   I4 => x32_out_2,
   I5 => W_54_19_i_17_n_0,
   O => W_54_15_i_6_n_0
);
W_54_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_54_15_i_3_n_0,
   I1 => W_54_15_i_10_n_0,
   I2 => x32_out_24,
   I3 => x32_out_31,
   I4 => x32_out_1,
   I5 => W_54_15_i_11_n_0,
   O => W_54_15_i_7_n_0
);
W_54_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_54_15_i_4_n_0,
   I1 => W_54_15_i_12_n_0,
   I2 => x32_out_23,
   I3 => x32_out_30,
   I4 => x32_out_0,
   I5 => W_54_15_i_13_n_0,
   O => W_54_15_i_8_n_0
);
W_54_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_54_15_i_5_n_0,
   I1 => W_54_15_i_14_n_0,
   I2 => x32_out_22,
   I3 => x32_out_29,
   I4 => x32_out_31,
   I5 => W_54_15_i_15_n_0,
   O => W_54_15_i_9_n_0
);
W_54_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x74_out_18,
   I1 => x47_out_18,
   I2 => x71_out_4,
   I3 => x71_out_25,
   I4 => x71_out_21,
   O => W_54_19_i_10_n_0
);
W_54_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x47_out_17,
   I1 => x71_out_20,
   I2 => x71_out_24,
   I3 => x71_out_3,
   I4 => x74_out_17,
   O => W_54_19_i_11_n_0
);
W_54_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x74_out_17,
   I1 => x47_out_17,
   I2 => x71_out_3,
   I3 => x71_out_24,
   I4 => x71_out_20,
   O => W_54_19_i_12_n_0
);
W_54_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x47_out_16,
   I1 => x71_out_19,
   I2 => x71_out_23,
   I3 => x71_out_2,
   I4 => x74_out_16,
   O => W_54_19_i_13_n_0
);
W_54_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x74_out_16,
   I1 => x47_out_16,
   I2 => x71_out_2,
   I3 => x71_out_23,
   I4 => x71_out_19,
   O => W_54_19_i_14_n_0
);
W_54_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x47_out_15,
   I1 => x71_out_18,
   I2 => x71_out_22,
   I3 => x71_out_1,
   I4 => x74_out_15,
   O => W_54_19_i_15_n_0
);
W_54_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x74_out_15,
   I1 => x47_out_15,
   I2 => x71_out_1,
   I3 => x71_out_22,
   I4 => x71_out_18,
   O => W_54_19_i_16_n_0
);
W_54_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x47_out_14,
   I1 => x71_out_17,
   I2 => x71_out_21,
   I3 => x71_out_0,
   I4 => x74_out_14,
   O => W_54_19_i_17_n_0
);
W_54_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x32_out_28,
   I1 => x32_out_3,
   I2 => x32_out_5,
   I3 => W_54_19_i_10_n_0,
   I4 => W_54_19_i_11_n_0,
   O => W_54_19_i_2_n_0
);
W_54_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x32_out_27,
   I1 => x32_out_2,
   I2 => x32_out_4,
   I3 => W_54_19_i_12_n_0,
   I4 => W_54_19_i_13_n_0,
   O => W_54_19_i_3_n_0
);
W_54_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x32_out_26,
   I1 => x32_out_1,
   I2 => x32_out_3,
   I3 => W_54_19_i_14_n_0,
   I4 => W_54_19_i_15_n_0,
   O => W_54_19_i_4_n_0
);
W_54_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x32_out_25,
   I1 => x32_out_0,
   I2 => x32_out_2,
   I3 => W_54_19_i_16_n_0,
   I4 => W_54_19_i_17_n_0,
   O => W_54_19_i_5_n_0
);
W_54_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_54_19_i_2_n_0,
   I1 => W_54_23_i_16_n_0,
   I2 => x32_out_29,
   I3 => x32_out_4,
   I4 => x32_out_6,
   I5 => W_54_23_i_17_n_0,
   O => W_54_19_i_6_n_0
);
W_54_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_54_19_i_3_n_0,
   I1 => W_54_19_i_10_n_0,
   I2 => x32_out_28,
   I3 => x32_out_3,
   I4 => x32_out_5,
   I5 => W_54_19_i_11_n_0,
   O => W_54_19_i_7_n_0
);
W_54_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_54_19_i_4_n_0,
   I1 => W_54_19_i_12_n_0,
   I2 => x32_out_27,
   I3 => x32_out_2,
   I4 => x32_out_4,
   I5 => W_54_19_i_13_n_0,
   O => W_54_19_i_8_n_0
);
W_54_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_54_19_i_5_n_0,
   I1 => W_54_19_i_14_n_0,
   I2 => x32_out_26,
   I3 => x32_out_1,
   I4 => x32_out_3,
   I5 => W_54_19_i_15_n_0,
   O => W_54_19_i_9_n_0
);
W_54_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x74_out_22,
   I1 => x47_out_22,
   I2 => x71_out_8,
   I3 => x71_out_29,
   I4 => x71_out_25,
   O => W_54_23_i_10_n_0
);
W_54_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x47_out_21,
   I1 => x71_out_24,
   I2 => x71_out_28,
   I3 => x71_out_7,
   I4 => x74_out_21,
   O => W_54_23_i_11_n_0
);
W_54_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x74_out_21,
   I1 => x47_out_21,
   I2 => x71_out_7,
   I3 => x71_out_28,
   I4 => x71_out_24,
   O => W_54_23_i_12_n_0
);
W_54_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x47_out_20,
   I1 => x71_out_23,
   I2 => x71_out_27,
   I3 => x71_out_6,
   I4 => x74_out_20,
   O => W_54_23_i_13_n_0
);
W_54_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x74_out_20,
   I1 => x47_out_20,
   I2 => x71_out_6,
   I3 => x71_out_27,
   I4 => x71_out_23,
   O => W_54_23_i_14_n_0
);
W_54_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x47_out_19,
   I1 => x71_out_22,
   I2 => x71_out_26,
   I3 => x71_out_5,
   I4 => x74_out_19,
   O => W_54_23_i_15_n_0
);
W_54_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x74_out_19,
   I1 => x47_out_19,
   I2 => x71_out_5,
   I3 => x71_out_26,
   I4 => x71_out_22,
   O => W_54_23_i_16_n_0
);
W_54_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x47_out_18,
   I1 => x71_out_21,
   I2 => x71_out_25,
   I3 => x71_out_4,
   I4 => x74_out_18,
   O => W_54_23_i_17_n_0
);
W_54_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x32_out_7,
   I1 => x32_out_9,
   I2 => W_54_23_i_10_n_0,
   I3 => W_54_23_i_11_n_0,
   O => W_54_23_i_2_n_0
);
W_54_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x32_out_31,
   I1 => x32_out_6,
   I2 => x32_out_8,
   I3 => W_54_23_i_12_n_0,
   I4 => W_54_23_i_13_n_0,
   O => W_54_23_i_3_n_0
);
W_54_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x32_out_30,
   I1 => x32_out_5,
   I2 => x32_out_7,
   I3 => W_54_23_i_14_n_0,
   I4 => W_54_23_i_15_n_0,
   O => W_54_23_i_4_n_0
);
W_54_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x32_out_29,
   I1 => x32_out_4,
   I2 => x32_out_6,
   I3 => W_54_23_i_16_n_0,
   I4 => W_54_23_i_17_n_0,
   O => W_54_23_i_5_n_0
);
W_54_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x32_out_8,
   I1 => x32_out_10,
   I2 => W_54_27_i_16_n_0,
   I3 => W_54_27_i_17_n_0,
   I4 => W_54_23_i_2_n_0,
   O => W_54_23_i_6_n_0
);
W_54_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x32_out_7,
   I1 => x32_out_9,
   I2 => W_54_23_i_10_n_0,
   I3 => W_54_23_i_11_n_0,
   I4 => W_54_23_i_3_n_0,
   O => W_54_23_i_7_n_0
);
W_54_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_54_23_i_4_n_0,
   I1 => W_54_23_i_12_n_0,
   I2 => x32_out_31,
   I3 => x32_out_6,
   I4 => x32_out_8,
   I5 => W_54_23_i_13_n_0,
   O => W_54_23_i_8_n_0
);
W_54_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_54_23_i_5_n_0,
   I1 => W_54_23_i_14_n_0,
   I2 => x32_out_30,
   I3 => x32_out_5,
   I4 => x32_out_7,
   I5 => W_54_23_i_15_n_0,
   O => W_54_23_i_9_n_0
);
W_54_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x74_out_26,
   I1 => x47_out_26,
   I2 => x71_out_12,
   I3 => x71_out_1,
   I4 => x71_out_29,
   O => W_54_27_i_10_n_0
);
W_54_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x47_out_25,
   I1 => x71_out_28,
   I2 => x71_out_0,
   I3 => x71_out_11,
   I4 => x74_out_25,
   O => W_54_27_i_11_n_0
);
W_54_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x74_out_25,
   I1 => x47_out_25,
   I2 => x71_out_11,
   I3 => x71_out_0,
   I4 => x71_out_28,
   O => W_54_27_i_12_n_0
);
W_54_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x47_out_24,
   I1 => x71_out_27,
   I2 => x71_out_31,
   I3 => x71_out_10,
   I4 => x74_out_24,
   O => W_54_27_i_13_n_0
);
W_54_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x74_out_24,
   I1 => x47_out_24,
   I2 => x71_out_10,
   I3 => x71_out_31,
   I4 => x71_out_27,
   O => W_54_27_i_14_n_0
);
W_54_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x47_out_23,
   I1 => x71_out_26,
   I2 => x71_out_30,
   I3 => x71_out_9,
   I4 => x74_out_23,
   O => W_54_27_i_15_n_0
);
W_54_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x74_out_23,
   I1 => x47_out_23,
   I2 => x71_out_9,
   I3 => x71_out_30,
   I4 => x71_out_26,
   O => W_54_27_i_16_n_0
);
W_54_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x47_out_22,
   I1 => x71_out_25,
   I2 => x71_out_29,
   I3 => x71_out_8,
   I4 => x74_out_22,
   O => W_54_27_i_17_n_0
);
W_54_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x32_out_11,
   I1 => x32_out_13,
   I2 => W_54_27_i_10_n_0,
   I3 => W_54_27_i_11_n_0,
   O => W_54_27_i_2_n_0
);
W_54_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x32_out_10,
   I1 => x32_out_12,
   I2 => W_54_27_i_12_n_0,
   I3 => W_54_27_i_13_n_0,
   O => W_54_27_i_3_n_0
);
W_54_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x32_out_9,
   I1 => x32_out_11,
   I2 => W_54_27_i_14_n_0,
   I3 => W_54_27_i_15_n_0,
   O => W_54_27_i_4_n_0
);
W_54_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x32_out_8,
   I1 => x32_out_10,
   I2 => W_54_27_i_16_n_0,
   I3 => W_54_27_i_17_n_0,
   O => W_54_27_i_5_n_0
);
W_54_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x32_out_12,
   I1 => x32_out_14,
   I2 => W_54_31_i_13_n_0,
   I3 => W_54_31_i_14_n_0,
   I4 => W_54_27_i_2_n_0,
   O => W_54_27_i_6_n_0
);
W_54_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x32_out_11,
   I1 => x32_out_13,
   I2 => W_54_27_i_10_n_0,
   I3 => W_54_27_i_11_n_0,
   I4 => W_54_27_i_3_n_0,
   O => W_54_27_i_7_n_0
);
W_54_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x32_out_10,
   I1 => x32_out_12,
   I2 => W_54_27_i_12_n_0,
   I3 => W_54_27_i_13_n_0,
   I4 => W_54_27_i_4_n_0,
   O => W_54_27_i_8_n_0
);
W_54_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x32_out_9,
   I1 => x32_out_11,
   I2 => W_54_27_i_14_n_0,
   I3 => W_54_27_i_15_n_0,
   I4 => W_54_27_i_5_n_0,
   O => W_54_27_i_9_n_0
);
W_54_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x47_out_28,
   I1 => x71_out_31,
   I2 => x71_out_3,
   I3 => x71_out_14,
   I4 => x74_out_28,
   O => W_54_31_i_10_n_0
);
W_54_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x74_out_28,
   I1 => x47_out_28,
   I2 => x71_out_14,
   I3 => x71_out_3,
   I4 => x71_out_31,
   O => W_54_31_i_11_n_0
);
W_54_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x47_out_27,
   I1 => x71_out_30,
   I2 => x71_out_2,
   I3 => x71_out_13,
   I4 => x74_out_27,
   O => W_54_31_i_12_n_0
);
W_54_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x74_out_27,
   I1 => x47_out_27,
   I2 => x71_out_13,
   I3 => x71_out_2,
   I4 => x71_out_30,
   O => W_54_31_i_13_n_0
);
W_54_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x47_out_26,
   I1 => x71_out_29,
   I2 => x71_out_1,
   I3 => x71_out_12,
   I4 => x74_out_26,
   O => W_54_31_i_14_n_0
);
W_54_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x47_out_29,
   I1 => x71_out_4,
   I2 => x71_out_15,
   I3 => x74_out_29,
   O => W_54_31_i_15_n_0
);
W_54_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x32_out_17,
   I1 => x32_out_15,
   O => SIGMA_LCASE_183_out_0_30
);
W_54_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => x71_out_6,
   I1 => x71_out_17,
   I2 => x47_out_31,
   I3 => x74_out_31,
   I4 => x32_out_16,
   I5 => x32_out_18,
   O => W_54_31_i_17_n_0
);
W_54_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x71_out_16,
   I1 => x71_out_5,
   O => SIGMA_LCASE_079_out_30
);
W_54_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x74_out_30,
   I1 => x47_out_30,
   I2 => x71_out_16,
   I3 => x71_out_5,
   O => W_54_31_i_19_n_0
);
W_54_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x32_out_14,
   I1 => x32_out_16,
   I2 => W_54_31_i_9_n_0,
   I3 => W_54_31_i_10_n_0,
   O => W_54_31_i_2_n_0
);
W_54_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x32_out_13,
   I1 => x32_out_15,
   I2 => W_54_31_i_11_n_0,
   I3 => W_54_31_i_12_n_0,
   O => W_54_31_i_3_n_0
);
W_54_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x32_out_12,
   I1 => x32_out_14,
   I2 => W_54_31_i_13_n_0,
   I3 => W_54_31_i_14_n_0,
   O => W_54_31_i_4_n_0
);
W_54_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_54_31_i_15_n_0,
   I1 => SIGMA_LCASE_183_out_0_30,
   I2 => W_54_31_i_17_n_0,
   I3 => x47_out_30,
   I4 => SIGMA_LCASE_079_out_30,
   I5 => x74_out_30,
   O => W_54_31_i_5_n_0
);
W_54_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_54_31_i_2_n_0,
   I1 => W_54_31_i_19_n_0,
   I2 => x32_out_15,
   I3 => x32_out_17,
   I4 => W_54_31_i_15_n_0,
   O => W_54_31_i_6_n_0
);
W_54_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x32_out_14,
   I1 => x32_out_16,
   I2 => W_54_31_i_9_n_0,
   I3 => W_54_31_i_10_n_0,
   I4 => W_54_31_i_3_n_0,
   O => W_54_31_i_7_n_0
);
W_54_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x32_out_13,
   I1 => x32_out_15,
   I2 => W_54_31_i_11_n_0,
   I3 => W_54_31_i_12_n_0,
   I4 => W_54_31_i_4_n_0,
   O => W_54_31_i_8_n_0
);
W_54_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x74_out_29,
   I1 => x47_out_29,
   I2 => x71_out_15,
   I3 => x71_out_4,
   O => W_54_31_i_9_n_0
);
W_54_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x74_out_2,
   I1 => x47_out_2,
   I2 => x71_out_20,
   I3 => x71_out_9,
   I4 => x71_out_5,
   O => W_54_3_i_10_n_0
);
W_54_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x47_out_1,
   I1 => x71_out_4,
   I2 => x71_out_8,
   I3 => x71_out_19,
   I4 => x74_out_1,
   O => W_54_3_i_11_n_0
);
W_54_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x71_out_19,
   I1 => x71_out_8,
   I2 => x71_out_4,
   O => SIGMA_LCASE_079_out_1
);
W_54_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x32_out_21,
   I1 => x32_out_19,
   I2 => x32_out_12,
   O => SIGMA_LCASE_183_out_0_2
);
W_54_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x32_out_20,
   I1 => x32_out_18,
   I2 => x32_out_11,
   O => SIGMA_LCASE_183_out_1
);
W_54_3_i_15 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x74_out_1,
   I1 => x47_out_1,
   I2 => x71_out_19,
   I3 => x71_out_8,
   I4 => x71_out_4,
   O => W_54_3_i_15_n_0
);
W_54_3_i_16 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x71_out_18,
   I1 => x71_out_7,
   I2 => x71_out_3,
   O => SIGMA_LCASE_079_out_0
);
W_54_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x32_out_12,
   I1 => x32_out_19,
   I2 => x32_out_21,
   I3 => W_54_3_i_10_n_0,
   I4 => W_54_3_i_11_n_0,
   O => W_54_3_i_2_n_0
);
W_54_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_54_3_i_11_n_0,
   I1 => x32_out_21,
   I2 => x32_out_19,
   I3 => x32_out_12,
   I4 => W_54_3_i_10_n_0,
   O => W_54_3_i_3_n_0
);
W_54_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_079_out_1,
   I1 => x47_out_1,
   I2 => x74_out_1,
   I3 => x32_out_11,
   I4 => x32_out_18,
   I5 => x32_out_20,
   O => W_54_3_i_4_n_0
);
W_54_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x74_out_0,
   I1 => x47_out_0,
   I2 => x71_out_18,
   I3 => x71_out_7,
   I4 => x71_out_3,
   O => W_54_3_i_5_n_0
);
W_54_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_54_3_i_2_n_0,
   I1 => W_54_7_i_16_n_0,
   I2 => x32_out_13,
   I3 => x32_out_20,
   I4 => x32_out_22,
   I5 => W_54_7_i_17_n_0,
   O => W_54_3_i_6_n_0
);
W_54_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_54_3_i_10_n_0,
   I1 => SIGMA_LCASE_183_out_0_2,
   I2 => x74_out_1,
   I3 => x47_out_1,
   I4 => SIGMA_LCASE_079_out_1,
   I5 => SIGMA_LCASE_183_out_1,
   O => W_54_3_i_7_n_0
);
W_54_3_i_8 : LUT5
  generic map(
   INIT => X"99969666"
  )
 port map (
   I0 => SIGMA_LCASE_183_out_1,
   I1 => W_54_3_i_15_n_0,
   I2 => x74_out_0,
   I3 => SIGMA_LCASE_079_out_0,
   I4 => x47_out_0,
   O => W_54_3_i_8_n_0
);
W_54_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_54_3_i_5_n_0,
   I1 => x32_out_10,
   I2 => x32_out_17,
   I3 => x32_out_19,
   O => W_54_3_i_9_n_0
);
W_54_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x74_out_6,
   I1 => x47_out_6,
   I2 => x71_out_24,
   I3 => x71_out_13,
   I4 => x71_out_9,
   O => W_54_7_i_10_n_0
);
W_54_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x47_out_5,
   I1 => x71_out_8,
   I2 => x71_out_12,
   I3 => x71_out_23,
   I4 => x74_out_5,
   O => W_54_7_i_11_n_0
);
W_54_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x74_out_5,
   I1 => x47_out_5,
   I2 => x71_out_23,
   I3 => x71_out_12,
   I4 => x71_out_8,
   O => W_54_7_i_12_n_0
);
W_54_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x47_out_4,
   I1 => x71_out_7,
   I2 => x71_out_11,
   I3 => x71_out_22,
   I4 => x74_out_4,
   O => W_54_7_i_13_n_0
);
W_54_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x74_out_4,
   I1 => x47_out_4,
   I2 => x71_out_22,
   I3 => x71_out_11,
   I4 => x71_out_7,
   O => W_54_7_i_14_n_0
);
W_54_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x47_out_3,
   I1 => x71_out_6,
   I2 => x71_out_10,
   I3 => x71_out_21,
   I4 => x74_out_3,
   O => W_54_7_i_15_n_0
);
W_54_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x74_out_3,
   I1 => x47_out_3,
   I2 => x71_out_21,
   I3 => x71_out_10,
   I4 => x71_out_6,
   O => W_54_7_i_16_n_0
);
W_54_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x47_out_2,
   I1 => x71_out_5,
   I2 => x71_out_9,
   I3 => x71_out_20,
   I4 => x74_out_2,
   O => W_54_7_i_17_n_0
);
W_54_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x32_out_16,
   I1 => x32_out_23,
   I2 => x32_out_25,
   I3 => W_54_7_i_10_n_0,
   I4 => W_54_7_i_11_n_0,
   O => W_54_7_i_2_n_0
);
W_54_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x32_out_15,
   I1 => x32_out_22,
   I2 => x32_out_24,
   I3 => W_54_7_i_12_n_0,
   I4 => W_54_7_i_13_n_0,
   O => W_54_7_i_3_n_0
);
W_54_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x32_out_14,
   I1 => x32_out_21,
   I2 => x32_out_23,
   I3 => W_54_7_i_14_n_0,
   I4 => W_54_7_i_15_n_0,
   O => W_54_7_i_4_n_0
);
W_54_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x32_out_13,
   I1 => x32_out_20,
   I2 => x32_out_22,
   I3 => W_54_7_i_16_n_0,
   I4 => W_54_7_i_17_n_0,
   O => W_54_7_i_5_n_0
);
W_54_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_54_7_i_2_n_0,
   I1 => W_54_11_i_16_n_0,
   I2 => x32_out_17,
   I3 => x32_out_24,
   I4 => x32_out_26,
   I5 => W_54_11_i_17_n_0,
   O => W_54_7_i_6_n_0
);
W_54_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_54_7_i_3_n_0,
   I1 => W_54_7_i_10_n_0,
   I2 => x32_out_16,
   I3 => x32_out_23,
   I4 => x32_out_25,
   I5 => W_54_7_i_11_n_0,
   O => W_54_7_i_7_n_0
);
W_54_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_54_7_i_4_n_0,
   I1 => W_54_7_i_12_n_0,
   I2 => x32_out_15,
   I3 => x32_out_22,
   I4 => x32_out_24,
   I5 => W_54_7_i_13_n_0,
   O => W_54_7_i_8_n_0
);
W_54_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_54_7_i_5_n_0,
   I1 => W_54_7_i_14_n_0,
   I2 => x32_out_14,
   I3 => x32_out_21,
   I4 => x32_out_23,
   I5 => W_54_7_i_15_n_0,
   O => W_54_7_i_9_n_0
);
W_55_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x71_out_10,
   I1 => x44_out_10,
   I2 => x68_out_28,
   I3 => x68_out_17,
   I4 => x68_out_13,
   O => W_55_11_i_10_n_0
);
W_55_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x44_out_9,
   I1 => x68_out_12,
   I2 => x68_out_16,
   I3 => x68_out_27,
   I4 => x71_out_9,
   O => W_55_11_i_11_n_0
);
W_55_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x71_out_9,
   I1 => x44_out_9,
   I2 => x68_out_27,
   I3 => x68_out_16,
   I4 => x68_out_12,
   O => W_55_11_i_12_n_0
);
W_55_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x44_out_8,
   I1 => x68_out_11,
   I2 => x68_out_15,
   I3 => x68_out_26,
   I4 => x71_out_8,
   O => W_55_11_i_13_n_0
);
W_55_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x71_out_8,
   I1 => x44_out_8,
   I2 => x68_out_26,
   I3 => x68_out_15,
   I4 => x68_out_11,
   O => W_55_11_i_14_n_0
);
W_55_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x44_out_7,
   I1 => x68_out_10,
   I2 => x68_out_14,
   I3 => x68_out_25,
   I4 => x71_out_7,
   O => W_55_11_i_15_n_0
);
W_55_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x71_out_7,
   I1 => x44_out_7,
   I2 => x68_out_25,
   I3 => x68_out_14,
   I4 => x68_out_10,
   O => W_55_11_i_16_n_0
);
W_55_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x44_out_6,
   I1 => x68_out_9,
   I2 => x68_out_13,
   I3 => x68_out_24,
   I4 => x71_out_6,
   O => W_55_11_i_17_n_0
);
W_55_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x29_out_20,
   I1 => x29_out_27,
   I2 => x29_out_29,
   I3 => W_55_11_i_10_n_0,
   I4 => W_55_11_i_11_n_0,
   O => W_55_11_i_2_n_0
);
W_55_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x29_out_19,
   I1 => x29_out_26,
   I2 => x29_out_28,
   I3 => W_55_11_i_12_n_0,
   I4 => W_55_11_i_13_n_0,
   O => W_55_11_i_3_n_0
);
W_55_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x29_out_18,
   I1 => x29_out_25,
   I2 => x29_out_27,
   I3 => W_55_11_i_14_n_0,
   I4 => W_55_11_i_15_n_0,
   O => W_55_11_i_4_n_0
);
W_55_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x29_out_17,
   I1 => x29_out_24,
   I2 => x29_out_26,
   I3 => W_55_11_i_16_n_0,
   I4 => W_55_11_i_17_n_0,
   O => W_55_11_i_5_n_0
);
W_55_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_55_11_i_2_n_0,
   I1 => W_55_15_i_16_n_0,
   I2 => x29_out_21,
   I3 => x29_out_28,
   I4 => x29_out_30,
   I5 => W_55_15_i_17_n_0,
   O => W_55_11_i_6_n_0
);
W_55_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_55_11_i_3_n_0,
   I1 => W_55_11_i_10_n_0,
   I2 => x29_out_20,
   I3 => x29_out_27,
   I4 => x29_out_29,
   I5 => W_55_11_i_11_n_0,
   O => W_55_11_i_7_n_0
);
W_55_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_55_11_i_4_n_0,
   I1 => W_55_11_i_12_n_0,
   I2 => x29_out_19,
   I3 => x29_out_26,
   I4 => x29_out_28,
   I5 => W_55_11_i_13_n_0,
   O => W_55_11_i_8_n_0
);
W_55_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_55_11_i_5_n_0,
   I1 => W_55_11_i_14_n_0,
   I2 => x29_out_18,
   I3 => x29_out_25,
   I4 => x29_out_27,
   I5 => W_55_11_i_15_n_0,
   O => W_55_11_i_9_n_0
);
W_55_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x71_out_14,
   I1 => x44_out_14,
   I2 => x68_out_0,
   I3 => x68_out_21,
   I4 => x68_out_17,
   O => W_55_15_i_10_n_0
);
W_55_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x44_out_13,
   I1 => x68_out_16,
   I2 => x68_out_20,
   I3 => x68_out_31,
   I4 => x71_out_13,
   O => W_55_15_i_11_n_0
);
W_55_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x71_out_13,
   I1 => x44_out_13,
   I2 => x68_out_31,
   I3 => x68_out_20,
   I4 => x68_out_16,
   O => W_55_15_i_12_n_0
);
W_55_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x44_out_12,
   I1 => x68_out_15,
   I2 => x68_out_19,
   I3 => x68_out_30,
   I4 => x71_out_12,
   O => W_55_15_i_13_n_0
);
W_55_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x71_out_12,
   I1 => x44_out_12,
   I2 => x68_out_30,
   I3 => x68_out_19,
   I4 => x68_out_15,
   O => W_55_15_i_14_n_0
);
W_55_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x44_out_11,
   I1 => x68_out_14,
   I2 => x68_out_18,
   I3 => x68_out_29,
   I4 => x71_out_11,
   O => W_55_15_i_15_n_0
);
W_55_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x71_out_11,
   I1 => x44_out_11,
   I2 => x68_out_29,
   I3 => x68_out_18,
   I4 => x68_out_14,
   O => W_55_15_i_16_n_0
);
W_55_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x44_out_10,
   I1 => x68_out_13,
   I2 => x68_out_17,
   I3 => x68_out_28,
   I4 => x71_out_10,
   O => W_55_15_i_17_n_0
);
W_55_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x29_out_24,
   I1 => x29_out_31,
   I2 => x29_out_1,
   I3 => W_55_15_i_10_n_0,
   I4 => W_55_15_i_11_n_0,
   O => W_55_15_i_2_n_0
);
W_55_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x29_out_23,
   I1 => x29_out_30,
   I2 => x29_out_0,
   I3 => W_55_15_i_12_n_0,
   I4 => W_55_15_i_13_n_0,
   O => W_55_15_i_3_n_0
);
W_55_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x29_out_22,
   I1 => x29_out_29,
   I2 => x29_out_31,
   I3 => W_55_15_i_14_n_0,
   I4 => W_55_15_i_15_n_0,
   O => W_55_15_i_4_n_0
);
W_55_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x29_out_21,
   I1 => x29_out_28,
   I2 => x29_out_30,
   I3 => W_55_15_i_16_n_0,
   I4 => W_55_15_i_17_n_0,
   O => W_55_15_i_5_n_0
);
W_55_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_55_15_i_2_n_0,
   I1 => W_55_19_i_16_n_0,
   I2 => x29_out_25,
   I3 => x29_out_0,
   I4 => x29_out_2,
   I5 => W_55_19_i_17_n_0,
   O => W_55_15_i_6_n_0
);
W_55_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_55_15_i_3_n_0,
   I1 => W_55_15_i_10_n_0,
   I2 => x29_out_24,
   I3 => x29_out_31,
   I4 => x29_out_1,
   I5 => W_55_15_i_11_n_0,
   O => W_55_15_i_7_n_0
);
W_55_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_55_15_i_4_n_0,
   I1 => W_55_15_i_12_n_0,
   I2 => x29_out_23,
   I3 => x29_out_30,
   I4 => x29_out_0,
   I5 => W_55_15_i_13_n_0,
   O => W_55_15_i_8_n_0
);
W_55_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_55_15_i_5_n_0,
   I1 => W_55_15_i_14_n_0,
   I2 => x29_out_22,
   I3 => x29_out_29,
   I4 => x29_out_31,
   I5 => W_55_15_i_15_n_0,
   O => W_55_15_i_9_n_0
);
W_55_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x71_out_18,
   I1 => x44_out_18,
   I2 => x68_out_4,
   I3 => x68_out_25,
   I4 => x68_out_21,
   O => W_55_19_i_10_n_0
);
W_55_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x44_out_17,
   I1 => x68_out_20,
   I2 => x68_out_24,
   I3 => x68_out_3,
   I4 => x71_out_17,
   O => W_55_19_i_11_n_0
);
W_55_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x71_out_17,
   I1 => x44_out_17,
   I2 => x68_out_3,
   I3 => x68_out_24,
   I4 => x68_out_20,
   O => W_55_19_i_12_n_0
);
W_55_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x44_out_16,
   I1 => x68_out_19,
   I2 => x68_out_23,
   I3 => x68_out_2,
   I4 => x71_out_16,
   O => W_55_19_i_13_n_0
);
W_55_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x71_out_16,
   I1 => x44_out_16,
   I2 => x68_out_2,
   I3 => x68_out_23,
   I4 => x68_out_19,
   O => W_55_19_i_14_n_0
);
W_55_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x44_out_15,
   I1 => x68_out_18,
   I2 => x68_out_22,
   I3 => x68_out_1,
   I4 => x71_out_15,
   O => W_55_19_i_15_n_0
);
W_55_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x71_out_15,
   I1 => x44_out_15,
   I2 => x68_out_1,
   I3 => x68_out_22,
   I4 => x68_out_18,
   O => W_55_19_i_16_n_0
);
W_55_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x44_out_14,
   I1 => x68_out_17,
   I2 => x68_out_21,
   I3 => x68_out_0,
   I4 => x71_out_14,
   O => W_55_19_i_17_n_0
);
W_55_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x29_out_28,
   I1 => x29_out_3,
   I2 => x29_out_5,
   I3 => W_55_19_i_10_n_0,
   I4 => W_55_19_i_11_n_0,
   O => W_55_19_i_2_n_0
);
W_55_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x29_out_27,
   I1 => x29_out_2,
   I2 => x29_out_4,
   I3 => W_55_19_i_12_n_0,
   I4 => W_55_19_i_13_n_0,
   O => W_55_19_i_3_n_0
);
W_55_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x29_out_26,
   I1 => x29_out_1,
   I2 => x29_out_3,
   I3 => W_55_19_i_14_n_0,
   I4 => W_55_19_i_15_n_0,
   O => W_55_19_i_4_n_0
);
W_55_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x29_out_25,
   I1 => x29_out_0,
   I2 => x29_out_2,
   I3 => W_55_19_i_16_n_0,
   I4 => W_55_19_i_17_n_0,
   O => W_55_19_i_5_n_0
);
W_55_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_55_19_i_2_n_0,
   I1 => W_55_23_i_16_n_0,
   I2 => x29_out_29,
   I3 => x29_out_4,
   I4 => x29_out_6,
   I5 => W_55_23_i_17_n_0,
   O => W_55_19_i_6_n_0
);
W_55_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_55_19_i_3_n_0,
   I1 => W_55_19_i_10_n_0,
   I2 => x29_out_28,
   I3 => x29_out_3,
   I4 => x29_out_5,
   I5 => W_55_19_i_11_n_0,
   O => W_55_19_i_7_n_0
);
W_55_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_55_19_i_4_n_0,
   I1 => W_55_19_i_12_n_0,
   I2 => x29_out_27,
   I3 => x29_out_2,
   I4 => x29_out_4,
   I5 => W_55_19_i_13_n_0,
   O => W_55_19_i_8_n_0
);
W_55_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_55_19_i_5_n_0,
   I1 => W_55_19_i_14_n_0,
   I2 => x29_out_26,
   I3 => x29_out_1,
   I4 => x29_out_3,
   I5 => W_55_19_i_15_n_0,
   O => W_55_19_i_9_n_0
);
W_55_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x71_out_22,
   I1 => x44_out_22,
   I2 => x68_out_8,
   I3 => x68_out_29,
   I4 => x68_out_25,
   O => W_55_23_i_10_n_0
);
W_55_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x44_out_21,
   I1 => x68_out_24,
   I2 => x68_out_28,
   I3 => x68_out_7,
   I4 => x71_out_21,
   O => W_55_23_i_11_n_0
);
W_55_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x71_out_21,
   I1 => x44_out_21,
   I2 => x68_out_7,
   I3 => x68_out_28,
   I4 => x68_out_24,
   O => W_55_23_i_12_n_0
);
W_55_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x44_out_20,
   I1 => x68_out_23,
   I2 => x68_out_27,
   I3 => x68_out_6,
   I4 => x71_out_20,
   O => W_55_23_i_13_n_0
);
W_55_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x71_out_20,
   I1 => x44_out_20,
   I2 => x68_out_6,
   I3 => x68_out_27,
   I4 => x68_out_23,
   O => W_55_23_i_14_n_0
);
W_55_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x44_out_19,
   I1 => x68_out_22,
   I2 => x68_out_26,
   I3 => x68_out_5,
   I4 => x71_out_19,
   O => W_55_23_i_15_n_0
);
W_55_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x71_out_19,
   I1 => x44_out_19,
   I2 => x68_out_5,
   I3 => x68_out_26,
   I4 => x68_out_22,
   O => W_55_23_i_16_n_0
);
W_55_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x44_out_18,
   I1 => x68_out_21,
   I2 => x68_out_25,
   I3 => x68_out_4,
   I4 => x71_out_18,
   O => W_55_23_i_17_n_0
);
W_55_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x29_out_7,
   I1 => x29_out_9,
   I2 => W_55_23_i_10_n_0,
   I3 => W_55_23_i_11_n_0,
   O => W_55_23_i_2_n_0
);
W_55_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x29_out_31,
   I1 => x29_out_6,
   I2 => x29_out_8,
   I3 => W_55_23_i_12_n_0,
   I4 => W_55_23_i_13_n_0,
   O => W_55_23_i_3_n_0
);
W_55_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x29_out_30,
   I1 => x29_out_5,
   I2 => x29_out_7,
   I3 => W_55_23_i_14_n_0,
   I4 => W_55_23_i_15_n_0,
   O => W_55_23_i_4_n_0
);
W_55_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x29_out_29,
   I1 => x29_out_4,
   I2 => x29_out_6,
   I3 => W_55_23_i_16_n_0,
   I4 => W_55_23_i_17_n_0,
   O => W_55_23_i_5_n_0
);
W_55_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x29_out_8,
   I1 => x29_out_10,
   I2 => W_55_27_i_16_n_0,
   I3 => W_55_27_i_17_n_0,
   I4 => W_55_23_i_2_n_0,
   O => W_55_23_i_6_n_0
);
W_55_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x29_out_7,
   I1 => x29_out_9,
   I2 => W_55_23_i_10_n_0,
   I3 => W_55_23_i_11_n_0,
   I4 => W_55_23_i_3_n_0,
   O => W_55_23_i_7_n_0
);
W_55_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_55_23_i_4_n_0,
   I1 => W_55_23_i_12_n_0,
   I2 => x29_out_31,
   I3 => x29_out_6,
   I4 => x29_out_8,
   I5 => W_55_23_i_13_n_0,
   O => W_55_23_i_8_n_0
);
W_55_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_55_23_i_5_n_0,
   I1 => W_55_23_i_14_n_0,
   I2 => x29_out_30,
   I3 => x29_out_5,
   I4 => x29_out_7,
   I5 => W_55_23_i_15_n_0,
   O => W_55_23_i_9_n_0
);
W_55_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x71_out_26,
   I1 => x44_out_26,
   I2 => x68_out_12,
   I3 => x68_out_1,
   I4 => x68_out_29,
   O => W_55_27_i_10_n_0
);
W_55_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x44_out_25,
   I1 => x68_out_28,
   I2 => x68_out_0,
   I3 => x68_out_11,
   I4 => x71_out_25,
   O => W_55_27_i_11_n_0
);
W_55_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x71_out_25,
   I1 => x44_out_25,
   I2 => x68_out_11,
   I3 => x68_out_0,
   I4 => x68_out_28,
   O => W_55_27_i_12_n_0
);
W_55_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x44_out_24,
   I1 => x68_out_27,
   I2 => x68_out_31,
   I3 => x68_out_10,
   I4 => x71_out_24,
   O => W_55_27_i_13_n_0
);
W_55_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x71_out_24,
   I1 => x44_out_24,
   I2 => x68_out_10,
   I3 => x68_out_31,
   I4 => x68_out_27,
   O => W_55_27_i_14_n_0
);
W_55_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x44_out_23,
   I1 => x68_out_26,
   I2 => x68_out_30,
   I3 => x68_out_9,
   I4 => x71_out_23,
   O => W_55_27_i_15_n_0
);
W_55_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x71_out_23,
   I1 => x44_out_23,
   I2 => x68_out_9,
   I3 => x68_out_30,
   I4 => x68_out_26,
   O => W_55_27_i_16_n_0
);
W_55_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x44_out_22,
   I1 => x68_out_25,
   I2 => x68_out_29,
   I3 => x68_out_8,
   I4 => x71_out_22,
   O => W_55_27_i_17_n_0
);
W_55_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x29_out_11,
   I1 => x29_out_13,
   I2 => W_55_27_i_10_n_0,
   I3 => W_55_27_i_11_n_0,
   O => W_55_27_i_2_n_0
);
W_55_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x29_out_10,
   I1 => x29_out_12,
   I2 => W_55_27_i_12_n_0,
   I3 => W_55_27_i_13_n_0,
   O => W_55_27_i_3_n_0
);
W_55_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x29_out_9,
   I1 => x29_out_11,
   I2 => W_55_27_i_14_n_0,
   I3 => W_55_27_i_15_n_0,
   O => W_55_27_i_4_n_0
);
W_55_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x29_out_8,
   I1 => x29_out_10,
   I2 => W_55_27_i_16_n_0,
   I3 => W_55_27_i_17_n_0,
   O => W_55_27_i_5_n_0
);
W_55_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x29_out_12,
   I1 => x29_out_14,
   I2 => W_55_31_i_13_n_0,
   I3 => W_55_31_i_14_n_0,
   I4 => W_55_27_i_2_n_0,
   O => W_55_27_i_6_n_0
);
W_55_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x29_out_11,
   I1 => x29_out_13,
   I2 => W_55_27_i_10_n_0,
   I3 => W_55_27_i_11_n_0,
   I4 => W_55_27_i_3_n_0,
   O => W_55_27_i_7_n_0
);
W_55_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x29_out_10,
   I1 => x29_out_12,
   I2 => W_55_27_i_12_n_0,
   I3 => W_55_27_i_13_n_0,
   I4 => W_55_27_i_4_n_0,
   O => W_55_27_i_8_n_0
);
W_55_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x29_out_9,
   I1 => x29_out_11,
   I2 => W_55_27_i_14_n_0,
   I3 => W_55_27_i_15_n_0,
   I4 => W_55_27_i_5_n_0,
   O => W_55_27_i_9_n_0
);
W_55_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x44_out_28,
   I1 => x68_out_31,
   I2 => x68_out_3,
   I3 => x68_out_14,
   I4 => x71_out_28,
   O => W_55_31_i_10_n_0
);
W_55_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x71_out_28,
   I1 => x44_out_28,
   I2 => x68_out_14,
   I3 => x68_out_3,
   I4 => x68_out_31,
   O => W_55_31_i_11_n_0
);
W_55_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x44_out_27,
   I1 => x68_out_30,
   I2 => x68_out_2,
   I3 => x68_out_13,
   I4 => x71_out_27,
   O => W_55_31_i_12_n_0
);
W_55_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x71_out_27,
   I1 => x44_out_27,
   I2 => x68_out_13,
   I3 => x68_out_2,
   I4 => x68_out_30,
   O => W_55_31_i_13_n_0
);
W_55_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x44_out_26,
   I1 => x68_out_29,
   I2 => x68_out_1,
   I3 => x68_out_12,
   I4 => x71_out_26,
   O => W_55_31_i_14_n_0
);
W_55_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x44_out_29,
   I1 => x68_out_4,
   I2 => x68_out_15,
   I3 => x71_out_29,
   O => W_55_31_i_15_n_0
);
W_55_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x29_out_17,
   I1 => x29_out_15,
   O => SIGMA_LCASE_175_out_0_30
);
W_55_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => x68_out_6,
   I1 => x68_out_17,
   I2 => x44_out_31,
   I3 => x71_out_31,
   I4 => x29_out_16,
   I5 => x29_out_18,
   O => W_55_31_i_17_n_0
);
W_55_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x68_out_16,
   I1 => x68_out_5,
   O => SIGMA_LCASE_071_out_30
);
W_55_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x71_out_30,
   I1 => x44_out_30,
   I2 => x68_out_16,
   I3 => x68_out_5,
   O => W_55_31_i_19_n_0
);
W_55_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x29_out_14,
   I1 => x29_out_16,
   I2 => W_55_31_i_9_n_0,
   I3 => W_55_31_i_10_n_0,
   O => W_55_31_i_2_n_0
);
W_55_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x29_out_13,
   I1 => x29_out_15,
   I2 => W_55_31_i_11_n_0,
   I3 => W_55_31_i_12_n_0,
   O => W_55_31_i_3_n_0
);
W_55_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x29_out_12,
   I1 => x29_out_14,
   I2 => W_55_31_i_13_n_0,
   I3 => W_55_31_i_14_n_0,
   O => W_55_31_i_4_n_0
);
W_55_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_55_31_i_15_n_0,
   I1 => SIGMA_LCASE_175_out_0_30,
   I2 => W_55_31_i_17_n_0,
   I3 => x44_out_30,
   I4 => SIGMA_LCASE_071_out_30,
   I5 => x71_out_30,
   O => W_55_31_i_5_n_0
);
W_55_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_55_31_i_2_n_0,
   I1 => W_55_31_i_19_n_0,
   I2 => x29_out_15,
   I3 => x29_out_17,
   I4 => W_55_31_i_15_n_0,
   O => W_55_31_i_6_n_0
);
W_55_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x29_out_14,
   I1 => x29_out_16,
   I2 => W_55_31_i_9_n_0,
   I3 => W_55_31_i_10_n_0,
   I4 => W_55_31_i_3_n_0,
   O => W_55_31_i_7_n_0
);
W_55_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x29_out_13,
   I1 => x29_out_15,
   I2 => W_55_31_i_11_n_0,
   I3 => W_55_31_i_12_n_0,
   I4 => W_55_31_i_4_n_0,
   O => W_55_31_i_8_n_0
);
W_55_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x71_out_29,
   I1 => x44_out_29,
   I2 => x68_out_15,
   I3 => x68_out_4,
   O => W_55_31_i_9_n_0
);
W_55_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x71_out_2,
   I1 => x44_out_2,
   I2 => x68_out_20,
   I3 => x68_out_9,
   I4 => x68_out_5,
   O => W_55_3_i_10_n_0
);
W_55_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x44_out_1,
   I1 => x68_out_4,
   I2 => x68_out_8,
   I3 => x68_out_19,
   I4 => x71_out_1,
   O => W_55_3_i_11_n_0
);
W_55_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x68_out_19,
   I1 => x68_out_8,
   I2 => x68_out_4,
   O => SIGMA_LCASE_071_out_1
);
W_55_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x29_out_21,
   I1 => x29_out_19,
   I2 => x29_out_12,
   O => SIGMA_LCASE_175_out_0_2
);
W_55_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x29_out_20,
   I1 => x29_out_18,
   I2 => x29_out_11,
   O => SIGMA_LCASE_175_out_1
);
W_55_3_i_15 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x71_out_1,
   I1 => x44_out_1,
   I2 => x68_out_19,
   I3 => x68_out_8,
   I4 => x68_out_4,
   O => W_55_3_i_15_n_0
);
W_55_3_i_16 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x68_out_18,
   I1 => x68_out_7,
   I2 => x68_out_3,
   O => SIGMA_LCASE_071_out_0
);
W_55_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x29_out_12,
   I1 => x29_out_19,
   I2 => x29_out_21,
   I3 => W_55_3_i_10_n_0,
   I4 => W_55_3_i_11_n_0,
   O => W_55_3_i_2_n_0
);
W_55_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_55_3_i_11_n_0,
   I1 => x29_out_21,
   I2 => x29_out_19,
   I3 => x29_out_12,
   I4 => W_55_3_i_10_n_0,
   O => W_55_3_i_3_n_0
);
W_55_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_071_out_1,
   I1 => x44_out_1,
   I2 => x71_out_1,
   I3 => x29_out_11,
   I4 => x29_out_18,
   I5 => x29_out_20,
   O => W_55_3_i_4_n_0
);
W_55_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x71_out_0,
   I1 => x44_out_0,
   I2 => x68_out_18,
   I3 => x68_out_7,
   I4 => x68_out_3,
   O => W_55_3_i_5_n_0
);
W_55_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_55_3_i_2_n_0,
   I1 => W_55_7_i_16_n_0,
   I2 => x29_out_13,
   I3 => x29_out_20,
   I4 => x29_out_22,
   I5 => W_55_7_i_17_n_0,
   O => W_55_3_i_6_n_0
);
W_55_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_55_3_i_10_n_0,
   I1 => SIGMA_LCASE_175_out_0_2,
   I2 => x71_out_1,
   I3 => x44_out_1,
   I4 => SIGMA_LCASE_071_out_1,
   I5 => SIGMA_LCASE_175_out_1,
   O => W_55_3_i_7_n_0
);
W_55_3_i_8 : LUT5
  generic map(
   INIT => X"99969666"
  )
 port map (
   I0 => SIGMA_LCASE_175_out_1,
   I1 => W_55_3_i_15_n_0,
   I2 => x71_out_0,
   I3 => SIGMA_LCASE_071_out_0,
   I4 => x44_out_0,
   O => W_55_3_i_8_n_0
);
W_55_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_55_3_i_5_n_0,
   I1 => x29_out_10,
   I2 => x29_out_17,
   I3 => x29_out_19,
   O => W_55_3_i_9_n_0
);
W_55_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x71_out_6,
   I1 => x44_out_6,
   I2 => x68_out_24,
   I3 => x68_out_13,
   I4 => x68_out_9,
   O => W_55_7_i_10_n_0
);
W_55_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x44_out_5,
   I1 => x68_out_8,
   I2 => x68_out_12,
   I3 => x68_out_23,
   I4 => x71_out_5,
   O => W_55_7_i_11_n_0
);
W_55_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x71_out_5,
   I1 => x44_out_5,
   I2 => x68_out_23,
   I3 => x68_out_12,
   I4 => x68_out_8,
   O => W_55_7_i_12_n_0
);
W_55_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x44_out_4,
   I1 => x68_out_7,
   I2 => x68_out_11,
   I3 => x68_out_22,
   I4 => x71_out_4,
   O => W_55_7_i_13_n_0
);
W_55_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x71_out_4,
   I1 => x44_out_4,
   I2 => x68_out_22,
   I3 => x68_out_11,
   I4 => x68_out_7,
   O => W_55_7_i_14_n_0
);
W_55_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x44_out_3,
   I1 => x68_out_6,
   I2 => x68_out_10,
   I3 => x68_out_21,
   I4 => x71_out_3,
   O => W_55_7_i_15_n_0
);
W_55_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x71_out_3,
   I1 => x44_out_3,
   I2 => x68_out_21,
   I3 => x68_out_10,
   I4 => x68_out_6,
   O => W_55_7_i_16_n_0
);
W_55_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x44_out_2,
   I1 => x68_out_5,
   I2 => x68_out_9,
   I3 => x68_out_20,
   I4 => x71_out_2,
   O => W_55_7_i_17_n_0
);
W_55_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x29_out_16,
   I1 => x29_out_23,
   I2 => x29_out_25,
   I3 => W_55_7_i_10_n_0,
   I4 => W_55_7_i_11_n_0,
   O => W_55_7_i_2_n_0
);
W_55_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x29_out_15,
   I1 => x29_out_22,
   I2 => x29_out_24,
   I3 => W_55_7_i_12_n_0,
   I4 => W_55_7_i_13_n_0,
   O => W_55_7_i_3_n_0
);
W_55_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x29_out_14,
   I1 => x29_out_21,
   I2 => x29_out_23,
   I3 => W_55_7_i_14_n_0,
   I4 => W_55_7_i_15_n_0,
   O => W_55_7_i_4_n_0
);
W_55_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x29_out_13,
   I1 => x29_out_20,
   I2 => x29_out_22,
   I3 => W_55_7_i_16_n_0,
   I4 => W_55_7_i_17_n_0,
   O => W_55_7_i_5_n_0
);
W_55_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_55_7_i_2_n_0,
   I1 => W_55_11_i_16_n_0,
   I2 => x29_out_17,
   I3 => x29_out_24,
   I4 => x29_out_26,
   I5 => W_55_11_i_17_n_0,
   O => W_55_7_i_6_n_0
);
W_55_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_55_7_i_3_n_0,
   I1 => W_55_7_i_10_n_0,
   I2 => x29_out_16,
   I3 => x29_out_23,
   I4 => x29_out_25,
   I5 => W_55_7_i_11_n_0,
   O => W_55_7_i_7_n_0
);
W_55_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_55_7_i_4_n_0,
   I1 => W_55_7_i_12_n_0,
   I2 => x29_out_15,
   I3 => x29_out_22,
   I4 => x29_out_24,
   I5 => W_55_7_i_13_n_0,
   O => W_55_7_i_8_n_0
);
W_55_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_55_7_i_5_n_0,
   I1 => W_55_7_i_14_n_0,
   I2 => x29_out_14,
   I3 => x29_out_21,
   I4 => x29_out_23,
   I5 => W_55_7_i_15_n_0,
   O => W_55_7_i_9_n_0
);
W_56_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x68_out_10,
   I1 => x41_out_10,
   I2 => x65_out_28,
   I3 => x65_out_17,
   I4 => x65_out_13,
   O => W_56_11_i_10_n_0
);
W_56_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x41_out_9,
   I1 => x65_out_12,
   I2 => x65_out_16,
   I3 => x65_out_27,
   I4 => x68_out_9,
   O => W_56_11_i_11_n_0
);
W_56_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x68_out_9,
   I1 => x41_out_9,
   I2 => x65_out_27,
   I3 => x65_out_16,
   I4 => x65_out_12,
   O => W_56_11_i_12_n_0
);
W_56_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x41_out_8,
   I1 => x65_out_11,
   I2 => x65_out_15,
   I3 => x65_out_26,
   I4 => x68_out_8,
   O => W_56_11_i_13_n_0
);
W_56_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x68_out_8,
   I1 => x41_out_8,
   I2 => x65_out_26,
   I3 => x65_out_15,
   I4 => x65_out_11,
   O => W_56_11_i_14_n_0
);
W_56_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x41_out_7,
   I1 => x65_out_10,
   I2 => x65_out_14,
   I3 => x65_out_25,
   I4 => x68_out_7,
   O => W_56_11_i_15_n_0
);
W_56_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x68_out_7,
   I1 => x41_out_7,
   I2 => x65_out_25,
   I3 => x65_out_14,
   I4 => x65_out_10,
   O => W_56_11_i_16_n_0
);
W_56_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x41_out_6,
   I1 => x65_out_9,
   I2 => x65_out_13,
   I3 => x65_out_24,
   I4 => x68_out_6,
   O => W_56_11_i_17_n_0
);
W_56_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x26_out_20,
   I1 => x26_out_27,
   I2 => x26_out_29,
   I3 => W_56_11_i_10_n_0,
   I4 => W_56_11_i_11_n_0,
   O => W_56_11_i_2_n_0
);
W_56_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x26_out_19,
   I1 => x26_out_26,
   I2 => x26_out_28,
   I3 => W_56_11_i_12_n_0,
   I4 => W_56_11_i_13_n_0,
   O => W_56_11_i_3_n_0
);
W_56_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x26_out_18,
   I1 => x26_out_25,
   I2 => x26_out_27,
   I3 => W_56_11_i_14_n_0,
   I4 => W_56_11_i_15_n_0,
   O => W_56_11_i_4_n_0
);
W_56_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x26_out_17,
   I1 => x26_out_24,
   I2 => x26_out_26,
   I3 => W_56_11_i_16_n_0,
   I4 => W_56_11_i_17_n_0,
   O => W_56_11_i_5_n_0
);
W_56_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_56_11_i_2_n_0,
   I1 => W_56_15_i_16_n_0,
   I2 => x26_out_21,
   I3 => x26_out_28,
   I4 => x26_out_30,
   I5 => W_56_15_i_17_n_0,
   O => W_56_11_i_6_n_0
);
W_56_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_56_11_i_3_n_0,
   I1 => W_56_11_i_10_n_0,
   I2 => x26_out_20,
   I3 => x26_out_27,
   I4 => x26_out_29,
   I5 => W_56_11_i_11_n_0,
   O => W_56_11_i_7_n_0
);
W_56_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_56_11_i_4_n_0,
   I1 => W_56_11_i_12_n_0,
   I2 => x26_out_19,
   I3 => x26_out_26,
   I4 => x26_out_28,
   I5 => W_56_11_i_13_n_0,
   O => W_56_11_i_8_n_0
);
W_56_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_56_11_i_5_n_0,
   I1 => W_56_11_i_14_n_0,
   I2 => x26_out_18,
   I3 => x26_out_25,
   I4 => x26_out_27,
   I5 => W_56_11_i_15_n_0,
   O => W_56_11_i_9_n_0
);
W_56_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x68_out_14,
   I1 => x41_out_14,
   I2 => x65_out_0,
   I3 => x65_out_21,
   I4 => x65_out_17,
   O => W_56_15_i_10_n_0
);
W_56_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x41_out_13,
   I1 => x65_out_16,
   I2 => x65_out_20,
   I3 => x65_out_31,
   I4 => x68_out_13,
   O => W_56_15_i_11_n_0
);
W_56_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x68_out_13,
   I1 => x41_out_13,
   I2 => x65_out_31,
   I3 => x65_out_20,
   I4 => x65_out_16,
   O => W_56_15_i_12_n_0
);
W_56_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x41_out_12,
   I1 => x65_out_15,
   I2 => x65_out_19,
   I3 => x65_out_30,
   I4 => x68_out_12,
   O => W_56_15_i_13_n_0
);
W_56_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x68_out_12,
   I1 => x41_out_12,
   I2 => x65_out_30,
   I3 => x65_out_19,
   I4 => x65_out_15,
   O => W_56_15_i_14_n_0
);
W_56_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x41_out_11,
   I1 => x65_out_14,
   I2 => x65_out_18,
   I3 => x65_out_29,
   I4 => x68_out_11,
   O => W_56_15_i_15_n_0
);
W_56_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x68_out_11,
   I1 => x41_out_11,
   I2 => x65_out_29,
   I3 => x65_out_18,
   I4 => x65_out_14,
   O => W_56_15_i_16_n_0
);
W_56_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x41_out_10,
   I1 => x65_out_13,
   I2 => x65_out_17,
   I3 => x65_out_28,
   I4 => x68_out_10,
   O => W_56_15_i_17_n_0
);
W_56_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x26_out_24,
   I1 => x26_out_31,
   I2 => x26_out_1,
   I3 => W_56_15_i_10_n_0,
   I4 => W_56_15_i_11_n_0,
   O => W_56_15_i_2_n_0
);
W_56_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x26_out_23,
   I1 => x26_out_30,
   I2 => x26_out_0,
   I3 => W_56_15_i_12_n_0,
   I4 => W_56_15_i_13_n_0,
   O => W_56_15_i_3_n_0
);
W_56_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x26_out_22,
   I1 => x26_out_29,
   I2 => x26_out_31,
   I3 => W_56_15_i_14_n_0,
   I4 => W_56_15_i_15_n_0,
   O => W_56_15_i_4_n_0
);
W_56_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x26_out_21,
   I1 => x26_out_28,
   I2 => x26_out_30,
   I3 => W_56_15_i_16_n_0,
   I4 => W_56_15_i_17_n_0,
   O => W_56_15_i_5_n_0
);
W_56_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_56_15_i_2_n_0,
   I1 => W_56_19_i_16_n_0,
   I2 => x26_out_25,
   I3 => x26_out_0,
   I4 => x26_out_2,
   I5 => W_56_19_i_17_n_0,
   O => W_56_15_i_6_n_0
);
W_56_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_56_15_i_3_n_0,
   I1 => W_56_15_i_10_n_0,
   I2 => x26_out_24,
   I3 => x26_out_31,
   I4 => x26_out_1,
   I5 => W_56_15_i_11_n_0,
   O => W_56_15_i_7_n_0
);
W_56_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_56_15_i_4_n_0,
   I1 => W_56_15_i_12_n_0,
   I2 => x26_out_23,
   I3 => x26_out_30,
   I4 => x26_out_0,
   I5 => W_56_15_i_13_n_0,
   O => W_56_15_i_8_n_0
);
W_56_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_56_15_i_5_n_0,
   I1 => W_56_15_i_14_n_0,
   I2 => x26_out_22,
   I3 => x26_out_29,
   I4 => x26_out_31,
   I5 => W_56_15_i_15_n_0,
   O => W_56_15_i_9_n_0
);
W_56_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x68_out_18,
   I1 => x41_out_18,
   I2 => x65_out_4,
   I3 => x65_out_25,
   I4 => x65_out_21,
   O => W_56_19_i_10_n_0
);
W_56_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x41_out_17,
   I1 => x65_out_20,
   I2 => x65_out_24,
   I3 => x65_out_3,
   I4 => x68_out_17,
   O => W_56_19_i_11_n_0
);
W_56_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x68_out_17,
   I1 => x41_out_17,
   I2 => x65_out_3,
   I3 => x65_out_24,
   I4 => x65_out_20,
   O => W_56_19_i_12_n_0
);
W_56_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x41_out_16,
   I1 => x65_out_19,
   I2 => x65_out_23,
   I3 => x65_out_2,
   I4 => x68_out_16,
   O => W_56_19_i_13_n_0
);
W_56_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x68_out_16,
   I1 => x41_out_16,
   I2 => x65_out_2,
   I3 => x65_out_23,
   I4 => x65_out_19,
   O => W_56_19_i_14_n_0
);
W_56_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x41_out_15,
   I1 => x65_out_18,
   I2 => x65_out_22,
   I3 => x65_out_1,
   I4 => x68_out_15,
   O => W_56_19_i_15_n_0
);
W_56_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x68_out_15,
   I1 => x41_out_15,
   I2 => x65_out_1,
   I3 => x65_out_22,
   I4 => x65_out_18,
   O => W_56_19_i_16_n_0
);
W_56_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x41_out_14,
   I1 => x65_out_17,
   I2 => x65_out_21,
   I3 => x65_out_0,
   I4 => x68_out_14,
   O => W_56_19_i_17_n_0
);
W_56_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x26_out_28,
   I1 => x26_out_3,
   I2 => x26_out_5,
   I3 => W_56_19_i_10_n_0,
   I4 => W_56_19_i_11_n_0,
   O => W_56_19_i_2_n_0
);
W_56_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x26_out_27,
   I1 => x26_out_2,
   I2 => x26_out_4,
   I3 => W_56_19_i_12_n_0,
   I4 => W_56_19_i_13_n_0,
   O => W_56_19_i_3_n_0
);
W_56_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x26_out_26,
   I1 => x26_out_1,
   I2 => x26_out_3,
   I3 => W_56_19_i_14_n_0,
   I4 => W_56_19_i_15_n_0,
   O => W_56_19_i_4_n_0
);
W_56_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x26_out_25,
   I1 => x26_out_0,
   I2 => x26_out_2,
   I3 => W_56_19_i_16_n_0,
   I4 => W_56_19_i_17_n_0,
   O => W_56_19_i_5_n_0
);
W_56_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_56_19_i_2_n_0,
   I1 => W_56_23_i_16_n_0,
   I2 => x26_out_29,
   I3 => x26_out_4,
   I4 => x26_out_6,
   I5 => W_56_23_i_17_n_0,
   O => W_56_19_i_6_n_0
);
W_56_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_56_19_i_3_n_0,
   I1 => W_56_19_i_10_n_0,
   I2 => x26_out_28,
   I3 => x26_out_3,
   I4 => x26_out_5,
   I5 => W_56_19_i_11_n_0,
   O => W_56_19_i_7_n_0
);
W_56_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_56_19_i_4_n_0,
   I1 => W_56_19_i_12_n_0,
   I2 => x26_out_27,
   I3 => x26_out_2,
   I4 => x26_out_4,
   I5 => W_56_19_i_13_n_0,
   O => W_56_19_i_8_n_0
);
W_56_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_56_19_i_5_n_0,
   I1 => W_56_19_i_14_n_0,
   I2 => x26_out_26,
   I3 => x26_out_1,
   I4 => x26_out_3,
   I5 => W_56_19_i_15_n_0,
   O => W_56_19_i_9_n_0
);
W_56_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x68_out_22,
   I1 => x41_out_22,
   I2 => x65_out_8,
   I3 => x65_out_29,
   I4 => x65_out_25,
   O => W_56_23_i_10_n_0
);
W_56_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x41_out_21,
   I1 => x65_out_24,
   I2 => x65_out_28,
   I3 => x65_out_7,
   I4 => x68_out_21,
   O => W_56_23_i_11_n_0
);
W_56_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x68_out_21,
   I1 => x41_out_21,
   I2 => x65_out_7,
   I3 => x65_out_28,
   I4 => x65_out_24,
   O => W_56_23_i_12_n_0
);
W_56_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x41_out_20,
   I1 => x65_out_23,
   I2 => x65_out_27,
   I3 => x65_out_6,
   I4 => x68_out_20,
   O => W_56_23_i_13_n_0
);
W_56_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x68_out_20,
   I1 => x41_out_20,
   I2 => x65_out_6,
   I3 => x65_out_27,
   I4 => x65_out_23,
   O => W_56_23_i_14_n_0
);
W_56_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x41_out_19,
   I1 => x65_out_22,
   I2 => x65_out_26,
   I3 => x65_out_5,
   I4 => x68_out_19,
   O => W_56_23_i_15_n_0
);
W_56_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x68_out_19,
   I1 => x41_out_19,
   I2 => x65_out_5,
   I3 => x65_out_26,
   I4 => x65_out_22,
   O => W_56_23_i_16_n_0
);
W_56_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x41_out_18,
   I1 => x65_out_21,
   I2 => x65_out_25,
   I3 => x65_out_4,
   I4 => x68_out_18,
   O => W_56_23_i_17_n_0
);
W_56_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x26_out_7,
   I1 => x26_out_9,
   I2 => W_56_23_i_10_n_0,
   I3 => W_56_23_i_11_n_0,
   O => W_56_23_i_2_n_0
);
W_56_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x26_out_31,
   I1 => x26_out_6,
   I2 => x26_out_8,
   I3 => W_56_23_i_12_n_0,
   I4 => W_56_23_i_13_n_0,
   O => W_56_23_i_3_n_0
);
W_56_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x26_out_30,
   I1 => x26_out_5,
   I2 => x26_out_7,
   I3 => W_56_23_i_14_n_0,
   I4 => W_56_23_i_15_n_0,
   O => W_56_23_i_4_n_0
);
W_56_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x26_out_29,
   I1 => x26_out_4,
   I2 => x26_out_6,
   I3 => W_56_23_i_16_n_0,
   I4 => W_56_23_i_17_n_0,
   O => W_56_23_i_5_n_0
);
W_56_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x26_out_8,
   I1 => x26_out_10,
   I2 => W_56_27_i_16_n_0,
   I3 => W_56_27_i_17_n_0,
   I4 => W_56_23_i_2_n_0,
   O => W_56_23_i_6_n_0
);
W_56_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x26_out_7,
   I1 => x26_out_9,
   I2 => W_56_23_i_10_n_0,
   I3 => W_56_23_i_11_n_0,
   I4 => W_56_23_i_3_n_0,
   O => W_56_23_i_7_n_0
);
W_56_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_56_23_i_4_n_0,
   I1 => W_56_23_i_12_n_0,
   I2 => x26_out_31,
   I3 => x26_out_6,
   I4 => x26_out_8,
   I5 => W_56_23_i_13_n_0,
   O => W_56_23_i_8_n_0
);
W_56_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_56_23_i_5_n_0,
   I1 => W_56_23_i_14_n_0,
   I2 => x26_out_30,
   I3 => x26_out_5,
   I4 => x26_out_7,
   I5 => W_56_23_i_15_n_0,
   O => W_56_23_i_9_n_0
);
W_56_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x68_out_26,
   I1 => x41_out_26,
   I2 => x65_out_12,
   I3 => x65_out_1,
   I4 => x65_out_29,
   O => W_56_27_i_10_n_0
);
W_56_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x41_out_25,
   I1 => x65_out_28,
   I2 => x65_out_0,
   I3 => x65_out_11,
   I4 => x68_out_25,
   O => W_56_27_i_11_n_0
);
W_56_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x68_out_25,
   I1 => x41_out_25,
   I2 => x65_out_11,
   I3 => x65_out_0,
   I4 => x65_out_28,
   O => W_56_27_i_12_n_0
);
W_56_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x41_out_24,
   I1 => x65_out_27,
   I2 => x65_out_31,
   I3 => x65_out_10,
   I4 => x68_out_24,
   O => W_56_27_i_13_n_0
);
W_56_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x68_out_24,
   I1 => x41_out_24,
   I2 => x65_out_10,
   I3 => x65_out_31,
   I4 => x65_out_27,
   O => W_56_27_i_14_n_0
);
W_56_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x41_out_23,
   I1 => x65_out_26,
   I2 => x65_out_30,
   I3 => x65_out_9,
   I4 => x68_out_23,
   O => W_56_27_i_15_n_0
);
W_56_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x68_out_23,
   I1 => x41_out_23,
   I2 => x65_out_9,
   I3 => x65_out_30,
   I4 => x65_out_26,
   O => W_56_27_i_16_n_0
);
W_56_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x41_out_22,
   I1 => x65_out_25,
   I2 => x65_out_29,
   I3 => x65_out_8,
   I4 => x68_out_22,
   O => W_56_27_i_17_n_0
);
W_56_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x26_out_11,
   I1 => x26_out_13,
   I2 => W_56_27_i_10_n_0,
   I3 => W_56_27_i_11_n_0,
   O => W_56_27_i_2_n_0
);
W_56_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x26_out_10,
   I1 => x26_out_12,
   I2 => W_56_27_i_12_n_0,
   I3 => W_56_27_i_13_n_0,
   O => W_56_27_i_3_n_0
);
W_56_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x26_out_9,
   I1 => x26_out_11,
   I2 => W_56_27_i_14_n_0,
   I3 => W_56_27_i_15_n_0,
   O => W_56_27_i_4_n_0
);
W_56_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x26_out_8,
   I1 => x26_out_10,
   I2 => W_56_27_i_16_n_0,
   I3 => W_56_27_i_17_n_0,
   O => W_56_27_i_5_n_0
);
W_56_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x26_out_12,
   I1 => x26_out_14,
   I2 => W_56_31_i_13_n_0,
   I3 => W_56_31_i_14_n_0,
   I4 => W_56_27_i_2_n_0,
   O => W_56_27_i_6_n_0
);
W_56_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x26_out_11,
   I1 => x26_out_13,
   I2 => W_56_27_i_10_n_0,
   I3 => W_56_27_i_11_n_0,
   I4 => W_56_27_i_3_n_0,
   O => W_56_27_i_7_n_0
);
W_56_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x26_out_10,
   I1 => x26_out_12,
   I2 => W_56_27_i_12_n_0,
   I3 => W_56_27_i_13_n_0,
   I4 => W_56_27_i_4_n_0,
   O => W_56_27_i_8_n_0
);
W_56_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x26_out_9,
   I1 => x26_out_11,
   I2 => W_56_27_i_14_n_0,
   I3 => W_56_27_i_15_n_0,
   I4 => W_56_27_i_5_n_0,
   O => W_56_27_i_9_n_0
);
W_56_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x41_out_28,
   I1 => x65_out_31,
   I2 => x65_out_3,
   I3 => x65_out_14,
   I4 => x68_out_28,
   O => W_56_31_i_10_n_0
);
W_56_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x68_out_28,
   I1 => x41_out_28,
   I2 => x65_out_14,
   I3 => x65_out_3,
   I4 => x65_out_31,
   O => W_56_31_i_11_n_0
);
W_56_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x41_out_27,
   I1 => x65_out_30,
   I2 => x65_out_2,
   I3 => x65_out_13,
   I4 => x68_out_27,
   O => W_56_31_i_12_n_0
);
W_56_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x68_out_27,
   I1 => x41_out_27,
   I2 => x65_out_13,
   I3 => x65_out_2,
   I4 => x65_out_30,
   O => W_56_31_i_13_n_0
);
W_56_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x41_out_26,
   I1 => x65_out_29,
   I2 => x65_out_1,
   I3 => x65_out_12,
   I4 => x68_out_26,
   O => W_56_31_i_14_n_0
);
W_56_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x41_out_29,
   I1 => x65_out_4,
   I2 => x65_out_15,
   I3 => x68_out_29,
   O => W_56_31_i_15_n_0
);
W_56_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x26_out_17,
   I1 => x26_out_15,
   O => SIGMA_LCASE_167_out_0_30
);
W_56_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => x65_out_6,
   I1 => x65_out_17,
   I2 => x41_out_31,
   I3 => x68_out_31,
   I4 => x26_out_16,
   I5 => x26_out_18,
   O => W_56_31_i_17_n_0
);
W_56_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x65_out_16,
   I1 => x65_out_5,
   O => SIGMA_LCASE_063_out_30
);
W_56_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x68_out_30,
   I1 => x41_out_30,
   I2 => x65_out_16,
   I3 => x65_out_5,
   O => W_56_31_i_19_n_0
);
W_56_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x26_out_14,
   I1 => x26_out_16,
   I2 => W_56_31_i_9_n_0,
   I3 => W_56_31_i_10_n_0,
   O => W_56_31_i_2_n_0
);
W_56_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x26_out_13,
   I1 => x26_out_15,
   I2 => W_56_31_i_11_n_0,
   I3 => W_56_31_i_12_n_0,
   O => W_56_31_i_3_n_0
);
W_56_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x26_out_12,
   I1 => x26_out_14,
   I2 => W_56_31_i_13_n_0,
   I3 => W_56_31_i_14_n_0,
   O => W_56_31_i_4_n_0
);
W_56_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_56_31_i_15_n_0,
   I1 => SIGMA_LCASE_167_out_0_30,
   I2 => W_56_31_i_17_n_0,
   I3 => x41_out_30,
   I4 => SIGMA_LCASE_063_out_30,
   I5 => x68_out_30,
   O => W_56_31_i_5_n_0
);
W_56_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_56_31_i_2_n_0,
   I1 => W_56_31_i_19_n_0,
   I2 => x26_out_15,
   I3 => x26_out_17,
   I4 => W_56_31_i_15_n_0,
   O => W_56_31_i_6_n_0
);
W_56_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x26_out_14,
   I1 => x26_out_16,
   I2 => W_56_31_i_9_n_0,
   I3 => W_56_31_i_10_n_0,
   I4 => W_56_31_i_3_n_0,
   O => W_56_31_i_7_n_0
);
W_56_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x26_out_13,
   I1 => x26_out_15,
   I2 => W_56_31_i_11_n_0,
   I3 => W_56_31_i_12_n_0,
   I4 => W_56_31_i_4_n_0,
   O => W_56_31_i_8_n_0
);
W_56_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x68_out_29,
   I1 => x41_out_29,
   I2 => x65_out_15,
   I3 => x65_out_4,
   O => W_56_31_i_9_n_0
);
W_56_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x68_out_2,
   I1 => x41_out_2,
   I2 => x65_out_20,
   I3 => x65_out_9,
   I4 => x65_out_5,
   O => W_56_3_i_10_n_0
);
W_56_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x41_out_1,
   I1 => x65_out_4,
   I2 => x65_out_8,
   I3 => x65_out_19,
   I4 => x68_out_1,
   O => W_56_3_i_11_n_0
);
W_56_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x65_out_19,
   I1 => x65_out_8,
   I2 => x65_out_4,
   O => SIGMA_LCASE_063_out_1
);
W_56_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x26_out_21,
   I1 => x26_out_19,
   I2 => x26_out_12,
   O => SIGMA_LCASE_167_out_0_2
);
W_56_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x26_out_20,
   I1 => x26_out_18,
   I2 => x26_out_11,
   O => SIGMA_LCASE_167_out_1
);
W_56_3_i_15 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x68_out_1,
   I1 => x41_out_1,
   I2 => x65_out_19,
   I3 => x65_out_8,
   I4 => x65_out_4,
   O => W_56_3_i_15_n_0
);
W_56_3_i_16 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x65_out_18,
   I1 => x65_out_7,
   I2 => x65_out_3,
   O => SIGMA_LCASE_063_out_0
);
W_56_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x26_out_12,
   I1 => x26_out_19,
   I2 => x26_out_21,
   I3 => W_56_3_i_10_n_0,
   I4 => W_56_3_i_11_n_0,
   O => W_56_3_i_2_n_0
);
W_56_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_56_3_i_11_n_0,
   I1 => x26_out_21,
   I2 => x26_out_19,
   I3 => x26_out_12,
   I4 => W_56_3_i_10_n_0,
   O => W_56_3_i_3_n_0
);
W_56_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_063_out_1,
   I1 => x41_out_1,
   I2 => x68_out_1,
   I3 => x26_out_11,
   I4 => x26_out_18,
   I5 => x26_out_20,
   O => W_56_3_i_4_n_0
);
W_56_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x68_out_0,
   I1 => x41_out_0,
   I2 => x65_out_18,
   I3 => x65_out_7,
   I4 => x65_out_3,
   O => W_56_3_i_5_n_0
);
W_56_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_56_3_i_2_n_0,
   I1 => W_56_7_i_16_n_0,
   I2 => x26_out_13,
   I3 => x26_out_20,
   I4 => x26_out_22,
   I5 => W_56_7_i_17_n_0,
   O => W_56_3_i_6_n_0
);
W_56_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_56_3_i_10_n_0,
   I1 => SIGMA_LCASE_167_out_0_2,
   I2 => x68_out_1,
   I3 => x41_out_1,
   I4 => SIGMA_LCASE_063_out_1,
   I5 => SIGMA_LCASE_167_out_1,
   O => W_56_3_i_7_n_0
);
W_56_3_i_8 : LUT5
  generic map(
   INIT => X"99969666"
  )
 port map (
   I0 => SIGMA_LCASE_167_out_1,
   I1 => W_56_3_i_15_n_0,
   I2 => x68_out_0,
   I3 => SIGMA_LCASE_063_out_0,
   I4 => x41_out_0,
   O => W_56_3_i_8_n_0
);
W_56_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_56_3_i_5_n_0,
   I1 => x26_out_10,
   I2 => x26_out_17,
   I3 => x26_out_19,
   O => W_56_3_i_9_n_0
);
W_56_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x68_out_6,
   I1 => x41_out_6,
   I2 => x65_out_24,
   I3 => x65_out_13,
   I4 => x65_out_9,
   O => W_56_7_i_10_n_0
);
W_56_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x41_out_5,
   I1 => x65_out_8,
   I2 => x65_out_12,
   I3 => x65_out_23,
   I4 => x68_out_5,
   O => W_56_7_i_11_n_0
);
W_56_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x68_out_5,
   I1 => x41_out_5,
   I2 => x65_out_23,
   I3 => x65_out_12,
   I4 => x65_out_8,
   O => W_56_7_i_12_n_0
);
W_56_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x41_out_4,
   I1 => x65_out_7,
   I2 => x65_out_11,
   I3 => x65_out_22,
   I4 => x68_out_4,
   O => W_56_7_i_13_n_0
);
W_56_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x68_out_4,
   I1 => x41_out_4,
   I2 => x65_out_22,
   I3 => x65_out_11,
   I4 => x65_out_7,
   O => W_56_7_i_14_n_0
);
W_56_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x41_out_3,
   I1 => x65_out_6,
   I2 => x65_out_10,
   I3 => x65_out_21,
   I4 => x68_out_3,
   O => W_56_7_i_15_n_0
);
W_56_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x68_out_3,
   I1 => x41_out_3,
   I2 => x65_out_21,
   I3 => x65_out_10,
   I4 => x65_out_6,
   O => W_56_7_i_16_n_0
);
W_56_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x41_out_2,
   I1 => x65_out_5,
   I2 => x65_out_9,
   I3 => x65_out_20,
   I4 => x68_out_2,
   O => W_56_7_i_17_n_0
);
W_56_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x26_out_16,
   I1 => x26_out_23,
   I2 => x26_out_25,
   I3 => W_56_7_i_10_n_0,
   I4 => W_56_7_i_11_n_0,
   O => W_56_7_i_2_n_0
);
W_56_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x26_out_15,
   I1 => x26_out_22,
   I2 => x26_out_24,
   I3 => W_56_7_i_12_n_0,
   I4 => W_56_7_i_13_n_0,
   O => W_56_7_i_3_n_0
);
W_56_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x26_out_14,
   I1 => x26_out_21,
   I2 => x26_out_23,
   I3 => W_56_7_i_14_n_0,
   I4 => W_56_7_i_15_n_0,
   O => W_56_7_i_4_n_0
);
W_56_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x26_out_13,
   I1 => x26_out_20,
   I2 => x26_out_22,
   I3 => W_56_7_i_16_n_0,
   I4 => W_56_7_i_17_n_0,
   O => W_56_7_i_5_n_0
);
W_56_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_56_7_i_2_n_0,
   I1 => W_56_11_i_16_n_0,
   I2 => x26_out_17,
   I3 => x26_out_24,
   I4 => x26_out_26,
   I5 => W_56_11_i_17_n_0,
   O => W_56_7_i_6_n_0
);
W_56_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_56_7_i_3_n_0,
   I1 => W_56_7_i_10_n_0,
   I2 => x26_out_16,
   I3 => x26_out_23,
   I4 => x26_out_25,
   I5 => W_56_7_i_11_n_0,
   O => W_56_7_i_7_n_0
);
W_56_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_56_7_i_4_n_0,
   I1 => W_56_7_i_12_n_0,
   I2 => x26_out_15,
   I3 => x26_out_22,
   I4 => x26_out_24,
   I5 => W_56_7_i_13_n_0,
   O => W_56_7_i_8_n_0
);
W_56_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_56_7_i_5_n_0,
   I1 => W_56_7_i_14_n_0,
   I2 => x26_out_14,
   I3 => x26_out_21,
   I4 => x26_out_23,
   I5 => W_56_7_i_15_n_0,
   O => W_56_7_i_9_n_0
);
W_57_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x65_out_10,
   I1 => x38_out_10,
   I2 => x62_out_28,
   I3 => x62_out_17,
   I4 => x62_out_13,
   O => W_57_11_i_10_n_0
);
W_57_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x38_out_9,
   I1 => x62_out_12,
   I2 => x62_out_16,
   I3 => x62_out_27,
   I4 => x65_out_9,
   O => W_57_11_i_11_n_0
);
W_57_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x65_out_9,
   I1 => x38_out_9,
   I2 => x62_out_27,
   I3 => x62_out_16,
   I4 => x62_out_12,
   O => W_57_11_i_12_n_0
);
W_57_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x38_out_8,
   I1 => x62_out_11,
   I2 => x62_out_15,
   I3 => x62_out_26,
   I4 => x65_out_8,
   O => W_57_11_i_13_n_0
);
W_57_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x65_out_8,
   I1 => x38_out_8,
   I2 => x62_out_26,
   I3 => x62_out_15,
   I4 => x62_out_11,
   O => W_57_11_i_14_n_0
);
W_57_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x38_out_7,
   I1 => x62_out_10,
   I2 => x62_out_14,
   I3 => x62_out_25,
   I4 => x65_out_7,
   O => W_57_11_i_15_n_0
);
W_57_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x65_out_7,
   I1 => x38_out_7,
   I2 => x62_out_25,
   I3 => x62_out_14,
   I4 => x62_out_10,
   O => W_57_11_i_16_n_0
);
W_57_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x38_out_6,
   I1 => x62_out_9,
   I2 => x62_out_13,
   I3 => x62_out_24,
   I4 => x65_out_6,
   O => W_57_11_i_17_n_0
);
W_57_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x23_out_20,
   I1 => x23_out_27,
   I2 => x23_out_29,
   I3 => W_57_11_i_10_n_0,
   I4 => W_57_11_i_11_n_0,
   O => W_57_11_i_2_n_0
);
W_57_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x23_out_19,
   I1 => x23_out_26,
   I2 => x23_out_28,
   I3 => W_57_11_i_12_n_0,
   I4 => W_57_11_i_13_n_0,
   O => W_57_11_i_3_n_0
);
W_57_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x23_out_18,
   I1 => x23_out_25,
   I2 => x23_out_27,
   I3 => W_57_11_i_14_n_0,
   I4 => W_57_11_i_15_n_0,
   O => W_57_11_i_4_n_0
);
W_57_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x23_out_17,
   I1 => x23_out_24,
   I2 => x23_out_26,
   I3 => W_57_11_i_16_n_0,
   I4 => W_57_11_i_17_n_0,
   O => W_57_11_i_5_n_0
);
W_57_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_57_11_i_2_n_0,
   I1 => W_57_15_i_16_n_0,
   I2 => x23_out_21,
   I3 => x23_out_28,
   I4 => x23_out_30,
   I5 => W_57_15_i_17_n_0,
   O => W_57_11_i_6_n_0
);
W_57_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_57_11_i_3_n_0,
   I1 => W_57_11_i_10_n_0,
   I2 => x23_out_20,
   I3 => x23_out_27,
   I4 => x23_out_29,
   I5 => W_57_11_i_11_n_0,
   O => W_57_11_i_7_n_0
);
W_57_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_57_11_i_4_n_0,
   I1 => W_57_11_i_12_n_0,
   I2 => x23_out_19,
   I3 => x23_out_26,
   I4 => x23_out_28,
   I5 => W_57_11_i_13_n_0,
   O => W_57_11_i_8_n_0
);
W_57_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_57_11_i_5_n_0,
   I1 => W_57_11_i_14_n_0,
   I2 => x23_out_18,
   I3 => x23_out_25,
   I4 => x23_out_27,
   I5 => W_57_11_i_15_n_0,
   O => W_57_11_i_9_n_0
);
W_57_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x65_out_14,
   I1 => x38_out_14,
   I2 => x62_out_0,
   I3 => x62_out_21,
   I4 => x62_out_17,
   O => W_57_15_i_10_n_0
);
W_57_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x38_out_13,
   I1 => x62_out_16,
   I2 => x62_out_20,
   I3 => x62_out_31,
   I4 => x65_out_13,
   O => W_57_15_i_11_n_0
);
W_57_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x65_out_13,
   I1 => x38_out_13,
   I2 => x62_out_31,
   I3 => x62_out_20,
   I4 => x62_out_16,
   O => W_57_15_i_12_n_0
);
W_57_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x38_out_12,
   I1 => x62_out_15,
   I2 => x62_out_19,
   I3 => x62_out_30,
   I4 => x65_out_12,
   O => W_57_15_i_13_n_0
);
W_57_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x65_out_12,
   I1 => x38_out_12,
   I2 => x62_out_30,
   I3 => x62_out_19,
   I4 => x62_out_15,
   O => W_57_15_i_14_n_0
);
W_57_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x38_out_11,
   I1 => x62_out_14,
   I2 => x62_out_18,
   I3 => x62_out_29,
   I4 => x65_out_11,
   O => W_57_15_i_15_n_0
);
W_57_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x65_out_11,
   I1 => x38_out_11,
   I2 => x62_out_29,
   I3 => x62_out_18,
   I4 => x62_out_14,
   O => W_57_15_i_16_n_0
);
W_57_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x38_out_10,
   I1 => x62_out_13,
   I2 => x62_out_17,
   I3 => x62_out_28,
   I4 => x65_out_10,
   O => W_57_15_i_17_n_0
);
W_57_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x23_out_24,
   I1 => x23_out_31,
   I2 => x23_out_1,
   I3 => W_57_15_i_10_n_0,
   I4 => W_57_15_i_11_n_0,
   O => W_57_15_i_2_n_0
);
W_57_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x23_out_23,
   I1 => x23_out_30,
   I2 => x23_out_0,
   I3 => W_57_15_i_12_n_0,
   I4 => W_57_15_i_13_n_0,
   O => W_57_15_i_3_n_0
);
W_57_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x23_out_22,
   I1 => x23_out_29,
   I2 => x23_out_31,
   I3 => W_57_15_i_14_n_0,
   I4 => W_57_15_i_15_n_0,
   O => W_57_15_i_4_n_0
);
W_57_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x23_out_21,
   I1 => x23_out_28,
   I2 => x23_out_30,
   I3 => W_57_15_i_16_n_0,
   I4 => W_57_15_i_17_n_0,
   O => W_57_15_i_5_n_0
);
W_57_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_57_15_i_2_n_0,
   I1 => W_57_19_i_16_n_0,
   I2 => x23_out_25,
   I3 => x23_out_0,
   I4 => x23_out_2,
   I5 => W_57_19_i_17_n_0,
   O => W_57_15_i_6_n_0
);
W_57_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_57_15_i_3_n_0,
   I1 => W_57_15_i_10_n_0,
   I2 => x23_out_24,
   I3 => x23_out_31,
   I4 => x23_out_1,
   I5 => W_57_15_i_11_n_0,
   O => W_57_15_i_7_n_0
);
W_57_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_57_15_i_4_n_0,
   I1 => W_57_15_i_12_n_0,
   I2 => x23_out_23,
   I3 => x23_out_30,
   I4 => x23_out_0,
   I5 => W_57_15_i_13_n_0,
   O => W_57_15_i_8_n_0
);
W_57_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_57_15_i_5_n_0,
   I1 => W_57_15_i_14_n_0,
   I2 => x23_out_22,
   I3 => x23_out_29,
   I4 => x23_out_31,
   I5 => W_57_15_i_15_n_0,
   O => W_57_15_i_9_n_0
);
W_57_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x65_out_18,
   I1 => x38_out_18,
   I2 => x62_out_4,
   I3 => x62_out_25,
   I4 => x62_out_21,
   O => W_57_19_i_10_n_0
);
W_57_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x38_out_17,
   I1 => x62_out_20,
   I2 => x62_out_24,
   I3 => x62_out_3,
   I4 => x65_out_17,
   O => W_57_19_i_11_n_0
);
W_57_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x65_out_17,
   I1 => x38_out_17,
   I2 => x62_out_3,
   I3 => x62_out_24,
   I4 => x62_out_20,
   O => W_57_19_i_12_n_0
);
W_57_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x38_out_16,
   I1 => x62_out_19,
   I2 => x62_out_23,
   I3 => x62_out_2,
   I4 => x65_out_16,
   O => W_57_19_i_13_n_0
);
W_57_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x65_out_16,
   I1 => x38_out_16,
   I2 => x62_out_2,
   I3 => x62_out_23,
   I4 => x62_out_19,
   O => W_57_19_i_14_n_0
);
W_57_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x38_out_15,
   I1 => x62_out_18,
   I2 => x62_out_22,
   I3 => x62_out_1,
   I4 => x65_out_15,
   O => W_57_19_i_15_n_0
);
W_57_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x65_out_15,
   I1 => x38_out_15,
   I2 => x62_out_1,
   I3 => x62_out_22,
   I4 => x62_out_18,
   O => W_57_19_i_16_n_0
);
W_57_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x38_out_14,
   I1 => x62_out_17,
   I2 => x62_out_21,
   I3 => x62_out_0,
   I4 => x65_out_14,
   O => W_57_19_i_17_n_0
);
W_57_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x23_out_28,
   I1 => x23_out_3,
   I2 => x23_out_5,
   I3 => W_57_19_i_10_n_0,
   I4 => W_57_19_i_11_n_0,
   O => W_57_19_i_2_n_0
);
W_57_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x23_out_27,
   I1 => x23_out_2,
   I2 => x23_out_4,
   I3 => W_57_19_i_12_n_0,
   I4 => W_57_19_i_13_n_0,
   O => W_57_19_i_3_n_0
);
W_57_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x23_out_26,
   I1 => x23_out_1,
   I2 => x23_out_3,
   I3 => W_57_19_i_14_n_0,
   I4 => W_57_19_i_15_n_0,
   O => W_57_19_i_4_n_0
);
W_57_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x23_out_25,
   I1 => x23_out_0,
   I2 => x23_out_2,
   I3 => W_57_19_i_16_n_0,
   I4 => W_57_19_i_17_n_0,
   O => W_57_19_i_5_n_0
);
W_57_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_57_19_i_2_n_0,
   I1 => W_57_23_i_16_n_0,
   I2 => x23_out_29,
   I3 => x23_out_4,
   I4 => x23_out_6,
   I5 => W_57_23_i_17_n_0,
   O => W_57_19_i_6_n_0
);
W_57_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_57_19_i_3_n_0,
   I1 => W_57_19_i_10_n_0,
   I2 => x23_out_28,
   I3 => x23_out_3,
   I4 => x23_out_5,
   I5 => W_57_19_i_11_n_0,
   O => W_57_19_i_7_n_0
);
W_57_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_57_19_i_4_n_0,
   I1 => W_57_19_i_12_n_0,
   I2 => x23_out_27,
   I3 => x23_out_2,
   I4 => x23_out_4,
   I5 => W_57_19_i_13_n_0,
   O => W_57_19_i_8_n_0
);
W_57_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_57_19_i_5_n_0,
   I1 => W_57_19_i_14_n_0,
   I2 => x23_out_26,
   I3 => x23_out_1,
   I4 => x23_out_3,
   I5 => W_57_19_i_15_n_0,
   O => W_57_19_i_9_n_0
);
W_57_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x65_out_22,
   I1 => x38_out_22,
   I2 => x62_out_8,
   I3 => x62_out_29,
   I4 => x62_out_25,
   O => W_57_23_i_10_n_0
);
W_57_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x38_out_21,
   I1 => x62_out_24,
   I2 => x62_out_28,
   I3 => x62_out_7,
   I4 => x65_out_21,
   O => W_57_23_i_11_n_0
);
W_57_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x65_out_21,
   I1 => x38_out_21,
   I2 => x62_out_7,
   I3 => x62_out_28,
   I4 => x62_out_24,
   O => W_57_23_i_12_n_0
);
W_57_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x38_out_20,
   I1 => x62_out_23,
   I2 => x62_out_27,
   I3 => x62_out_6,
   I4 => x65_out_20,
   O => W_57_23_i_13_n_0
);
W_57_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x65_out_20,
   I1 => x38_out_20,
   I2 => x62_out_6,
   I3 => x62_out_27,
   I4 => x62_out_23,
   O => W_57_23_i_14_n_0
);
W_57_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x38_out_19,
   I1 => x62_out_22,
   I2 => x62_out_26,
   I3 => x62_out_5,
   I4 => x65_out_19,
   O => W_57_23_i_15_n_0
);
W_57_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x65_out_19,
   I1 => x38_out_19,
   I2 => x62_out_5,
   I3 => x62_out_26,
   I4 => x62_out_22,
   O => W_57_23_i_16_n_0
);
W_57_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x38_out_18,
   I1 => x62_out_21,
   I2 => x62_out_25,
   I3 => x62_out_4,
   I4 => x65_out_18,
   O => W_57_23_i_17_n_0
);
W_57_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x23_out_7,
   I1 => x23_out_9,
   I2 => W_57_23_i_10_n_0,
   I3 => W_57_23_i_11_n_0,
   O => W_57_23_i_2_n_0
);
W_57_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x23_out_31,
   I1 => x23_out_6,
   I2 => x23_out_8,
   I3 => W_57_23_i_12_n_0,
   I4 => W_57_23_i_13_n_0,
   O => W_57_23_i_3_n_0
);
W_57_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x23_out_30,
   I1 => x23_out_5,
   I2 => x23_out_7,
   I3 => W_57_23_i_14_n_0,
   I4 => W_57_23_i_15_n_0,
   O => W_57_23_i_4_n_0
);
W_57_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x23_out_29,
   I1 => x23_out_4,
   I2 => x23_out_6,
   I3 => W_57_23_i_16_n_0,
   I4 => W_57_23_i_17_n_0,
   O => W_57_23_i_5_n_0
);
W_57_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x23_out_8,
   I1 => x23_out_10,
   I2 => W_57_27_i_16_n_0,
   I3 => W_57_27_i_17_n_0,
   I4 => W_57_23_i_2_n_0,
   O => W_57_23_i_6_n_0
);
W_57_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x23_out_7,
   I1 => x23_out_9,
   I2 => W_57_23_i_10_n_0,
   I3 => W_57_23_i_11_n_0,
   I4 => W_57_23_i_3_n_0,
   O => W_57_23_i_7_n_0
);
W_57_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_57_23_i_4_n_0,
   I1 => W_57_23_i_12_n_0,
   I2 => x23_out_31,
   I3 => x23_out_6,
   I4 => x23_out_8,
   I5 => W_57_23_i_13_n_0,
   O => W_57_23_i_8_n_0
);
W_57_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_57_23_i_5_n_0,
   I1 => W_57_23_i_14_n_0,
   I2 => x23_out_30,
   I3 => x23_out_5,
   I4 => x23_out_7,
   I5 => W_57_23_i_15_n_0,
   O => W_57_23_i_9_n_0
);
W_57_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x65_out_26,
   I1 => x38_out_26,
   I2 => x62_out_12,
   I3 => x62_out_1,
   I4 => x62_out_29,
   O => W_57_27_i_10_n_0
);
W_57_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x38_out_25,
   I1 => x62_out_28,
   I2 => x62_out_0,
   I3 => x62_out_11,
   I4 => x65_out_25,
   O => W_57_27_i_11_n_0
);
W_57_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x65_out_25,
   I1 => x38_out_25,
   I2 => x62_out_11,
   I3 => x62_out_0,
   I4 => x62_out_28,
   O => W_57_27_i_12_n_0
);
W_57_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x38_out_24,
   I1 => x62_out_27,
   I2 => x62_out_31,
   I3 => x62_out_10,
   I4 => x65_out_24,
   O => W_57_27_i_13_n_0
);
W_57_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x65_out_24,
   I1 => x38_out_24,
   I2 => x62_out_10,
   I3 => x62_out_31,
   I4 => x62_out_27,
   O => W_57_27_i_14_n_0
);
W_57_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x38_out_23,
   I1 => x62_out_26,
   I2 => x62_out_30,
   I3 => x62_out_9,
   I4 => x65_out_23,
   O => W_57_27_i_15_n_0
);
W_57_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x65_out_23,
   I1 => x38_out_23,
   I2 => x62_out_9,
   I3 => x62_out_30,
   I4 => x62_out_26,
   O => W_57_27_i_16_n_0
);
W_57_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x38_out_22,
   I1 => x62_out_25,
   I2 => x62_out_29,
   I3 => x62_out_8,
   I4 => x65_out_22,
   O => W_57_27_i_17_n_0
);
W_57_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x23_out_11,
   I1 => x23_out_13,
   I2 => W_57_27_i_10_n_0,
   I3 => W_57_27_i_11_n_0,
   O => W_57_27_i_2_n_0
);
W_57_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x23_out_10,
   I1 => x23_out_12,
   I2 => W_57_27_i_12_n_0,
   I3 => W_57_27_i_13_n_0,
   O => W_57_27_i_3_n_0
);
W_57_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x23_out_9,
   I1 => x23_out_11,
   I2 => W_57_27_i_14_n_0,
   I3 => W_57_27_i_15_n_0,
   O => W_57_27_i_4_n_0
);
W_57_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x23_out_8,
   I1 => x23_out_10,
   I2 => W_57_27_i_16_n_0,
   I3 => W_57_27_i_17_n_0,
   O => W_57_27_i_5_n_0
);
W_57_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x23_out_12,
   I1 => x23_out_14,
   I2 => W_57_31_i_13_n_0,
   I3 => W_57_31_i_14_n_0,
   I4 => W_57_27_i_2_n_0,
   O => W_57_27_i_6_n_0
);
W_57_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x23_out_11,
   I1 => x23_out_13,
   I2 => W_57_27_i_10_n_0,
   I3 => W_57_27_i_11_n_0,
   I4 => W_57_27_i_3_n_0,
   O => W_57_27_i_7_n_0
);
W_57_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x23_out_10,
   I1 => x23_out_12,
   I2 => W_57_27_i_12_n_0,
   I3 => W_57_27_i_13_n_0,
   I4 => W_57_27_i_4_n_0,
   O => W_57_27_i_8_n_0
);
W_57_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x23_out_9,
   I1 => x23_out_11,
   I2 => W_57_27_i_14_n_0,
   I3 => W_57_27_i_15_n_0,
   I4 => W_57_27_i_5_n_0,
   O => W_57_27_i_9_n_0
);
W_57_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x38_out_28,
   I1 => x62_out_31,
   I2 => x62_out_3,
   I3 => x62_out_14,
   I4 => x65_out_28,
   O => W_57_31_i_10_n_0
);
W_57_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x65_out_28,
   I1 => x38_out_28,
   I2 => x62_out_14,
   I3 => x62_out_3,
   I4 => x62_out_31,
   O => W_57_31_i_11_n_0
);
W_57_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x38_out_27,
   I1 => x62_out_30,
   I2 => x62_out_2,
   I3 => x62_out_13,
   I4 => x65_out_27,
   O => W_57_31_i_12_n_0
);
W_57_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x65_out_27,
   I1 => x38_out_27,
   I2 => x62_out_13,
   I3 => x62_out_2,
   I4 => x62_out_30,
   O => W_57_31_i_13_n_0
);
W_57_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x38_out_26,
   I1 => x62_out_29,
   I2 => x62_out_1,
   I3 => x62_out_12,
   I4 => x65_out_26,
   O => W_57_31_i_14_n_0
);
W_57_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x38_out_29,
   I1 => x62_out_4,
   I2 => x62_out_15,
   I3 => x65_out_29,
   O => W_57_31_i_15_n_0
);
W_57_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x23_out_17,
   I1 => x23_out_15,
   O => SIGMA_LCASE_159_out_0_30
);
W_57_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => x62_out_6,
   I1 => x62_out_17,
   I2 => x38_out_31,
   I3 => x65_out_31,
   I4 => x23_out_16,
   I5 => x23_out_18,
   O => W_57_31_i_17_n_0
);
W_57_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x62_out_16,
   I1 => x62_out_5,
   O => SIGMA_LCASE_055_out_30
);
W_57_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x65_out_30,
   I1 => x38_out_30,
   I2 => x62_out_16,
   I3 => x62_out_5,
   O => W_57_31_i_19_n_0
);
W_57_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x23_out_14,
   I1 => x23_out_16,
   I2 => W_57_31_i_9_n_0,
   I3 => W_57_31_i_10_n_0,
   O => W_57_31_i_2_n_0
);
W_57_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x23_out_13,
   I1 => x23_out_15,
   I2 => W_57_31_i_11_n_0,
   I3 => W_57_31_i_12_n_0,
   O => W_57_31_i_3_n_0
);
W_57_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x23_out_12,
   I1 => x23_out_14,
   I2 => W_57_31_i_13_n_0,
   I3 => W_57_31_i_14_n_0,
   O => W_57_31_i_4_n_0
);
W_57_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_57_31_i_15_n_0,
   I1 => SIGMA_LCASE_159_out_0_30,
   I2 => W_57_31_i_17_n_0,
   I3 => x38_out_30,
   I4 => SIGMA_LCASE_055_out_30,
   I5 => x65_out_30,
   O => W_57_31_i_5_n_0
);
W_57_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_57_31_i_2_n_0,
   I1 => W_57_31_i_19_n_0,
   I2 => x23_out_15,
   I3 => x23_out_17,
   I4 => W_57_31_i_15_n_0,
   O => W_57_31_i_6_n_0
);
W_57_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x23_out_14,
   I1 => x23_out_16,
   I2 => W_57_31_i_9_n_0,
   I3 => W_57_31_i_10_n_0,
   I4 => W_57_31_i_3_n_0,
   O => W_57_31_i_7_n_0
);
W_57_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x23_out_13,
   I1 => x23_out_15,
   I2 => W_57_31_i_11_n_0,
   I3 => W_57_31_i_12_n_0,
   I4 => W_57_31_i_4_n_0,
   O => W_57_31_i_8_n_0
);
W_57_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x65_out_29,
   I1 => x38_out_29,
   I2 => x62_out_15,
   I3 => x62_out_4,
   O => W_57_31_i_9_n_0
);
W_57_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x65_out_2,
   I1 => x38_out_2,
   I2 => x62_out_20,
   I3 => x62_out_9,
   I4 => x62_out_5,
   O => W_57_3_i_10_n_0
);
W_57_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x38_out_1,
   I1 => x62_out_4,
   I2 => x62_out_8,
   I3 => x62_out_19,
   I4 => x65_out_1,
   O => W_57_3_i_11_n_0
);
W_57_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x62_out_19,
   I1 => x62_out_8,
   I2 => x62_out_4,
   O => SIGMA_LCASE_055_out_1
);
W_57_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x23_out_21,
   I1 => x23_out_19,
   I2 => x23_out_12,
   O => SIGMA_LCASE_159_out_0_2
);
W_57_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x23_out_20,
   I1 => x23_out_18,
   I2 => x23_out_11,
   O => SIGMA_LCASE_159_out_1
);
W_57_3_i_15 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x65_out_1,
   I1 => x38_out_1,
   I2 => x62_out_19,
   I3 => x62_out_8,
   I4 => x62_out_4,
   O => W_57_3_i_15_n_0
);
W_57_3_i_16 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x62_out_18,
   I1 => x62_out_7,
   I2 => x62_out_3,
   O => SIGMA_LCASE_055_out_0
);
W_57_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x23_out_12,
   I1 => x23_out_19,
   I2 => x23_out_21,
   I3 => W_57_3_i_10_n_0,
   I4 => W_57_3_i_11_n_0,
   O => W_57_3_i_2_n_0
);
W_57_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_57_3_i_11_n_0,
   I1 => x23_out_21,
   I2 => x23_out_19,
   I3 => x23_out_12,
   I4 => W_57_3_i_10_n_0,
   O => W_57_3_i_3_n_0
);
W_57_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_055_out_1,
   I1 => x38_out_1,
   I2 => x65_out_1,
   I3 => x23_out_11,
   I4 => x23_out_18,
   I5 => x23_out_20,
   O => W_57_3_i_4_n_0
);
W_57_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x65_out_0,
   I1 => x38_out_0,
   I2 => x62_out_18,
   I3 => x62_out_7,
   I4 => x62_out_3,
   O => W_57_3_i_5_n_0
);
W_57_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_57_3_i_2_n_0,
   I1 => W_57_7_i_16_n_0,
   I2 => x23_out_13,
   I3 => x23_out_20,
   I4 => x23_out_22,
   I5 => W_57_7_i_17_n_0,
   O => W_57_3_i_6_n_0
);
W_57_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_57_3_i_10_n_0,
   I1 => SIGMA_LCASE_159_out_0_2,
   I2 => x65_out_1,
   I3 => x38_out_1,
   I4 => SIGMA_LCASE_055_out_1,
   I5 => SIGMA_LCASE_159_out_1,
   O => W_57_3_i_7_n_0
);
W_57_3_i_8 : LUT5
  generic map(
   INIT => X"99969666"
  )
 port map (
   I0 => SIGMA_LCASE_159_out_1,
   I1 => W_57_3_i_15_n_0,
   I2 => x65_out_0,
   I3 => SIGMA_LCASE_055_out_0,
   I4 => x38_out_0,
   O => W_57_3_i_8_n_0
);
W_57_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_57_3_i_5_n_0,
   I1 => x23_out_10,
   I2 => x23_out_17,
   I3 => x23_out_19,
   O => W_57_3_i_9_n_0
);
W_57_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x65_out_6,
   I1 => x38_out_6,
   I2 => x62_out_24,
   I3 => x62_out_13,
   I4 => x62_out_9,
   O => W_57_7_i_10_n_0
);
W_57_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x38_out_5,
   I1 => x62_out_8,
   I2 => x62_out_12,
   I3 => x62_out_23,
   I4 => x65_out_5,
   O => W_57_7_i_11_n_0
);
W_57_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x65_out_5,
   I1 => x38_out_5,
   I2 => x62_out_23,
   I3 => x62_out_12,
   I4 => x62_out_8,
   O => W_57_7_i_12_n_0
);
W_57_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x38_out_4,
   I1 => x62_out_7,
   I2 => x62_out_11,
   I3 => x62_out_22,
   I4 => x65_out_4,
   O => W_57_7_i_13_n_0
);
W_57_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x65_out_4,
   I1 => x38_out_4,
   I2 => x62_out_22,
   I3 => x62_out_11,
   I4 => x62_out_7,
   O => W_57_7_i_14_n_0
);
W_57_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x38_out_3,
   I1 => x62_out_6,
   I2 => x62_out_10,
   I3 => x62_out_21,
   I4 => x65_out_3,
   O => W_57_7_i_15_n_0
);
W_57_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x65_out_3,
   I1 => x38_out_3,
   I2 => x62_out_21,
   I3 => x62_out_10,
   I4 => x62_out_6,
   O => W_57_7_i_16_n_0
);
W_57_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x38_out_2,
   I1 => x62_out_5,
   I2 => x62_out_9,
   I3 => x62_out_20,
   I4 => x65_out_2,
   O => W_57_7_i_17_n_0
);
W_57_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x23_out_16,
   I1 => x23_out_23,
   I2 => x23_out_25,
   I3 => W_57_7_i_10_n_0,
   I4 => W_57_7_i_11_n_0,
   O => W_57_7_i_2_n_0
);
W_57_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x23_out_15,
   I1 => x23_out_22,
   I2 => x23_out_24,
   I3 => W_57_7_i_12_n_0,
   I4 => W_57_7_i_13_n_0,
   O => W_57_7_i_3_n_0
);
W_57_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x23_out_14,
   I1 => x23_out_21,
   I2 => x23_out_23,
   I3 => W_57_7_i_14_n_0,
   I4 => W_57_7_i_15_n_0,
   O => W_57_7_i_4_n_0
);
W_57_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x23_out_13,
   I1 => x23_out_20,
   I2 => x23_out_22,
   I3 => W_57_7_i_16_n_0,
   I4 => W_57_7_i_17_n_0,
   O => W_57_7_i_5_n_0
);
W_57_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_57_7_i_2_n_0,
   I1 => W_57_11_i_16_n_0,
   I2 => x23_out_17,
   I3 => x23_out_24,
   I4 => x23_out_26,
   I5 => W_57_11_i_17_n_0,
   O => W_57_7_i_6_n_0
);
W_57_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_57_7_i_3_n_0,
   I1 => W_57_7_i_10_n_0,
   I2 => x23_out_16,
   I3 => x23_out_23,
   I4 => x23_out_25,
   I5 => W_57_7_i_11_n_0,
   O => W_57_7_i_7_n_0
);
W_57_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_57_7_i_4_n_0,
   I1 => W_57_7_i_12_n_0,
   I2 => x23_out_15,
   I3 => x23_out_22,
   I4 => x23_out_24,
   I5 => W_57_7_i_13_n_0,
   O => W_57_7_i_8_n_0
);
W_57_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_57_7_i_5_n_0,
   I1 => W_57_7_i_14_n_0,
   I2 => x23_out_14,
   I3 => x23_out_21,
   I4 => x23_out_23,
   I5 => W_57_7_i_15_n_0,
   O => W_57_7_i_9_n_0
);
W_58_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x62_out_10,
   I1 => x35_out_10,
   I2 => x59_out_28,
   I3 => x59_out_17,
   I4 => x59_out_13,
   O => W_58_11_i_10_n_0
);
W_58_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x35_out_9,
   I1 => x59_out_12,
   I2 => x59_out_16,
   I3 => x59_out_27,
   I4 => x62_out_9,
   O => W_58_11_i_11_n_0
);
W_58_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x62_out_9,
   I1 => x35_out_9,
   I2 => x59_out_27,
   I3 => x59_out_16,
   I4 => x59_out_12,
   O => W_58_11_i_12_n_0
);
W_58_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x35_out_8,
   I1 => x59_out_11,
   I2 => x59_out_15,
   I3 => x59_out_26,
   I4 => x62_out_8,
   O => W_58_11_i_13_n_0
);
W_58_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x62_out_8,
   I1 => x35_out_8,
   I2 => x59_out_26,
   I3 => x59_out_15,
   I4 => x59_out_11,
   O => W_58_11_i_14_n_0
);
W_58_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x35_out_7,
   I1 => x59_out_10,
   I2 => x59_out_14,
   I3 => x59_out_25,
   I4 => x62_out_7,
   O => W_58_11_i_15_n_0
);
W_58_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x62_out_7,
   I1 => x35_out_7,
   I2 => x59_out_25,
   I3 => x59_out_14,
   I4 => x59_out_10,
   O => W_58_11_i_16_n_0
);
W_58_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x35_out_6,
   I1 => x59_out_9,
   I2 => x59_out_13,
   I3 => x59_out_24,
   I4 => x62_out_6,
   O => W_58_11_i_17_n_0
);
W_58_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x20_out_20,
   I1 => x20_out_27,
   I2 => x20_out_29,
   I3 => W_58_11_i_10_n_0,
   I4 => W_58_11_i_11_n_0,
   O => W_58_11_i_2_n_0
);
W_58_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x20_out_19,
   I1 => x20_out_26,
   I2 => x20_out_28,
   I3 => W_58_11_i_12_n_0,
   I4 => W_58_11_i_13_n_0,
   O => W_58_11_i_3_n_0
);
W_58_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x20_out_18,
   I1 => x20_out_25,
   I2 => x20_out_27,
   I3 => W_58_11_i_14_n_0,
   I4 => W_58_11_i_15_n_0,
   O => W_58_11_i_4_n_0
);
W_58_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x20_out_17,
   I1 => x20_out_24,
   I2 => x20_out_26,
   I3 => W_58_11_i_16_n_0,
   I4 => W_58_11_i_17_n_0,
   O => W_58_11_i_5_n_0
);
W_58_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_58_11_i_2_n_0,
   I1 => W_58_15_i_16_n_0,
   I2 => x20_out_21,
   I3 => x20_out_28,
   I4 => x20_out_30,
   I5 => W_58_15_i_17_n_0,
   O => W_58_11_i_6_n_0
);
W_58_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_58_11_i_3_n_0,
   I1 => W_58_11_i_10_n_0,
   I2 => x20_out_20,
   I3 => x20_out_27,
   I4 => x20_out_29,
   I5 => W_58_11_i_11_n_0,
   O => W_58_11_i_7_n_0
);
W_58_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_58_11_i_4_n_0,
   I1 => W_58_11_i_12_n_0,
   I2 => x20_out_19,
   I3 => x20_out_26,
   I4 => x20_out_28,
   I5 => W_58_11_i_13_n_0,
   O => W_58_11_i_8_n_0
);
W_58_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_58_11_i_5_n_0,
   I1 => W_58_11_i_14_n_0,
   I2 => x20_out_18,
   I3 => x20_out_25,
   I4 => x20_out_27,
   I5 => W_58_11_i_15_n_0,
   O => W_58_11_i_9_n_0
);
W_58_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x62_out_14,
   I1 => x35_out_14,
   I2 => x59_out_0,
   I3 => x59_out_21,
   I4 => x59_out_17,
   O => W_58_15_i_10_n_0
);
W_58_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x35_out_13,
   I1 => x59_out_16,
   I2 => x59_out_20,
   I3 => x59_out_31,
   I4 => x62_out_13,
   O => W_58_15_i_11_n_0
);
W_58_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x62_out_13,
   I1 => x35_out_13,
   I2 => x59_out_31,
   I3 => x59_out_20,
   I4 => x59_out_16,
   O => W_58_15_i_12_n_0
);
W_58_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x35_out_12,
   I1 => x59_out_15,
   I2 => x59_out_19,
   I3 => x59_out_30,
   I4 => x62_out_12,
   O => W_58_15_i_13_n_0
);
W_58_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x62_out_12,
   I1 => x35_out_12,
   I2 => x59_out_30,
   I3 => x59_out_19,
   I4 => x59_out_15,
   O => W_58_15_i_14_n_0
);
W_58_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x35_out_11,
   I1 => x59_out_14,
   I2 => x59_out_18,
   I3 => x59_out_29,
   I4 => x62_out_11,
   O => W_58_15_i_15_n_0
);
W_58_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x62_out_11,
   I1 => x35_out_11,
   I2 => x59_out_29,
   I3 => x59_out_18,
   I4 => x59_out_14,
   O => W_58_15_i_16_n_0
);
W_58_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x35_out_10,
   I1 => x59_out_13,
   I2 => x59_out_17,
   I3 => x59_out_28,
   I4 => x62_out_10,
   O => W_58_15_i_17_n_0
);
W_58_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x20_out_24,
   I1 => x20_out_31,
   I2 => x20_out_1,
   I3 => W_58_15_i_10_n_0,
   I4 => W_58_15_i_11_n_0,
   O => W_58_15_i_2_n_0
);
W_58_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x20_out_23,
   I1 => x20_out_30,
   I2 => x20_out_0,
   I3 => W_58_15_i_12_n_0,
   I4 => W_58_15_i_13_n_0,
   O => W_58_15_i_3_n_0
);
W_58_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x20_out_22,
   I1 => x20_out_29,
   I2 => x20_out_31,
   I3 => W_58_15_i_14_n_0,
   I4 => W_58_15_i_15_n_0,
   O => W_58_15_i_4_n_0
);
W_58_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x20_out_21,
   I1 => x20_out_28,
   I2 => x20_out_30,
   I3 => W_58_15_i_16_n_0,
   I4 => W_58_15_i_17_n_0,
   O => W_58_15_i_5_n_0
);
W_58_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_58_15_i_2_n_0,
   I1 => W_58_19_i_16_n_0,
   I2 => x20_out_25,
   I3 => x20_out_0,
   I4 => x20_out_2,
   I5 => W_58_19_i_17_n_0,
   O => W_58_15_i_6_n_0
);
W_58_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_58_15_i_3_n_0,
   I1 => W_58_15_i_10_n_0,
   I2 => x20_out_24,
   I3 => x20_out_31,
   I4 => x20_out_1,
   I5 => W_58_15_i_11_n_0,
   O => W_58_15_i_7_n_0
);
W_58_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_58_15_i_4_n_0,
   I1 => W_58_15_i_12_n_0,
   I2 => x20_out_23,
   I3 => x20_out_30,
   I4 => x20_out_0,
   I5 => W_58_15_i_13_n_0,
   O => W_58_15_i_8_n_0
);
W_58_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_58_15_i_5_n_0,
   I1 => W_58_15_i_14_n_0,
   I2 => x20_out_22,
   I3 => x20_out_29,
   I4 => x20_out_31,
   I5 => W_58_15_i_15_n_0,
   O => W_58_15_i_9_n_0
);
W_58_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x62_out_18,
   I1 => x35_out_18,
   I2 => x59_out_4,
   I3 => x59_out_25,
   I4 => x59_out_21,
   O => W_58_19_i_10_n_0
);
W_58_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x35_out_17,
   I1 => x59_out_20,
   I2 => x59_out_24,
   I3 => x59_out_3,
   I4 => x62_out_17,
   O => W_58_19_i_11_n_0
);
W_58_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x62_out_17,
   I1 => x35_out_17,
   I2 => x59_out_3,
   I3 => x59_out_24,
   I4 => x59_out_20,
   O => W_58_19_i_12_n_0
);
W_58_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x35_out_16,
   I1 => x59_out_19,
   I2 => x59_out_23,
   I3 => x59_out_2,
   I4 => x62_out_16,
   O => W_58_19_i_13_n_0
);
W_58_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x62_out_16,
   I1 => x35_out_16,
   I2 => x59_out_2,
   I3 => x59_out_23,
   I4 => x59_out_19,
   O => W_58_19_i_14_n_0
);
W_58_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x35_out_15,
   I1 => x59_out_18,
   I2 => x59_out_22,
   I3 => x59_out_1,
   I4 => x62_out_15,
   O => W_58_19_i_15_n_0
);
W_58_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x62_out_15,
   I1 => x35_out_15,
   I2 => x59_out_1,
   I3 => x59_out_22,
   I4 => x59_out_18,
   O => W_58_19_i_16_n_0
);
W_58_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x35_out_14,
   I1 => x59_out_17,
   I2 => x59_out_21,
   I3 => x59_out_0,
   I4 => x62_out_14,
   O => W_58_19_i_17_n_0
);
W_58_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x20_out_28,
   I1 => x20_out_3,
   I2 => x20_out_5,
   I3 => W_58_19_i_10_n_0,
   I4 => W_58_19_i_11_n_0,
   O => W_58_19_i_2_n_0
);
W_58_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x20_out_27,
   I1 => x20_out_2,
   I2 => x20_out_4,
   I3 => W_58_19_i_12_n_0,
   I4 => W_58_19_i_13_n_0,
   O => W_58_19_i_3_n_0
);
W_58_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x20_out_26,
   I1 => x20_out_1,
   I2 => x20_out_3,
   I3 => W_58_19_i_14_n_0,
   I4 => W_58_19_i_15_n_0,
   O => W_58_19_i_4_n_0
);
W_58_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x20_out_25,
   I1 => x20_out_0,
   I2 => x20_out_2,
   I3 => W_58_19_i_16_n_0,
   I4 => W_58_19_i_17_n_0,
   O => W_58_19_i_5_n_0
);
W_58_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_58_19_i_2_n_0,
   I1 => W_58_23_i_16_n_0,
   I2 => x20_out_29,
   I3 => x20_out_4,
   I4 => x20_out_6,
   I5 => W_58_23_i_17_n_0,
   O => W_58_19_i_6_n_0
);
W_58_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_58_19_i_3_n_0,
   I1 => W_58_19_i_10_n_0,
   I2 => x20_out_28,
   I3 => x20_out_3,
   I4 => x20_out_5,
   I5 => W_58_19_i_11_n_0,
   O => W_58_19_i_7_n_0
);
W_58_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_58_19_i_4_n_0,
   I1 => W_58_19_i_12_n_0,
   I2 => x20_out_27,
   I3 => x20_out_2,
   I4 => x20_out_4,
   I5 => W_58_19_i_13_n_0,
   O => W_58_19_i_8_n_0
);
W_58_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_58_19_i_5_n_0,
   I1 => W_58_19_i_14_n_0,
   I2 => x20_out_26,
   I3 => x20_out_1,
   I4 => x20_out_3,
   I5 => W_58_19_i_15_n_0,
   O => W_58_19_i_9_n_0
);
W_58_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x62_out_22,
   I1 => x35_out_22,
   I2 => x59_out_8,
   I3 => x59_out_29,
   I4 => x59_out_25,
   O => W_58_23_i_10_n_0
);
W_58_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x35_out_21,
   I1 => x59_out_24,
   I2 => x59_out_28,
   I3 => x59_out_7,
   I4 => x62_out_21,
   O => W_58_23_i_11_n_0
);
W_58_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x62_out_21,
   I1 => x35_out_21,
   I2 => x59_out_7,
   I3 => x59_out_28,
   I4 => x59_out_24,
   O => W_58_23_i_12_n_0
);
W_58_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x35_out_20,
   I1 => x59_out_23,
   I2 => x59_out_27,
   I3 => x59_out_6,
   I4 => x62_out_20,
   O => W_58_23_i_13_n_0
);
W_58_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x62_out_20,
   I1 => x35_out_20,
   I2 => x59_out_6,
   I3 => x59_out_27,
   I4 => x59_out_23,
   O => W_58_23_i_14_n_0
);
W_58_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x35_out_19,
   I1 => x59_out_22,
   I2 => x59_out_26,
   I3 => x59_out_5,
   I4 => x62_out_19,
   O => W_58_23_i_15_n_0
);
W_58_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x62_out_19,
   I1 => x35_out_19,
   I2 => x59_out_5,
   I3 => x59_out_26,
   I4 => x59_out_22,
   O => W_58_23_i_16_n_0
);
W_58_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x35_out_18,
   I1 => x59_out_21,
   I2 => x59_out_25,
   I3 => x59_out_4,
   I4 => x62_out_18,
   O => W_58_23_i_17_n_0
);
W_58_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x20_out_7,
   I1 => x20_out_9,
   I2 => W_58_23_i_10_n_0,
   I3 => W_58_23_i_11_n_0,
   O => W_58_23_i_2_n_0
);
W_58_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x20_out_31,
   I1 => x20_out_6,
   I2 => x20_out_8,
   I3 => W_58_23_i_12_n_0,
   I4 => W_58_23_i_13_n_0,
   O => W_58_23_i_3_n_0
);
W_58_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x20_out_30,
   I1 => x20_out_5,
   I2 => x20_out_7,
   I3 => W_58_23_i_14_n_0,
   I4 => W_58_23_i_15_n_0,
   O => W_58_23_i_4_n_0
);
W_58_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x20_out_29,
   I1 => x20_out_4,
   I2 => x20_out_6,
   I3 => W_58_23_i_16_n_0,
   I4 => W_58_23_i_17_n_0,
   O => W_58_23_i_5_n_0
);
W_58_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x20_out_8,
   I1 => x20_out_10,
   I2 => W_58_27_i_16_n_0,
   I3 => W_58_27_i_17_n_0,
   I4 => W_58_23_i_2_n_0,
   O => W_58_23_i_6_n_0
);
W_58_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x20_out_7,
   I1 => x20_out_9,
   I2 => W_58_23_i_10_n_0,
   I3 => W_58_23_i_11_n_0,
   I4 => W_58_23_i_3_n_0,
   O => W_58_23_i_7_n_0
);
W_58_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_58_23_i_4_n_0,
   I1 => W_58_23_i_12_n_0,
   I2 => x20_out_31,
   I3 => x20_out_6,
   I4 => x20_out_8,
   I5 => W_58_23_i_13_n_0,
   O => W_58_23_i_8_n_0
);
W_58_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_58_23_i_5_n_0,
   I1 => W_58_23_i_14_n_0,
   I2 => x20_out_30,
   I3 => x20_out_5,
   I4 => x20_out_7,
   I5 => W_58_23_i_15_n_0,
   O => W_58_23_i_9_n_0
);
W_58_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x62_out_26,
   I1 => x35_out_26,
   I2 => x59_out_12,
   I3 => x59_out_1,
   I4 => x59_out_29,
   O => W_58_27_i_10_n_0
);
W_58_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x35_out_25,
   I1 => x59_out_28,
   I2 => x59_out_0,
   I3 => x59_out_11,
   I4 => x62_out_25,
   O => W_58_27_i_11_n_0
);
W_58_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x62_out_25,
   I1 => x35_out_25,
   I2 => x59_out_11,
   I3 => x59_out_0,
   I4 => x59_out_28,
   O => W_58_27_i_12_n_0
);
W_58_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x35_out_24,
   I1 => x59_out_27,
   I2 => x59_out_31,
   I3 => x59_out_10,
   I4 => x62_out_24,
   O => W_58_27_i_13_n_0
);
W_58_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x62_out_24,
   I1 => x35_out_24,
   I2 => x59_out_10,
   I3 => x59_out_31,
   I4 => x59_out_27,
   O => W_58_27_i_14_n_0
);
W_58_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x35_out_23,
   I1 => x59_out_26,
   I2 => x59_out_30,
   I3 => x59_out_9,
   I4 => x62_out_23,
   O => W_58_27_i_15_n_0
);
W_58_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x62_out_23,
   I1 => x35_out_23,
   I2 => x59_out_9,
   I3 => x59_out_30,
   I4 => x59_out_26,
   O => W_58_27_i_16_n_0
);
W_58_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x35_out_22,
   I1 => x59_out_25,
   I2 => x59_out_29,
   I3 => x59_out_8,
   I4 => x62_out_22,
   O => W_58_27_i_17_n_0
);
W_58_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x20_out_11,
   I1 => x20_out_13,
   I2 => W_58_27_i_10_n_0,
   I3 => W_58_27_i_11_n_0,
   O => W_58_27_i_2_n_0
);
W_58_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x20_out_10,
   I1 => x20_out_12,
   I2 => W_58_27_i_12_n_0,
   I3 => W_58_27_i_13_n_0,
   O => W_58_27_i_3_n_0
);
W_58_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x20_out_9,
   I1 => x20_out_11,
   I2 => W_58_27_i_14_n_0,
   I3 => W_58_27_i_15_n_0,
   O => W_58_27_i_4_n_0
);
W_58_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x20_out_8,
   I1 => x20_out_10,
   I2 => W_58_27_i_16_n_0,
   I3 => W_58_27_i_17_n_0,
   O => W_58_27_i_5_n_0
);
W_58_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x20_out_12,
   I1 => x20_out_14,
   I2 => W_58_31_i_13_n_0,
   I3 => W_58_31_i_14_n_0,
   I4 => W_58_27_i_2_n_0,
   O => W_58_27_i_6_n_0
);
W_58_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x20_out_11,
   I1 => x20_out_13,
   I2 => W_58_27_i_10_n_0,
   I3 => W_58_27_i_11_n_0,
   I4 => W_58_27_i_3_n_0,
   O => W_58_27_i_7_n_0
);
W_58_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x20_out_10,
   I1 => x20_out_12,
   I2 => W_58_27_i_12_n_0,
   I3 => W_58_27_i_13_n_0,
   I4 => W_58_27_i_4_n_0,
   O => W_58_27_i_8_n_0
);
W_58_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x20_out_9,
   I1 => x20_out_11,
   I2 => W_58_27_i_14_n_0,
   I3 => W_58_27_i_15_n_0,
   I4 => W_58_27_i_5_n_0,
   O => W_58_27_i_9_n_0
);
W_58_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x35_out_28,
   I1 => x59_out_31,
   I2 => x59_out_3,
   I3 => x59_out_14,
   I4 => x62_out_28,
   O => W_58_31_i_10_n_0
);
W_58_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x62_out_28,
   I1 => x35_out_28,
   I2 => x59_out_14,
   I3 => x59_out_3,
   I4 => x59_out_31,
   O => W_58_31_i_11_n_0
);
W_58_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x35_out_27,
   I1 => x59_out_30,
   I2 => x59_out_2,
   I3 => x59_out_13,
   I4 => x62_out_27,
   O => W_58_31_i_12_n_0
);
W_58_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x62_out_27,
   I1 => x35_out_27,
   I2 => x59_out_13,
   I3 => x59_out_2,
   I4 => x59_out_30,
   O => W_58_31_i_13_n_0
);
W_58_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x35_out_26,
   I1 => x59_out_29,
   I2 => x59_out_1,
   I3 => x59_out_12,
   I4 => x62_out_26,
   O => W_58_31_i_14_n_0
);
W_58_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x35_out_29,
   I1 => x59_out_4,
   I2 => x59_out_15,
   I3 => x62_out_29,
   O => W_58_31_i_15_n_0
);
W_58_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x20_out_17,
   I1 => x20_out_15,
   O => SIGMA_LCASE_151_out_0_30
);
W_58_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => x59_out_6,
   I1 => x59_out_17,
   I2 => x35_out_31,
   I3 => x62_out_31,
   I4 => x20_out_16,
   I5 => x20_out_18,
   O => W_58_31_i_17_n_0
);
W_58_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x59_out_16,
   I1 => x59_out_5,
   O => SIGMA_LCASE_047_out_30
);
W_58_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x62_out_30,
   I1 => x35_out_30,
   I2 => x59_out_16,
   I3 => x59_out_5,
   O => W_58_31_i_19_n_0
);
W_58_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x20_out_14,
   I1 => x20_out_16,
   I2 => W_58_31_i_9_n_0,
   I3 => W_58_31_i_10_n_0,
   O => W_58_31_i_2_n_0
);
W_58_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x20_out_13,
   I1 => x20_out_15,
   I2 => W_58_31_i_11_n_0,
   I3 => W_58_31_i_12_n_0,
   O => W_58_31_i_3_n_0
);
W_58_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x20_out_12,
   I1 => x20_out_14,
   I2 => W_58_31_i_13_n_0,
   I3 => W_58_31_i_14_n_0,
   O => W_58_31_i_4_n_0
);
W_58_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_58_31_i_15_n_0,
   I1 => SIGMA_LCASE_151_out_0_30,
   I2 => W_58_31_i_17_n_0,
   I3 => x35_out_30,
   I4 => SIGMA_LCASE_047_out_30,
   I5 => x62_out_30,
   O => W_58_31_i_5_n_0
);
W_58_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_58_31_i_2_n_0,
   I1 => W_58_31_i_19_n_0,
   I2 => x20_out_15,
   I3 => x20_out_17,
   I4 => W_58_31_i_15_n_0,
   O => W_58_31_i_6_n_0
);
W_58_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x20_out_14,
   I1 => x20_out_16,
   I2 => W_58_31_i_9_n_0,
   I3 => W_58_31_i_10_n_0,
   I4 => W_58_31_i_3_n_0,
   O => W_58_31_i_7_n_0
);
W_58_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x20_out_13,
   I1 => x20_out_15,
   I2 => W_58_31_i_11_n_0,
   I3 => W_58_31_i_12_n_0,
   I4 => W_58_31_i_4_n_0,
   O => W_58_31_i_8_n_0
);
W_58_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x62_out_29,
   I1 => x35_out_29,
   I2 => x59_out_15,
   I3 => x59_out_4,
   O => W_58_31_i_9_n_0
);
W_58_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x62_out_2,
   I1 => x35_out_2,
   I2 => x59_out_20,
   I3 => x59_out_9,
   I4 => x59_out_5,
   O => W_58_3_i_10_n_0
);
W_58_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x35_out_1,
   I1 => x59_out_4,
   I2 => x59_out_8,
   I3 => x59_out_19,
   I4 => x62_out_1,
   O => W_58_3_i_11_n_0
);
W_58_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x59_out_19,
   I1 => x59_out_8,
   I2 => x59_out_4,
   O => SIGMA_LCASE_047_out_1
);
W_58_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x20_out_21,
   I1 => x20_out_19,
   I2 => x20_out_12,
   O => SIGMA_LCASE_151_out_0_2
);
W_58_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x20_out_20,
   I1 => x20_out_18,
   I2 => x20_out_11,
   O => SIGMA_LCASE_151_out_1
);
W_58_3_i_15 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x62_out_1,
   I1 => x35_out_1,
   I2 => x59_out_19,
   I3 => x59_out_8,
   I4 => x59_out_4,
   O => W_58_3_i_15_n_0
);
W_58_3_i_16 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x59_out_18,
   I1 => x59_out_7,
   I2 => x59_out_3,
   O => SIGMA_LCASE_047_out_0
);
W_58_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x20_out_12,
   I1 => x20_out_19,
   I2 => x20_out_21,
   I3 => W_58_3_i_10_n_0,
   I4 => W_58_3_i_11_n_0,
   O => W_58_3_i_2_n_0
);
W_58_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_58_3_i_11_n_0,
   I1 => x20_out_21,
   I2 => x20_out_19,
   I3 => x20_out_12,
   I4 => W_58_3_i_10_n_0,
   O => W_58_3_i_3_n_0
);
W_58_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_047_out_1,
   I1 => x35_out_1,
   I2 => x62_out_1,
   I3 => x20_out_11,
   I4 => x20_out_18,
   I5 => x20_out_20,
   O => W_58_3_i_4_n_0
);
W_58_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x62_out_0,
   I1 => x35_out_0,
   I2 => x59_out_18,
   I3 => x59_out_7,
   I4 => x59_out_3,
   O => W_58_3_i_5_n_0
);
W_58_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_58_3_i_2_n_0,
   I1 => W_58_7_i_16_n_0,
   I2 => x20_out_13,
   I3 => x20_out_20,
   I4 => x20_out_22,
   I5 => W_58_7_i_17_n_0,
   O => W_58_3_i_6_n_0
);
W_58_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_58_3_i_10_n_0,
   I1 => SIGMA_LCASE_151_out_0_2,
   I2 => x62_out_1,
   I3 => x35_out_1,
   I4 => SIGMA_LCASE_047_out_1,
   I5 => SIGMA_LCASE_151_out_1,
   O => W_58_3_i_7_n_0
);
W_58_3_i_8 : LUT5
  generic map(
   INIT => X"99969666"
  )
 port map (
   I0 => SIGMA_LCASE_151_out_1,
   I1 => W_58_3_i_15_n_0,
   I2 => x62_out_0,
   I3 => SIGMA_LCASE_047_out_0,
   I4 => x35_out_0,
   O => W_58_3_i_8_n_0
);
W_58_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_58_3_i_5_n_0,
   I1 => x20_out_10,
   I2 => x20_out_17,
   I3 => x20_out_19,
   O => W_58_3_i_9_n_0
);
W_58_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x62_out_6,
   I1 => x35_out_6,
   I2 => x59_out_24,
   I3 => x59_out_13,
   I4 => x59_out_9,
   O => W_58_7_i_10_n_0
);
W_58_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x35_out_5,
   I1 => x59_out_8,
   I2 => x59_out_12,
   I3 => x59_out_23,
   I4 => x62_out_5,
   O => W_58_7_i_11_n_0
);
W_58_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x62_out_5,
   I1 => x35_out_5,
   I2 => x59_out_23,
   I3 => x59_out_12,
   I4 => x59_out_8,
   O => W_58_7_i_12_n_0
);
W_58_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x35_out_4,
   I1 => x59_out_7,
   I2 => x59_out_11,
   I3 => x59_out_22,
   I4 => x62_out_4,
   O => W_58_7_i_13_n_0
);
W_58_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x62_out_4,
   I1 => x35_out_4,
   I2 => x59_out_22,
   I3 => x59_out_11,
   I4 => x59_out_7,
   O => W_58_7_i_14_n_0
);
W_58_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x35_out_3,
   I1 => x59_out_6,
   I2 => x59_out_10,
   I3 => x59_out_21,
   I4 => x62_out_3,
   O => W_58_7_i_15_n_0
);
W_58_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x62_out_3,
   I1 => x35_out_3,
   I2 => x59_out_21,
   I3 => x59_out_10,
   I4 => x59_out_6,
   O => W_58_7_i_16_n_0
);
W_58_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x35_out_2,
   I1 => x59_out_5,
   I2 => x59_out_9,
   I3 => x59_out_20,
   I4 => x62_out_2,
   O => W_58_7_i_17_n_0
);
W_58_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x20_out_16,
   I1 => x20_out_23,
   I2 => x20_out_25,
   I3 => W_58_7_i_10_n_0,
   I4 => W_58_7_i_11_n_0,
   O => W_58_7_i_2_n_0
);
W_58_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x20_out_15,
   I1 => x20_out_22,
   I2 => x20_out_24,
   I3 => W_58_7_i_12_n_0,
   I4 => W_58_7_i_13_n_0,
   O => W_58_7_i_3_n_0
);
W_58_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x20_out_14,
   I1 => x20_out_21,
   I2 => x20_out_23,
   I3 => W_58_7_i_14_n_0,
   I4 => W_58_7_i_15_n_0,
   O => W_58_7_i_4_n_0
);
W_58_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x20_out_13,
   I1 => x20_out_20,
   I2 => x20_out_22,
   I3 => W_58_7_i_16_n_0,
   I4 => W_58_7_i_17_n_0,
   O => W_58_7_i_5_n_0
);
W_58_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_58_7_i_2_n_0,
   I1 => W_58_11_i_16_n_0,
   I2 => x20_out_17,
   I3 => x20_out_24,
   I4 => x20_out_26,
   I5 => W_58_11_i_17_n_0,
   O => W_58_7_i_6_n_0
);
W_58_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_58_7_i_3_n_0,
   I1 => W_58_7_i_10_n_0,
   I2 => x20_out_16,
   I3 => x20_out_23,
   I4 => x20_out_25,
   I5 => W_58_7_i_11_n_0,
   O => W_58_7_i_7_n_0
);
W_58_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_58_7_i_4_n_0,
   I1 => W_58_7_i_12_n_0,
   I2 => x20_out_15,
   I3 => x20_out_22,
   I4 => x20_out_24,
   I5 => W_58_7_i_13_n_0,
   O => W_58_7_i_8_n_0
);
W_58_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_58_7_i_5_n_0,
   I1 => W_58_7_i_14_n_0,
   I2 => x20_out_14,
   I3 => x20_out_21,
   I4 => x20_out_23,
   I5 => W_58_7_i_15_n_0,
   O => W_58_7_i_9_n_0
);
W_59_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x59_out_10,
   I1 => x32_out_10,
   I2 => x56_out_28,
   I3 => x56_out_17,
   I4 => x56_out_13,
   O => W_59_11_i_10_n_0
);
W_59_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x32_out_9,
   I1 => x56_out_12,
   I2 => x56_out_16,
   I3 => x56_out_27,
   I4 => x59_out_9,
   O => W_59_11_i_11_n_0
);
W_59_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x59_out_9,
   I1 => x32_out_9,
   I2 => x56_out_27,
   I3 => x56_out_16,
   I4 => x56_out_12,
   O => W_59_11_i_12_n_0
);
W_59_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x32_out_8,
   I1 => x56_out_11,
   I2 => x56_out_15,
   I3 => x56_out_26,
   I4 => x59_out_8,
   O => W_59_11_i_13_n_0
);
W_59_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x59_out_8,
   I1 => x32_out_8,
   I2 => x56_out_26,
   I3 => x56_out_15,
   I4 => x56_out_11,
   O => W_59_11_i_14_n_0
);
W_59_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x32_out_7,
   I1 => x56_out_10,
   I2 => x56_out_14,
   I3 => x56_out_25,
   I4 => x59_out_7,
   O => W_59_11_i_15_n_0
);
W_59_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x59_out_7,
   I1 => x32_out_7,
   I2 => x56_out_25,
   I3 => x56_out_14,
   I4 => x56_out_10,
   O => W_59_11_i_16_n_0
);
W_59_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x32_out_6,
   I1 => x56_out_9,
   I2 => x56_out_13,
   I3 => x56_out_24,
   I4 => x59_out_6,
   O => W_59_11_i_17_n_0
);
W_59_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x17_out_20,
   I1 => x17_out_27,
   I2 => x17_out_29,
   I3 => W_59_11_i_10_n_0,
   I4 => W_59_11_i_11_n_0,
   O => W_59_11_i_2_n_0
);
W_59_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x17_out_19,
   I1 => x17_out_26,
   I2 => x17_out_28,
   I3 => W_59_11_i_12_n_0,
   I4 => W_59_11_i_13_n_0,
   O => W_59_11_i_3_n_0
);
W_59_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x17_out_18,
   I1 => x17_out_25,
   I2 => x17_out_27,
   I3 => W_59_11_i_14_n_0,
   I4 => W_59_11_i_15_n_0,
   O => W_59_11_i_4_n_0
);
W_59_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x17_out_17,
   I1 => x17_out_24,
   I2 => x17_out_26,
   I3 => W_59_11_i_16_n_0,
   I4 => W_59_11_i_17_n_0,
   O => W_59_11_i_5_n_0
);
W_59_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_59_11_i_2_n_0,
   I1 => W_59_15_i_16_n_0,
   I2 => x17_out_21,
   I3 => x17_out_28,
   I4 => x17_out_30,
   I5 => W_59_15_i_17_n_0,
   O => W_59_11_i_6_n_0
);
W_59_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_59_11_i_3_n_0,
   I1 => W_59_11_i_10_n_0,
   I2 => x17_out_20,
   I3 => x17_out_27,
   I4 => x17_out_29,
   I5 => W_59_11_i_11_n_0,
   O => W_59_11_i_7_n_0
);
W_59_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_59_11_i_4_n_0,
   I1 => W_59_11_i_12_n_0,
   I2 => x17_out_19,
   I3 => x17_out_26,
   I4 => x17_out_28,
   I5 => W_59_11_i_13_n_0,
   O => W_59_11_i_8_n_0
);
W_59_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_59_11_i_5_n_0,
   I1 => W_59_11_i_14_n_0,
   I2 => x17_out_18,
   I3 => x17_out_25,
   I4 => x17_out_27,
   I5 => W_59_11_i_15_n_0,
   O => W_59_11_i_9_n_0
);
W_59_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x59_out_14,
   I1 => x32_out_14,
   I2 => x56_out_0,
   I3 => x56_out_21,
   I4 => x56_out_17,
   O => W_59_15_i_10_n_0
);
W_59_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x32_out_13,
   I1 => x56_out_16,
   I2 => x56_out_20,
   I3 => x56_out_31,
   I4 => x59_out_13,
   O => W_59_15_i_11_n_0
);
W_59_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x59_out_13,
   I1 => x32_out_13,
   I2 => x56_out_31,
   I3 => x56_out_20,
   I4 => x56_out_16,
   O => W_59_15_i_12_n_0
);
W_59_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x32_out_12,
   I1 => x56_out_15,
   I2 => x56_out_19,
   I3 => x56_out_30,
   I4 => x59_out_12,
   O => W_59_15_i_13_n_0
);
W_59_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x59_out_12,
   I1 => x32_out_12,
   I2 => x56_out_30,
   I3 => x56_out_19,
   I4 => x56_out_15,
   O => W_59_15_i_14_n_0
);
W_59_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x32_out_11,
   I1 => x56_out_14,
   I2 => x56_out_18,
   I3 => x56_out_29,
   I4 => x59_out_11,
   O => W_59_15_i_15_n_0
);
W_59_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x59_out_11,
   I1 => x32_out_11,
   I2 => x56_out_29,
   I3 => x56_out_18,
   I4 => x56_out_14,
   O => W_59_15_i_16_n_0
);
W_59_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x32_out_10,
   I1 => x56_out_13,
   I2 => x56_out_17,
   I3 => x56_out_28,
   I4 => x59_out_10,
   O => W_59_15_i_17_n_0
);
W_59_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x17_out_24,
   I1 => x17_out_31,
   I2 => x17_out_1,
   I3 => W_59_15_i_10_n_0,
   I4 => W_59_15_i_11_n_0,
   O => W_59_15_i_2_n_0
);
W_59_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x17_out_23,
   I1 => x17_out_30,
   I2 => x17_out_0,
   I3 => W_59_15_i_12_n_0,
   I4 => W_59_15_i_13_n_0,
   O => W_59_15_i_3_n_0
);
W_59_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x17_out_22,
   I1 => x17_out_29,
   I2 => x17_out_31,
   I3 => W_59_15_i_14_n_0,
   I4 => W_59_15_i_15_n_0,
   O => W_59_15_i_4_n_0
);
W_59_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x17_out_21,
   I1 => x17_out_28,
   I2 => x17_out_30,
   I3 => W_59_15_i_16_n_0,
   I4 => W_59_15_i_17_n_0,
   O => W_59_15_i_5_n_0
);
W_59_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_59_15_i_2_n_0,
   I1 => W_59_19_i_16_n_0,
   I2 => x17_out_25,
   I3 => x17_out_0,
   I4 => x17_out_2,
   I5 => W_59_19_i_17_n_0,
   O => W_59_15_i_6_n_0
);
W_59_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_59_15_i_3_n_0,
   I1 => W_59_15_i_10_n_0,
   I2 => x17_out_24,
   I3 => x17_out_31,
   I4 => x17_out_1,
   I5 => W_59_15_i_11_n_0,
   O => W_59_15_i_7_n_0
);
W_59_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_59_15_i_4_n_0,
   I1 => W_59_15_i_12_n_0,
   I2 => x17_out_23,
   I3 => x17_out_30,
   I4 => x17_out_0,
   I5 => W_59_15_i_13_n_0,
   O => W_59_15_i_8_n_0
);
W_59_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_59_15_i_5_n_0,
   I1 => W_59_15_i_14_n_0,
   I2 => x17_out_22,
   I3 => x17_out_29,
   I4 => x17_out_31,
   I5 => W_59_15_i_15_n_0,
   O => W_59_15_i_9_n_0
);
W_59_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x59_out_18,
   I1 => x32_out_18,
   I2 => x56_out_4,
   I3 => x56_out_25,
   I4 => x56_out_21,
   O => W_59_19_i_10_n_0
);
W_59_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x32_out_17,
   I1 => x56_out_20,
   I2 => x56_out_24,
   I3 => x56_out_3,
   I4 => x59_out_17,
   O => W_59_19_i_11_n_0
);
W_59_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x59_out_17,
   I1 => x32_out_17,
   I2 => x56_out_3,
   I3 => x56_out_24,
   I4 => x56_out_20,
   O => W_59_19_i_12_n_0
);
W_59_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x32_out_16,
   I1 => x56_out_19,
   I2 => x56_out_23,
   I3 => x56_out_2,
   I4 => x59_out_16,
   O => W_59_19_i_13_n_0
);
W_59_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x59_out_16,
   I1 => x32_out_16,
   I2 => x56_out_2,
   I3 => x56_out_23,
   I4 => x56_out_19,
   O => W_59_19_i_14_n_0
);
W_59_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x32_out_15,
   I1 => x56_out_18,
   I2 => x56_out_22,
   I3 => x56_out_1,
   I4 => x59_out_15,
   O => W_59_19_i_15_n_0
);
W_59_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x59_out_15,
   I1 => x32_out_15,
   I2 => x56_out_1,
   I3 => x56_out_22,
   I4 => x56_out_18,
   O => W_59_19_i_16_n_0
);
W_59_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x32_out_14,
   I1 => x56_out_17,
   I2 => x56_out_21,
   I3 => x56_out_0,
   I4 => x59_out_14,
   O => W_59_19_i_17_n_0
);
W_59_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x17_out_28,
   I1 => x17_out_3,
   I2 => x17_out_5,
   I3 => W_59_19_i_10_n_0,
   I4 => W_59_19_i_11_n_0,
   O => W_59_19_i_2_n_0
);
W_59_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x17_out_27,
   I1 => x17_out_2,
   I2 => x17_out_4,
   I3 => W_59_19_i_12_n_0,
   I4 => W_59_19_i_13_n_0,
   O => W_59_19_i_3_n_0
);
W_59_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x17_out_26,
   I1 => x17_out_1,
   I2 => x17_out_3,
   I3 => W_59_19_i_14_n_0,
   I4 => W_59_19_i_15_n_0,
   O => W_59_19_i_4_n_0
);
W_59_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x17_out_25,
   I1 => x17_out_0,
   I2 => x17_out_2,
   I3 => W_59_19_i_16_n_0,
   I4 => W_59_19_i_17_n_0,
   O => W_59_19_i_5_n_0
);
W_59_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_59_19_i_2_n_0,
   I1 => W_59_23_i_16_n_0,
   I2 => x17_out_29,
   I3 => x17_out_4,
   I4 => x17_out_6,
   I5 => W_59_23_i_17_n_0,
   O => W_59_19_i_6_n_0
);
W_59_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_59_19_i_3_n_0,
   I1 => W_59_19_i_10_n_0,
   I2 => x17_out_28,
   I3 => x17_out_3,
   I4 => x17_out_5,
   I5 => W_59_19_i_11_n_0,
   O => W_59_19_i_7_n_0
);
W_59_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_59_19_i_4_n_0,
   I1 => W_59_19_i_12_n_0,
   I2 => x17_out_27,
   I3 => x17_out_2,
   I4 => x17_out_4,
   I5 => W_59_19_i_13_n_0,
   O => W_59_19_i_8_n_0
);
W_59_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_59_19_i_5_n_0,
   I1 => W_59_19_i_14_n_0,
   I2 => x17_out_26,
   I3 => x17_out_1,
   I4 => x17_out_3,
   I5 => W_59_19_i_15_n_0,
   O => W_59_19_i_9_n_0
);
W_59_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x59_out_22,
   I1 => x32_out_22,
   I2 => x56_out_8,
   I3 => x56_out_29,
   I4 => x56_out_25,
   O => W_59_23_i_10_n_0
);
W_59_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x32_out_21,
   I1 => x56_out_24,
   I2 => x56_out_28,
   I3 => x56_out_7,
   I4 => x59_out_21,
   O => W_59_23_i_11_n_0
);
W_59_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x59_out_21,
   I1 => x32_out_21,
   I2 => x56_out_7,
   I3 => x56_out_28,
   I4 => x56_out_24,
   O => W_59_23_i_12_n_0
);
W_59_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x32_out_20,
   I1 => x56_out_23,
   I2 => x56_out_27,
   I3 => x56_out_6,
   I4 => x59_out_20,
   O => W_59_23_i_13_n_0
);
W_59_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x59_out_20,
   I1 => x32_out_20,
   I2 => x56_out_6,
   I3 => x56_out_27,
   I4 => x56_out_23,
   O => W_59_23_i_14_n_0
);
W_59_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x32_out_19,
   I1 => x56_out_22,
   I2 => x56_out_26,
   I3 => x56_out_5,
   I4 => x59_out_19,
   O => W_59_23_i_15_n_0
);
W_59_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x59_out_19,
   I1 => x32_out_19,
   I2 => x56_out_5,
   I3 => x56_out_26,
   I4 => x56_out_22,
   O => W_59_23_i_16_n_0
);
W_59_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x32_out_18,
   I1 => x56_out_21,
   I2 => x56_out_25,
   I3 => x56_out_4,
   I4 => x59_out_18,
   O => W_59_23_i_17_n_0
);
W_59_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x17_out_7,
   I1 => x17_out_9,
   I2 => W_59_23_i_10_n_0,
   I3 => W_59_23_i_11_n_0,
   O => W_59_23_i_2_n_0
);
W_59_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x17_out_31,
   I1 => x17_out_6,
   I2 => x17_out_8,
   I3 => W_59_23_i_12_n_0,
   I4 => W_59_23_i_13_n_0,
   O => W_59_23_i_3_n_0
);
W_59_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x17_out_30,
   I1 => x17_out_5,
   I2 => x17_out_7,
   I3 => W_59_23_i_14_n_0,
   I4 => W_59_23_i_15_n_0,
   O => W_59_23_i_4_n_0
);
W_59_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x17_out_29,
   I1 => x17_out_4,
   I2 => x17_out_6,
   I3 => W_59_23_i_16_n_0,
   I4 => W_59_23_i_17_n_0,
   O => W_59_23_i_5_n_0
);
W_59_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x17_out_8,
   I1 => x17_out_10,
   I2 => W_59_27_i_16_n_0,
   I3 => W_59_27_i_17_n_0,
   I4 => W_59_23_i_2_n_0,
   O => W_59_23_i_6_n_0
);
W_59_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x17_out_7,
   I1 => x17_out_9,
   I2 => W_59_23_i_10_n_0,
   I3 => W_59_23_i_11_n_0,
   I4 => W_59_23_i_3_n_0,
   O => W_59_23_i_7_n_0
);
W_59_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_59_23_i_4_n_0,
   I1 => W_59_23_i_12_n_0,
   I2 => x17_out_31,
   I3 => x17_out_6,
   I4 => x17_out_8,
   I5 => W_59_23_i_13_n_0,
   O => W_59_23_i_8_n_0
);
W_59_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_59_23_i_5_n_0,
   I1 => W_59_23_i_14_n_0,
   I2 => x17_out_30,
   I3 => x17_out_5,
   I4 => x17_out_7,
   I5 => W_59_23_i_15_n_0,
   O => W_59_23_i_9_n_0
);
W_59_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x59_out_26,
   I1 => x32_out_26,
   I2 => x56_out_12,
   I3 => x56_out_1,
   I4 => x56_out_29,
   O => W_59_27_i_10_n_0
);
W_59_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x32_out_25,
   I1 => x56_out_28,
   I2 => x56_out_0,
   I3 => x56_out_11,
   I4 => x59_out_25,
   O => W_59_27_i_11_n_0
);
W_59_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x59_out_25,
   I1 => x32_out_25,
   I2 => x56_out_11,
   I3 => x56_out_0,
   I4 => x56_out_28,
   O => W_59_27_i_12_n_0
);
W_59_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x32_out_24,
   I1 => x56_out_27,
   I2 => x56_out_31,
   I3 => x56_out_10,
   I4 => x59_out_24,
   O => W_59_27_i_13_n_0
);
W_59_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x59_out_24,
   I1 => x32_out_24,
   I2 => x56_out_10,
   I3 => x56_out_31,
   I4 => x56_out_27,
   O => W_59_27_i_14_n_0
);
W_59_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x32_out_23,
   I1 => x56_out_26,
   I2 => x56_out_30,
   I3 => x56_out_9,
   I4 => x59_out_23,
   O => W_59_27_i_15_n_0
);
W_59_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x59_out_23,
   I1 => x32_out_23,
   I2 => x56_out_9,
   I3 => x56_out_30,
   I4 => x56_out_26,
   O => W_59_27_i_16_n_0
);
W_59_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x32_out_22,
   I1 => x56_out_25,
   I2 => x56_out_29,
   I3 => x56_out_8,
   I4 => x59_out_22,
   O => W_59_27_i_17_n_0
);
W_59_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x17_out_11,
   I1 => x17_out_13,
   I2 => W_59_27_i_10_n_0,
   I3 => W_59_27_i_11_n_0,
   O => W_59_27_i_2_n_0
);
W_59_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x17_out_10,
   I1 => x17_out_12,
   I2 => W_59_27_i_12_n_0,
   I3 => W_59_27_i_13_n_0,
   O => W_59_27_i_3_n_0
);
W_59_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x17_out_9,
   I1 => x17_out_11,
   I2 => W_59_27_i_14_n_0,
   I3 => W_59_27_i_15_n_0,
   O => W_59_27_i_4_n_0
);
W_59_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x17_out_8,
   I1 => x17_out_10,
   I2 => W_59_27_i_16_n_0,
   I3 => W_59_27_i_17_n_0,
   O => W_59_27_i_5_n_0
);
W_59_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x17_out_12,
   I1 => x17_out_14,
   I2 => W_59_31_i_13_n_0,
   I3 => W_59_31_i_14_n_0,
   I4 => W_59_27_i_2_n_0,
   O => W_59_27_i_6_n_0
);
W_59_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x17_out_11,
   I1 => x17_out_13,
   I2 => W_59_27_i_10_n_0,
   I3 => W_59_27_i_11_n_0,
   I4 => W_59_27_i_3_n_0,
   O => W_59_27_i_7_n_0
);
W_59_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x17_out_10,
   I1 => x17_out_12,
   I2 => W_59_27_i_12_n_0,
   I3 => W_59_27_i_13_n_0,
   I4 => W_59_27_i_4_n_0,
   O => W_59_27_i_8_n_0
);
W_59_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x17_out_9,
   I1 => x17_out_11,
   I2 => W_59_27_i_14_n_0,
   I3 => W_59_27_i_15_n_0,
   I4 => W_59_27_i_5_n_0,
   O => W_59_27_i_9_n_0
);
W_59_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x32_out_28,
   I1 => x56_out_31,
   I2 => x56_out_3,
   I3 => x56_out_14,
   I4 => x59_out_28,
   O => W_59_31_i_10_n_0
);
W_59_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x59_out_28,
   I1 => x32_out_28,
   I2 => x56_out_14,
   I3 => x56_out_3,
   I4 => x56_out_31,
   O => W_59_31_i_11_n_0
);
W_59_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x32_out_27,
   I1 => x56_out_30,
   I2 => x56_out_2,
   I3 => x56_out_13,
   I4 => x59_out_27,
   O => W_59_31_i_12_n_0
);
W_59_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x59_out_27,
   I1 => x32_out_27,
   I2 => x56_out_13,
   I3 => x56_out_2,
   I4 => x56_out_30,
   O => W_59_31_i_13_n_0
);
W_59_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x32_out_26,
   I1 => x56_out_29,
   I2 => x56_out_1,
   I3 => x56_out_12,
   I4 => x59_out_26,
   O => W_59_31_i_14_n_0
);
W_59_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x32_out_29,
   I1 => x56_out_4,
   I2 => x56_out_15,
   I3 => x59_out_29,
   O => W_59_31_i_15_n_0
);
W_59_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x17_out_17,
   I1 => x17_out_15,
   O => SIGMA_LCASE_143_out_0_30
);
W_59_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => x56_out_6,
   I1 => x56_out_17,
   I2 => x32_out_31,
   I3 => x59_out_31,
   I4 => x17_out_16,
   I5 => x17_out_18,
   O => W_59_31_i_17_n_0
);
W_59_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x56_out_16,
   I1 => x56_out_5,
   O => SIGMA_LCASE_039_out_30
);
W_59_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x59_out_30,
   I1 => x32_out_30,
   I2 => x56_out_16,
   I3 => x56_out_5,
   O => W_59_31_i_19_n_0
);
W_59_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x17_out_14,
   I1 => x17_out_16,
   I2 => W_59_31_i_9_n_0,
   I3 => W_59_31_i_10_n_0,
   O => W_59_31_i_2_n_0
);
W_59_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x17_out_13,
   I1 => x17_out_15,
   I2 => W_59_31_i_11_n_0,
   I3 => W_59_31_i_12_n_0,
   O => W_59_31_i_3_n_0
);
W_59_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x17_out_12,
   I1 => x17_out_14,
   I2 => W_59_31_i_13_n_0,
   I3 => W_59_31_i_14_n_0,
   O => W_59_31_i_4_n_0
);
W_59_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_59_31_i_15_n_0,
   I1 => SIGMA_LCASE_143_out_0_30,
   I2 => W_59_31_i_17_n_0,
   I3 => x32_out_30,
   I4 => SIGMA_LCASE_039_out_30,
   I5 => x59_out_30,
   O => W_59_31_i_5_n_0
);
W_59_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_59_31_i_2_n_0,
   I1 => W_59_31_i_19_n_0,
   I2 => x17_out_15,
   I3 => x17_out_17,
   I4 => W_59_31_i_15_n_0,
   O => W_59_31_i_6_n_0
);
W_59_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x17_out_14,
   I1 => x17_out_16,
   I2 => W_59_31_i_9_n_0,
   I3 => W_59_31_i_10_n_0,
   I4 => W_59_31_i_3_n_0,
   O => W_59_31_i_7_n_0
);
W_59_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x17_out_13,
   I1 => x17_out_15,
   I2 => W_59_31_i_11_n_0,
   I3 => W_59_31_i_12_n_0,
   I4 => W_59_31_i_4_n_0,
   O => W_59_31_i_8_n_0
);
W_59_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x59_out_29,
   I1 => x32_out_29,
   I2 => x56_out_15,
   I3 => x56_out_4,
   O => W_59_31_i_9_n_0
);
W_59_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x59_out_2,
   I1 => x32_out_2,
   I2 => x56_out_20,
   I3 => x56_out_9,
   I4 => x56_out_5,
   O => W_59_3_i_10_n_0
);
W_59_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x32_out_1,
   I1 => x56_out_4,
   I2 => x56_out_8,
   I3 => x56_out_19,
   I4 => x59_out_1,
   O => W_59_3_i_11_n_0
);
W_59_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x56_out_19,
   I1 => x56_out_8,
   I2 => x56_out_4,
   O => SIGMA_LCASE_039_out_1
);
W_59_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x17_out_21,
   I1 => x17_out_19,
   I2 => x17_out_12,
   O => SIGMA_LCASE_143_out_0_2
);
W_59_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x17_out_20,
   I1 => x17_out_18,
   I2 => x17_out_11,
   O => SIGMA_LCASE_143_out_1
);
W_59_3_i_15 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x59_out_1,
   I1 => x32_out_1,
   I2 => x56_out_19,
   I3 => x56_out_8,
   I4 => x56_out_4,
   O => W_59_3_i_15_n_0
);
W_59_3_i_16 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x56_out_18,
   I1 => x56_out_7,
   I2 => x56_out_3,
   O => SIGMA_LCASE_039_out_0
);
W_59_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x17_out_12,
   I1 => x17_out_19,
   I2 => x17_out_21,
   I3 => W_59_3_i_10_n_0,
   I4 => W_59_3_i_11_n_0,
   O => W_59_3_i_2_n_0
);
W_59_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_59_3_i_11_n_0,
   I1 => x17_out_21,
   I2 => x17_out_19,
   I3 => x17_out_12,
   I4 => W_59_3_i_10_n_0,
   O => W_59_3_i_3_n_0
);
W_59_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_039_out_1,
   I1 => x32_out_1,
   I2 => x59_out_1,
   I3 => x17_out_11,
   I4 => x17_out_18,
   I5 => x17_out_20,
   O => W_59_3_i_4_n_0
);
W_59_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x59_out_0,
   I1 => x32_out_0,
   I2 => x56_out_18,
   I3 => x56_out_7,
   I4 => x56_out_3,
   O => W_59_3_i_5_n_0
);
W_59_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_59_3_i_2_n_0,
   I1 => W_59_7_i_16_n_0,
   I2 => x17_out_13,
   I3 => x17_out_20,
   I4 => x17_out_22,
   I5 => W_59_7_i_17_n_0,
   O => W_59_3_i_6_n_0
);
W_59_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_59_3_i_10_n_0,
   I1 => SIGMA_LCASE_143_out_0_2,
   I2 => x59_out_1,
   I3 => x32_out_1,
   I4 => SIGMA_LCASE_039_out_1,
   I5 => SIGMA_LCASE_143_out_1,
   O => W_59_3_i_7_n_0
);
W_59_3_i_8 : LUT5
  generic map(
   INIT => X"99969666"
  )
 port map (
   I0 => SIGMA_LCASE_143_out_1,
   I1 => W_59_3_i_15_n_0,
   I2 => x59_out_0,
   I3 => SIGMA_LCASE_039_out_0,
   I4 => x32_out_0,
   O => W_59_3_i_8_n_0
);
W_59_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_59_3_i_5_n_0,
   I1 => x17_out_10,
   I2 => x17_out_17,
   I3 => x17_out_19,
   O => W_59_3_i_9_n_0
);
W_59_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x59_out_6,
   I1 => x32_out_6,
   I2 => x56_out_24,
   I3 => x56_out_13,
   I4 => x56_out_9,
   O => W_59_7_i_10_n_0
);
W_59_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x32_out_5,
   I1 => x56_out_8,
   I2 => x56_out_12,
   I3 => x56_out_23,
   I4 => x59_out_5,
   O => W_59_7_i_11_n_0
);
W_59_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x59_out_5,
   I1 => x32_out_5,
   I2 => x56_out_23,
   I3 => x56_out_12,
   I4 => x56_out_8,
   O => W_59_7_i_12_n_0
);
W_59_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x32_out_4,
   I1 => x56_out_7,
   I2 => x56_out_11,
   I3 => x56_out_22,
   I4 => x59_out_4,
   O => W_59_7_i_13_n_0
);
W_59_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x59_out_4,
   I1 => x32_out_4,
   I2 => x56_out_22,
   I3 => x56_out_11,
   I4 => x56_out_7,
   O => W_59_7_i_14_n_0
);
W_59_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x32_out_3,
   I1 => x56_out_6,
   I2 => x56_out_10,
   I3 => x56_out_21,
   I4 => x59_out_3,
   O => W_59_7_i_15_n_0
);
W_59_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x59_out_3,
   I1 => x32_out_3,
   I2 => x56_out_21,
   I3 => x56_out_10,
   I4 => x56_out_6,
   O => W_59_7_i_16_n_0
);
W_59_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x32_out_2,
   I1 => x56_out_5,
   I2 => x56_out_9,
   I3 => x56_out_20,
   I4 => x59_out_2,
   O => W_59_7_i_17_n_0
);
W_59_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x17_out_16,
   I1 => x17_out_23,
   I2 => x17_out_25,
   I3 => W_59_7_i_10_n_0,
   I4 => W_59_7_i_11_n_0,
   O => W_59_7_i_2_n_0
);
W_59_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x17_out_15,
   I1 => x17_out_22,
   I2 => x17_out_24,
   I3 => W_59_7_i_12_n_0,
   I4 => W_59_7_i_13_n_0,
   O => W_59_7_i_3_n_0
);
W_59_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x17_out_14,
   I1 => x17_out_21,
   I2 => x17_out_23,
   I3 => W_59_7_i_14_n_0,
   I4 => W_59_7_i_15_n_0,
   O => W_59_7_i_4_n_0
);
W_59_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x17_out_13,
   I1 => x17_out_20,
   I2 => x17_out_22,
   I3 => W_59_7_i_16_n_0,
   I4 => W_59_7_i_17_n_0,
   O => W_59_7_i_5_n_0
);
W_59_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_59_7_i_2_n_0,
   I1 => W_59_11_i_16_n_0,
   I2 => x17_out_17,
   I3 => x17_out_24,
   I4 => x17_out_26,
   I5 => W_59_11_i_17_n_0,
   O => W_59_7_i_6_n_0
);
W_59_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_59_7_i_3_n_0,
   I1 => W_59_7_i_10_n_0,
   I2 => x17_out_16,
   I3 => x17_out_23,
   I4 => x17_out_25,
   I5 => W_59_7_i_11_n_0,
   O => W_59_7_i_7_n_0
);
W_59_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_59_7_i_4_n_0,
   I1 => W_59_7_i_12_n_0,
   I2 => x17_out_15,
   I3 => x17_out_22,
   I4 => x17_out_24,
   I5 => W_59_7_i_13_n_0,
   O => W_59_7_i_8_n_0
);
W_59_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_59_7_i_5_n_0,
   I1 => W_59_7_i_14_n_0,
   I2 => x17_out_14,
   I3 => x17_out_21,
   I4 => x17_out_23,
   I5 => W_59_7_i_15_n_0,
   O => W_59_7_i_9_n_0
);
W_60_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x56_out_10,
   I1 => x29_out_10,
   I2 => x53_out_28,
   I3 => x53_out_17,
   I4 => x53_out_13,
   O => W_60_11_i_10_n_0
);
W_60_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x29_out_9,
   I1 => x53_out_12,
   I2 => x53_out_16,
   I3 => x53_out_27,
   I4 => x56_out_9,
   O => W_60_11_i_11_n_0
);
W_60_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x56_out_9,
   I1 => x29_out_9,
   I2 => x53_out_27,
   I3 => x53_out_16,
   I4 => x53_out_12,
   O => W_60_11_i_12_n_0
);
W_60_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x29_out_8,
   I1 => x53_out_11,
   I2 => x53_out_15,
   I3 => x53_out_26,
   I4 => x56_out_8,
   O => W_60_11_i_13_n_0
);
W_60_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x56_out_8,
   I1 => x29_out_8,
   I2 => x53_out_26,
   I3 => x53_out_15,
   I4 => x53_out_11,
   O => W_60_11_i_14_n_0
);
W_60_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x29_out_7,
   I1 => x53_out_10,
   I2 => x53_out_14,
   I3 => x53_out_25,
   I4 => x56_out_7,
   O => W_60_11_i_15_n_0
);
W_60_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x56_out_7,
   I1 => x29_out_7,
   I2 => x53_out_25,
   I3 => x53_out_14,
   I4 => x53_out_10,
   O => W_60_11_i_16_n_0
);
W_60_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x29_out_6,
   I1 => x53_out_9,
   I2 => x53_out_13,
   I3 => x53_out_24,
   I4 => x56_out_6,
   O => W_60_11_i_17_n_0
);
W_60_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x14_out_20,
   I1 => x14_out_27,
   I2 => x14_out_29,
   I3 => W_60_11_i_10_n_0,
   I4 => W_60_11_i_11_n_0,
   O => W_60_11_i_2_n_0
);
W_60_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x14_out_19,
   I1 => x14_out_26,
   I2 => x14_out_28,
   I3 => W_60_11_i_12_n_0,
   I4 => W_60_11_i_13_n_0,
   O => W_60_11_i_3_n_0
);
W_60_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x14_out_18,
   I1 => x14_out_25,
   I2 => x14_out_27,
   I3 => W_60_11_i_14_n_0,
   I4 => W_60_11_i_15_n_0,
   O => W_60_11_i_4_n_0
);
W_60_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x14_out_17,
   I1 => x14_out_24,
   I2 => x14_out_26,
   I3 => W_60_11_i_16_n_0,
   I4 => W_60_11_i_17_n_0,
   O => W_60_11_i_5_n_0
);
W_60_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_60_11_i_2_n_0,
   I1 => W_60_15_i_16_n_0,
   I2 => x14_out_21,
   I3 => x14_out_28,
   I4 => x14_out_30,
   I5 => W_60_15_i_17_n_0,
   O => W_60_11_i_6_n_0
);
W_60_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_60_11_i_3_n_0,
   I1 => W_60_11_i_10_n_0,
   I2 => x14_out_20,
   I3 => x14_out_27,
   I4 => x14_out_29,
   I5 => W_60_11_i_11_n_0,
   O => W_60_11_i_7_n_0
);
W_60_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_60_11_i_4_n_0,
   I1 => W_60_11_i_12_n_0,
   I2 => x14_out_19,
   I3 => x14_out_26,
   I4 => x14_out_28,
   I5 => W_60_11_i_13_n_0,
   O => W_60_11_i_8_n_0
);
W_60_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_60_11_i_5_n_0,
   I1 => W_60_11_i_14_n_0,
   I2 => x14_out_18,
   I3 => x14_out_25,
   I4 => x14_out_27,
   I5 => W_60_11_i_15_n_0,
   O => W_60_11_i_9_n_0
);
W_60_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x56_out_14,
   I1 => x29_out_14,
   I2 => x53_out_0,
   I3 => x53_out_21,
   I4 => x53_out_17,
   O => W_60_15_i_10_n_0
);
W_60_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x29_out_13,
   I1 => x53_out_16,
   I2 => x53_out_20,
   I3 => x53_out_31,
   I4 => x56_out_13,
   O => W_60_15_i_11_n_0
);
W_60_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x56_out_13,
   I1 => x29_out_13,
   I2 => x53_out_31,
   I3 => x53_out_20,
   I4 => x53_out_16,
   O => W_60_15_i_12_n_0
);
W_60_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x29_out_12,
   I1 => x53_out_15,
   I2 => x53_out_19,
   I3 => x53_out_30,
   I4 => x56_out_12,
   O => W_60_15_i_13_n_0
);
W_60_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x56_out_12,
   I1 => x29_out_12,
   I2 => x53_out_30,
   I3 => x53_out_19,
   I4 => x53_out_15,
   O => W_60_15_i_14_n_0
);
W_60_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x29_out_11,
   I1 => x53_out_14,
   I2 => x53_out_18,
   I3 => x53_out_29,
   I4 => x56_out_11,
   O => W_60_15_i_15_n_0
);
W_60_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x56_out_11,
   I1 => x29_out_11,
   I2 => x53_out_29,
   I3 => x53_out_18,
   I4 => x53_out_14,
   O => W_60_15_i_16_n_0
);
W_60_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x29_out_10,
   I1 => x53_out_13,
   I2 => x53_out_17,
   I3 => x53_out_28,
   I4 => x56_out_10,
   O => W_60_15_i_17_n_0
);
W_60_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x14_out_24,
   I1 => x14_out_31,
   I2 => x14_out_1,
   I3 => W_60_15_i_10_n_0,
   I4 => W_60_15_i_11_n_0,
   O => W_60_15_i_2_n_0
);
W_60_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x14_out_23,
   I1 => x14_out_30,
   I2 => x14_out_0,
   I3 => W_60_15_i_12_n_0,
   I4 => W_60_15_i_13_n_0,
   O => W_60_15_i_3_n_0
);
W_60_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x14_out_22,
   I1 => x14_out_29,
   I2 => x14_out_31,
   I3 => W_60_15_i_14_n_0,
   I4 => W_60_15_i_15_n_0,
   O => W_60_15_i_4_n_0
);
W_60_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x14_out_21,
   I1 => x14_out_28,
   I2 => x14_out_30,
   I3 => W_60_15_i_16_n_0,
   I4 => W_60_15_i_17_n_0,
   O => W_60_15_i_5_n_0
);
W_60_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_60_15_i_2_n_0,
   I1 => W_60_19_i_16_n_0,
   I2 => x14_out_25,
   I3 => x14_out_0,
   I4 => x14_out_2,
   I5 => W_60_19_i_17_n_0,
   O => W_60_15_i_6_n_0
);
W_60_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_60_15_i_3_n_0,
   I1 => W_60_15_i_10_n_0,
   I2 => x14_out_24,
   I3 => x14_out_31,
   I4 => x14_out_1,
   I5 => W_60_15_i_11_n_0,
   O => W_60_15_i_7_n_0
);
W_60_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_60_15_i_4_n_0,
   I1 => W_60_15_i_12_n_0,
   I2 => x14_out_23,
   I3 => x14_out_30,
   I4 => x14_out_0,
   I5 => W_60_15_i_13_n_0,
   O => W_60_15_i_8_n_0
);
W_60_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_60_15_i_5_n_0,
   I1 => W_60_15_i_14_n_0,
   I2 => x14_out_22,
   I3 => x14_out_29,
   I4 => x14_out_31,
   I5 => W_60_15_i_15_n_0,
   O => W_60_15_i_9_n_0
);
W_60_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x56_out_18,
   I1 => x29_out_18,
   I2 => x53_out_4,
   I3 => x53_out_25,
   I4 => x53_out_21,
   O => W_60_19_i_10_n_0
);
W_60_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x29_out_17,
   I1 => x53_out_20,
   I2 => x53_out_24,
   I3 => x53_out_3,
   I4 => x56_out_17,
   O => W_60_19_i_11_n_0
);
W_60_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x56_out_17,
   I1 => x29_out_17,
   I2 => x53_out_3,
   I3 => x53_out_24,
   I4 => x53_out_20,
   O => W_60_19_i_12_n_0
);
W_60_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x29_out_16,
   I1 => x53_out_19,
   I2 => x53_out_23,
   I3 => x53_out_2,
   I4 => x56_out_16,
   O => W_60_19_i_13_n_0
);
W_60_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x56_out_16,
   I1 => x29_out_16,
   I2 => x53_out_2,
   I3 => x53_out_23,
   I4 => x53_out_19,
   O => W_60_19_i_14_n_0
);
W_60_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x29_out_15,
   I1 => x53_out_18,
   I2 => x53_out_22,
   I3 => x53_out_1,
   I4 => x56_out_15,
   O => W_60_19_i_15_n_0
);
W_60_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x56_out_15,
   I1 => x29_out_15,
   I2 => x53_out_1,
   I3 => x53_out_22,
   I4 => x53_out_18,
   O => W_60_19_i_16_n_0
);
W_60_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x29_out_14,
   I1 => x53_out_17,
   I2 => x53_out_21,
   I3 => x53_out_0,
   I4 => x56_out_14,
   O => W_60_19_i_17_n_0
);
W_60_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x14_out_28,
   I1 => x14_out_3,
   I2 => x14_out_5,
   I3 => W_60_19_i_10_n_0,
   I4 => W_60_19_i_11_n_0,
   O => W_60_19_i_2_n_0
);
W_60_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x14_out_27,
   I1 => x14_out_2,
   I2 => x14_out_4,
   I3 => W_60_19_i_12_n_0,
   I4 => W_60_19_i_13_n_0,
   O => W_60_19_i_3_n_0
);
W_60_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x14_out_26,
   I1 => x14_out_1,
   I2 => x14_out_3,
   I3 => W_60_19_i_14_n_0,
   I4 => W_60_19_i_15_n_0,
   O => W_60_19_i_4_n_0
);
W_60_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x14_out_25,
   I1 => x14_out_0,
   I2 => x14_out_2,
   I3 => W_60_19_i_16_n_0,
   I4 => W_60_19_i_17_n_0,
   O => W_60_19_i_5_n_0
);
W_60_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_60_19_i_2_n_0,
   I1 => W_60_23_i_16_n_0,
   I2 => x14_out_29,
   I3 => x14_out_4,
   I4 => x14_out_6,
   I5 => W_60_23_i_17_n_0,
   O => W_60_19_i_6_n_0
);
W_60_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_60_19_i_3_n_0,
   I1 => W_60_19_i_10_n_0,
   I2 => x14_out_28,
   I3 => x14_out_3,
   I4 => x14_out_5,
   I5 => W_60_19_i_11_n_0,
   O => W_60_19_i_7_n_0
);
W_60_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_60_19_i_4_n_0,
   I1 => W_60_19_i_12_n_0,
   I2 => x14_out_27,
   I3 => x14_out_2,
   I4 => x14_out_4,
   I5 => W_60_19_i_13_n_0,
   O => W_60_19_i_8_n_0
);
W_60_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_60_19_i_5_n_0,
   I1 => W_60_19_i_14_n_0,
   I2 => x14_out_26,
   I3 => x14_out_1,
   I4 => x14_out_3,
   I5 => W_60_19_i_15_n_0,
   O => W_60_19_i_9_n_0
);
W_60_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x56_out_22,
   I1 => x29_out_22,
   I2 => x53_out_8,
   I3 => x53_out_29,
   I4 => x53_out_25,
   O => W_60_23_i_10_n_0
);
W_60_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x29_out_21,
   I1 => x53_out_24,
   I2 => x53_out_28,
   I3 => x53_out_7,
   I4 => x56_out_21,
   O => W_60_23_i_11_n_0
);
W_60_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x56_out_21,
   I1 => x29_out_21,
   I2 => x53_out_7,
   I3 => x53_out_28,
   I4 => x53_out_24,
   O => W_60_23_i_12_n_0
);
W_60_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x29_out_20,
   I1 => x53_out_23,
   I2 => x53_out_27,
   I3 => x53_out_6,
   I4 => x56_out_20,
   O => W_60_23_i_13_n_0
);
W_60_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x56_out_20,
   I1 => x29_out_20,
   I2 => x53_out_6,
   I3 => x53_out_27,
   I4 => x53_out_23,
   O => W_60_23_i_14_n_0
);
W_60_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x29_out_19,
   I1 => x53_out_22,
   I2 => x53_out_26,
   I3 => x53_out_5,
   I4 => x56_out_19,
   O => W_60_23_i_15_n_0
);
W_60_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x56_out_19,
   I1 => x29_out_19,
   I2 => x53_out_5,
   I3 => x53_out_26,
   I4 => x53_out_22,
   O => W_60_23_i_16_n_0
);
W_60_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x29_out_18,
   I1 => x53_out_21,
   I2 => x53_out_25,
   I3 => x53_out_4,
   I4 => x56_out_18,
   O => W_60_23_i_17_n_0
);
W_60_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x14_out_7,
   I1 => x14_out_9,
   I2 => W_60_23_i_10_n_0,
   I3 => W_60_23_i_11_n_0,
   O => W_60_23_i_2_n_0
);
W_60_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x14_out_31,
   I1 => x14_out_6,
   I2 => x14_out_8,
   I3 => W_60_23_i_12_n_0,
   I4 => W_60_23_i_13_n_0,
   O => W_60_23_i_3_n_0
);
W_60_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x14_out_30,
   I1 => x14_out_5,
   I2 => x14_out_7,
   I3 => W_60_23_i_14_n_0,
   I4 => W_60_23_i_15_n_0,
   O => W_60_23_i_4_n_0
);
W_60_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x14_out_29,
   I1 => x14_out_4,
   I2 => x14_out_6,
   I3 => W_60_23_i_16_n_0,
   I4 => W_60_23_i_17_n_0,
   O => W_60_23_i_5_n_0
);
W_60_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x14_out_8,
   I1 => x14_out_10,
   I2 => W_60_27_i_16_n_0,
   I3 => W_60_27_i_17_n_0,
   I4 => W_60_23_i_2_n_0,
   O => W_60_23_i_6_n_0
);
W_60_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x14_out_7,
   I1 => x14_out_9,
   I2 => W_60_23_i_10_n_0,
   I3 => W_60_23_i_11_n_0,
   I4 => W_60_23_i_3_n_0,
   O => W_60_23_i_7_n_0
);
W_60_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_60_23_i_4_n_0,
   I1 => W_60_23_i_12_n_0,
   I2 => x14_out_31,
   I3 => x14_out_6,
   I4 => x14_out_8,
   I5 => W_60_23_i_13_n_0,
   O => W_60_23_i_8_n_0
);
W_60_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_60_23_i_5_n_0,
   I1 => W_60_23_i_14_n_0,
   I2 => x14_out_30,
   I3 => x14_out_5,
   I4 => x14_out_7,
   I5 => W_60_23_i_15_n_0,
   O => W_60_23_i_9_n_0
);
W_60_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x56_out_26,
   I1 => x29_out_26,
   I2 => x53_out_12,
   I3 => x53_out_1,
   I4 => x53_out_29,
   O => W_60_27_i_10_n_0
);
W_60_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x29_out_25,
   I1 => x53_out_28,
   I2 => x53_out_0,
   I3 => x53_out_11,
   I4 => x56_out_25,
   O => W_60_27_i_11_n_0
);
W_60_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x56_out_25,
   I1 => x29_out_25,
   I2 => x53_out_11,
   I3 => x53_out_0,
   I4 => x53_out_28,
   O => W_60_27_i_12_n_0
);
W_60_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x29_out_24,
   I1 => x53_out_27,
   I2 => x53_out_31,
   I3 => x53_out_10,
   I4 => x56_out_24,
   O => W_60_27_i_13_n_0
);
W_60_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x56_out_24,
   I1 => x29_out_24,
   I2 => x53_out_10,
   I3 => x53_out_31,
   I4 => x53_out_27,
   O => W_60_27_i_14_n_0
);
W_60_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x29_out_23,
   I1 => x53_out_26,
   I2 => x53_out_30,
   I3 => x53_out_9,
   I4 => x56_out_23,
   O => W_60_27_i_15_n_0
);
W_60_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x56_out_23,
   I1 => x29_out_23,
   I2 => x53_out_9,
   I3 => x53_out_30,
   I4 => x53_out_26,
   O => W_60_27_i_16_n_0
);
W_60_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x29_out_22,
   I1 => x53_out_25,
   I2 => x53_out_29,
   I3 => x53_out_8,
   I4 => x56_out_22,
   O => W_60_27_i_17_n_0
);
W_60_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x14_out_11,
   I1 => x14_out_13,
   I2 => W_60_27_i_10_n_0,
   I3 => W_60_27_i_11_n_0,
   O => W_60_27_i_2_n_0
);
W_60_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x14_out_10,
   I1 => x14_out_12,
   I2 => W_60_27_i_12_n_0,
   I3 => W_60_27_i_13_n_0,
   O => W_60_27_i_3_n_0
);
W_60_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x14_out_9,
   I1 => x14_out_11,
   I2 => W_60_27_i_14_n_0,
   I3 => W_60_27_i_15_n_0,
   O => W_60_27_i_4_n_0
);
W_60_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x14_out_8,
   I1 => x14_out_10,
   I2 => W_60_27_i_16_n_0,
   I3 => W_60_27_i_17_n_0,
   O => W_60_27_i_5_n_0
);
W_60_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x14_out_12,
   I1 => x14_out_14,
   I2 => W_60_31_i_13_n_0,
   I3 => W_60_31_i_14_n_0,
   I4 => W_60_27_i_2_n_0,
   O => W_60_27_i_6_n_0
);
W_60_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x14_out_11,
   I1 => x14_out_13,
   I2 => W_60_27_i_10_n_0,
   I3 => W_60_27_i_11_n_0,
   I4 => W_60_27_i_3_n_0,
   O => W_60_27_i_7_n_0
);
W_60_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x14_out_10,
   I1 => x14_out_12,
   I2 => W_60_27_i_12_n_0,
   I3 => W_60_27_i_13_n_0,
   I4 => W_60_27_i_4_n_0,
   O => W_60_27_i_8_n_0
);
W_60_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x14_out_9,
   I1 => x14_out_11,
   I2 => W_60_27_i_14_n_0,
   I3 => W_60_27_i_15_n_0,
   I4 => W_60_27_i_5_n_0,
   O => W_60_27_i_9_n_0
);
W_60_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x29_out_28,
   I1 => x53_out_31,
   I2 => x53_out_3,
   I3 => x53_out_14,
   I4 => x56_out_28,
   O => W_60_31_i_10_n_0
);
W_60_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x56_out_28,
   I1 => x29_out_28,
   I2 => x53_out_14,
   I3 => x53_out_3,
   I4 => x53_out_31,
   O => W_60_31_i_11_n_0
);
W_60_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x29_out_27,
   I1 => x53_out_30,
   I2 => x53_out_2,
   I3 => x53_out_13,
   I4 => x56_out_27,
   O => W_60_31_i_12_n_0
);
W_60_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x56_out_27,
   I1 => x29_out_27,
   I2 => x53_out_13,
   I3 => x53_out_2,
   I4 => x53_out_30,
   O => W_60_31_i_13_n_0
);
W_60_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x29_out_26,
   I1 => x53_out_29,
   I2 => x53_out_1,
   I3 => x53_out_12,
   I4 => x56_out_26,
   O => W_60_31_i_14_n_0
);
W_60_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x29_out_29,
   I1 => x53_out_4,
   I2 => x53_out_15,
   I3 => x56_out_29,
   O => W_60_31_i_15_n_0
);
W_60_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x14_out_17,
   I1 => x14_out_15,
   O => SIGMA_LCASE_135_out_0_30
);
W_60_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => x53_out_6,
   I1 => x53_out_17,
   I2 => x29_out_31,
   I3 => x56_out_31,
   I4 => x14_out_16,
   I5 => x14_out_18,
   O => W_60_31_i_17_n_0
);
W_60_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x53_out_16,
   I1 => x53_out_5,
   O => SIGMA_LCASE_031_out_30
);
W_60_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x56_out_30,
   I1 => x29_out_30,
   I2 => x53_out_16,
   I3 => x53_out_5,
   O => W_60_31_i_19_n_0
);
W_60_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x14_out_14,
   I1 => x14_out_16,
   I2 => W_60_31_i_9_n_0,
   I3 => W_60_31_i_10_n_0,
   O => W_60_31_i_2_n_0
);
W_60_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x14_out_13,
   I1 => x14_out_15,
   I2 => W_60_31_i_11_n_0,
   I3 => W_60_31_i_12_n_0,
   O => W_60_31_i_3_n_0
);
W_60_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x14_out_12,
   I1 => x14_out_14,
   I2 => W_60_31_i_13_n_0,
   I3 => W_60_31_i_14_n_0,
   O => W_60_31_i_4_n_0
);
W_60_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_60_31_i_15_n_0,
   I1 => SIGMA_LCASE_135_out_0_30,
   I2 => W_60_31_i_17_n_0,
   I3 => x29_out_30,
   I4 => SIGMA_LCASE_031_out_30,
   I5 => x56_out_30,
   O => W_60_31_i_5_n_0
);
W_60_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_60_31_i_2_n_0,
   I1 => W_60_31_i_19_n_0,
   I2 => x14_out_15,
   I3 => x14_out_17,
   I4 => W_60_31_i_15_n_0,
   O => W_60_31_i_6_n_0
);
W_60_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x14_out_14,
   I1 => x14_out_16,
   I2 => W_60_31_i_9_n_0,
   I3 => W_60_31_i_10_n_0,
   I4 => W_60_31_i_3_n_0,
   O => W_60_31_i_7_n_0
);
W_60_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x14_out_13,
   I1 => x14_out_15,
   I2 => W_60_31_i_11_n_0,
   I3 => W_60_31_i_12_n_0,
   I4 => W_60_31_i_4_n_0,
   O => W_60_31_i_8_n_0
);
W_60_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x56_out_29,
   I1 => x29_out_29,
   I2 => x53_out_15,
   I3 => x53_out_4,
   O => W_60_31_i_9_n_0
);
W_60_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x56_out_2,
   I1 => x29_out_2,
   I2 => x53_out_20,
   I3 => x53_out_9,
   I4 => x53_out_5,
   O => W_60_3_i_10_n_0
);
W_60_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x29_out_1,
   I1 => x53_out_4,
   I2 => x53_out_8,
   I3 => x53_out_19,
   I4 => x56_out_1,
   O => W_60_3_i_11_n_0
);
W_60_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x53_out_19,
   I1 => x53_out_8,
   I2 => x53_out_4,
   O => SIGMA_LCASE_031_out_1
);
W_60_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x14_out_21,
   I1 => x14_out_19,
   I2 => x14_out_12,
   O => SIGMA_LCASE_135_out_0_2
);
W_60_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x14_out_20,
   I1 => x14_out_18,
   I2 => x14_out_11,
   O => SIGMA_LCASE_135_out_1
);
W_60_3_i_15 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x56_out_1,
   I1 => x29_out_1,
   I2 => x53_out_19,
   I3 => x53_out_8,
   I4 => x53_out_4,
   O => W_60_3_i_15_n_0
);
W_60_3_i_16 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x53_out_18,
   I1 => x53_out_7,
   I2 => x53_out_3,
   O => SIGMA_LCASE_031_out_0
);
W_60_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x14_out_12,
   I1 => x14_out_19,
   I2 => x14_out_21,
   I3 => W_60_3_i_10_n_0,
   I4 => W_60_3_i_11_n_0,
   O => W_60_3_i_2_n_0
);
W_60_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_60_3_i_11_n_0,
   I1 => x14_out_21,
   I2 => x14_out_19,
   I3 => x14_out_12,
   I4 => W_60_3_i_10_n_0,
   O => W_60_3_i_3_n_0
);
W_60_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_031_out_1,
   I1 => x29_out_1,
   I2 => x56_out_1,
   I3 => x14_out_11,
   I4 => x14_out_18,
   I5 => x14_out_20,
   O => W_60_3_i_4_n_0
);
W_60_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x56_out_0,
   I1 => x29_out_0,
   I2 => x53_out_18,
   I3 => x53_out_7,
   I4 => x53_out_3,
   O => W_60_3_i_5_n_0
);
W_60_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_60_3_i_2_n_0,
   I1 => W_60_7_i_16_n_0,
   I2 => x14_out_13,
   I3 => x14_out_20,
   I4 => x14_out_22,
   I5 => W_60_7_i_17_n_0,
   O => W_60_3_i_6_n_0
);
W_60_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_60_3_i_10_n_0,
   I1 => SIGMA_LCASE_135_out_0_2,
   I2 => x56_out_1,
   I3 => x29_out_1,
   I4 => SIGMA_LCASE_031_out_1,
   I5 => SIGMA_LCASE_135_out_1,
   O => W_60_3_i_7_n_0
);
W_60_3_i_8 : LUT5
  generic map(
   INIT => X"99969666"
  )
 port map (
   I0 => SIGMA_LCASE_135_out_1,
   I1 => W_60_3_i_15_n_0,
   I2 => x56_out_0,
   I3 => SIGMA_LCASE_031_out_0,
   I4 => x29_out_0,
   O => W_60_3_i_8_n_0
);
W_60_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_60_3_i_5_n_0,
   I1 => x14_out_10,
   I2 => x14_out_17,
   I3 => x14_out_19,
   O => W_60_3_i_9_n_0
);
W_60_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x56_out_6,
   I1 => x29_out_6,
   I2 => x53_out_24,
   I3 => x53_out_13,
   I4 => x53_out_9,
   O => W_60_7_i_10_n_0
);
W_60_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x29_out_5,
   I1 => x53_out_8,
   I2 => x53_out_12,
   I3 => x53_out_23,
   I4 => x56_out_5,
   O => W_60_7_i_11_n_0
);
W_60_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x56_out_5,
   I1 => x29_out_5,
   I2 => x53_out_23,
   I3 => x53_out_12,
   I4 => x53_out_8,
   O => W_60_7_i_12_n_0
);
W_60_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x29_out_4,
   I1 => x53_out_7,
   I2 => x53_out_11,
   I3 => x53_out_22,
   I4 => x56_out_4,
   O => W_60_7_i_13_n_0
);
W_60_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x56_out_4,
   I1 => x29_out_4,
   I2 => x53_out_22,
   I3 => x53_out_11,
   I4 => x53_out_7,
   O => W_60_7_i_14_n_0
);
W_60_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x29_out_3,
   I1 => x53_out_6,
   I2 => x53_out_10,
   I3 => x53_out_21,
   I4 => x56_out_3,
   O => W_60_7_i_15_n_0
);
W_60_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x56_out_3,
   I1 => x29_out_3,
   I2 => x53_out_21,
   I3 => x53_out_10,
   I4 => x53_out_6,
   O => W_60_7_i_16_n_0
);
W_60_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x29_out_2,
   I1 => x53_out_5,
   I2 => x53_out_9,
   I3 => x53_out_20,
   I4 => x56_out_2,
   O => W_60_7_i_17_n_0
);
W_60_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x14_out_16,
   I1 => x14_out_23,
   I2 => x14_out_25,
   I3 => W_60_7_i_10_n_0,
   I4 => W_60_7_i_11_n_0,
   O => W_60_7_i_2_n_0
);
W_60_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x14_out_15,
   I1 => x14_out_22,
   I2 => x14_out_24,
   I3 => W_60_7_i_12_n_0,
   I4 => W_60_7_i_13_n_0,
   O => W_60_7_i_3_n_0
);
W_60_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x14_out_14,
   I1 => x14_out_21,
   I2 => x14_out_23,
   I3 => W_60_7_i_14_n_0,
   I4 => W_60_7_i_15_n_0,
   O => W_60_7_i_4_n_0
);
W_60_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x14_out_13,
   I1 => x14_out_20,
   I2 => x14_out_22,
   I3 => W_60_7_i_16_n_0,
   I4 => W_60_7_i_17_n_0,
   O => W_60_7_i_5_n_0
);
W_60_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_60_7_i_2_n_0,
   I1 => W_60_11_i_16_n_0,
   I2 => x14_out_17,
   I3 => x14_out_24,
   I4 => x14_out_26,
   I5 => W_60_11_i_17_n_0,
   O => W_60_7_i_6_n_0
);
W_60_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_60_7_i_3_n_0,
   I1 => W_60_7_i_10_n_0,
   I2 => x14_out_16,
   I3 => x14_out_23,
   I4 => x14_out_25,
   I5 => W_60_7_i_11_n_0,
   O => W_60_7_i_7_n_0
);
W_60_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_60_7_i_4_n_0,
   I1 => W_60_7_i_12_n_0,
   I2 => x14_out_15,
   I3 => x14_out_22,
   I4 => x14_out_24,
   I5 => W_60_7_i_13_n_0,
   O => W_60_7_i_8_n_0
);
W_60_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_60_7_i_5_n_0,
   I1 => W_60_7_i_14_n_0,
   I2 => x14_out_14,
   I3 => x14_out_21,
   I4 => x14_out_23,
   I5 => W_60_7_i_15_n_0,
   O => W_60_7_i_9_n_0
);
W_61_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x53_out_10,
   I1 => x26_out_10,
   I2 => x50_out_28,
   I3 => x50_out_17,
   I4 => x50_out_13,
   O => W_61_11_i_10_n_0
);
W_61_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x26_out_9,
   I1 => x50_out_12,
   I2 => x50_out_16,
   I3 => x50_out_27,
   I4 => x53_out_9,
   O => W_61_11_i_11_n_0
);
W_61_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x53_out_9,
   I1 => x26_out_9,
   I2 => x50_out_27,
   I3 => x50_out_16,
   I4 => x50_out_12,
   O => W_61_11_i_12_n_0
);
W_61_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x26_out_8,
   I1 => x50_out_11,
   I2 => x50_out_15,
   I3 => x50_out_26,
   I4 => x53_out_8,
   O => W_61_11_i_13_n_0
);
W_61_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x53_out_8,
   I1 => x26_out_8,
   I2 => x50_out_26,
   I3 => x50_out_15,
   I4 => x50_out_11,
   O => W_61_11_i_14_n_0
);
W_61_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x26_out_7,
   I1 => x50_out_10,
   I2 => x50_out_14,
   I3 => x50_out_25,
   I4 => x53_out_7,
   O => W_61_11_i_15_n_0
);
W_61_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x53_out_7,
   I1 => x26_out_7,
   I2 => x50_out_25,
   I3 => x50_out_14,
   I4 => x50_out_10,
   O => W_61_11_i_16_n_0
);
W_61_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x26_out_6,
   I1 => x50_out_9,
   I2 => x50_out_13,
   I3 => x50_out_24,
   I4 => x53_out_6,
   O => W_61_11_i_17_n_0
);
W_61_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x11_out_20,
   I1 => x11_out_27,
   I2 => x11_out_29,
   I3 => W_61_11_i_10_n_0,
   I4 => W_61_11_i_11_n_0,
   O => W_61_11_i_2_n_0
);
W_61_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x11_out_19,
   I1 => x11_out_26,
   I2 => x11_out_28,
   I3 => W_61_11_i_12_n_0,
   I4 => W_61_11_i_13_n_0,
   O => W_61_11_i_3_n_0
);
W_61_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x11_out_18,
   I1 => x11_out_25,
   I2 => x11_out_27,
   I3 => W_61_11_i_14_n_0,
   I4 => W_61_11_i_15_n_0,
   O => W_61_11_i_4_n_0
);
W_61_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x11_out_17,
   I1 => x11_out_24,
   I2 => x11_out_26,
   I3 => W_61_11_i_16_n_0,
   I4 => W_61_11_i_17_n_0,
   O => W_61_11_i_5_n_0
);
W_61_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_61_11_i_2_n_0,
   I1 => W_61_15_i_16_n_0,
   I2 => x11_out_21,
   I3 => x11_out_28,
   I4 => x11_out_30,
   I5 => W_61_15_i_17_n_0,
   O => W_61_11_i_6_n_0
);
W_61_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_61_11_i_3_n_0,
   I1 => W_61_11_i_10_n_0,
   I2 => x11_out_20,
   I3 => x11_out_27,
   I4 => x11_out_29,
   I5 => W_61_11_i_11_n_0,
   O => W_61_11_i_7_n_0
);
W_61_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_61_11_i_4_n_0,
   I1 => W_61_11_i_12_n_0,
   I2 => x11_out_19,
   I3 => x11_out_26,
   I4 => x11_out_28,
   I5 => W_61_11_i_13_n_0,
   O => W_61_11_i_8_n_0
);
W_61_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_61_11_i_5_n_0,
   I1 => W_61_11_i_14_n_0,
   I2 => x11_out_18,
   I3 => x11_out_25,
   I4 => x11_out_27,
   I5 => W_61_11_i_15_n_0,
   O => W_61_11_i_9_n_0
);
W_61_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x53_out_14,
   I1 => x26_out_14,
   I2 => x50_out_0,
   I3 => x50_out_21,
   I4 => x50_out_17,
   O => W_61_15_i_10_n_0
);
W_61_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x26_out_13,
   I1 => x50_out_16,
   I2 => x50_out_20,
   I3 => x50_out_31,
   I4 => x53_out_13,
   O => W_61_15_i_11_n_0
);
W_61_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x53_out_13,
   I1 => x26_out_13,
   I2 => x50_out_31,
   I3 => x50_out_20,
   I4 => x50_out_16,
   O => W_61_15_i_12_n_0
);
W_61_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x26_out_12,
   I1 => x50_out_15,
   I2 => x50_out_19,
   I3 => x50_out_30,
   I4 => x53_out_12,
   O => W_61_15_i_13_n_0
);
W_61_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x53_out_12,
   I1 => x26_out_12,
   I2 => x50_out_30,
   I3 => x50_out_19,
   I4 => x50_out_15,
   O => W_61_15_i_14_n_0
);
W_61_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x26_out_11,
   I1 => x50_out_14,
   I2 => x50_out_18,
   I3 => x50_out_29,
   I4 => x53_out_11,
   O => W_61_15_i_15_n_0
);
W_61_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x53_out_11,
   I1 => x26_out_11,
   I2 => x50_out_29,
   I3 => x50_out_18,
   I4 => x50_out_14,
   O => W_61_15_i_16_n_0
);
W_61_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x26_out_10,
   I1 => x50_out_13,
   I2 => x50_out_17,
   I3 => x50_out_28,
   I4 => x53_out_10,
   O => W_61_15_i_17_n_0
);
W_61_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x11_out_24,
   I1 => x11_out_31,
   I2 => x11_out_1,
   I3 => W_61_15_i_10_n_0,
   I4 => W_61_15_i_11_n_0,
   O => W_61_15_i_2_n_0
);
W_61_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x11_out_23,
   I1 => x11_out_30,
   I2 => x11_out_0,
   I3 => W_61_15_i_12_n_0,
   I4 => W_61_15_i_13_n_0,
   O => W_61_15_i_3_n_0
);
W_61_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x11_out_22,
   I1 => x11_out_29,
   I2 => x11_out_31,
   I3 => W_61_15_i_14_n_0,
   I4 => W_61_15_i_15_n_0,
   O => W_61_15_i_4_n_0
);
W_61_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x11_out_21,
   I1 => x11_out_28,
   I2 => x11_out_30,
   I3 => W_61_15_i_16_n_0,
   I4 => W_61_15_i_17_n_0,
   O => W_61_15_i_5_n_0
);
W_61_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_61_15_i_2_n_0,
   I1 => W_61_19_i_16_n_0,
   I2 => x11_out_25,
   I3 => x11_out_0,
   I4 => x11_out_2,
   I5 => W_61_19_i_17_n_0,
   O => W_61_15_i_6_n_0
);
W_61_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_61_15_i_3_n_0,
   I1 => W_61_15_i_10_n_0,
   I2 => x11_out_24,
   I3 => x11_out_31,
   I4 => x11_out_1,
   I5 => W_61_15_i_11_n_0,
   O => W_61_15_i_7_n_0
);
W_61_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_61_15_i_4_n_0,
   I1 => W_61_15_i_12_n_0,
   I2 => x11_out_23,
   I3 => x11_out_30,
   I4 => x11_out_0,
   I5 => W_61_15_i_13_n_0,
   O => W_61_15_i_8_n_0
);
W_61_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_61_15_i_5_n_0,
   I1 => W_61_15_i_14_n_0,
   I2 => x11_out_22,
   I3 => x11_out_29,
   I4 => x11_out_31,
   I5 => W_61_15_i_15_n_0,
   O => W_61_15_i_9_n_0
);
W_61_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x53_out_18,
   I1 => x26_out_18,
   I2 => x50_out_4,
   I3 => x50_out_25,
   I4 => x50_out_21,
   O => W_61_19_i_10_n_0
);
W_61_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x26_out_17,
   I1 => x50_out_20,
   I2 => x50_out_24,
   I3 => x50_out_3,
   I4 => x53_out_17,
   O => W_61_19_i_11_n_0
);
W_61_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x53_out_17,
   I1 => x26_out_17,
   I2 => x50_out_3,
   I3 => x50_out_24,
   I4 => x50_out_20,
   O => W_61_19_i_12_n_0
);
W_61_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x26_out_16,
   I1 => x50_out_19,
   I2 => x50_out_23,
   I3 => x50_out_2,
   I4 => x53_out_16,
   O => W_61_19_i_13_n_0
);
W_61_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x53_out_16,
   I1 => x26_out_16,
   I2 => x50_out_2,
   I3 => x50_out_23,
   I4 => x50_out_19,
   O => W_61_19_i_14_n_0
);
W_61_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x26_out_15,
   I1 => x50_out_18,
   I2 => x50_out_22,
   I3 => x50_out_1,
   I4 => x53_out_15,
   O => W_61_19_i_15_n_0
);
W_61_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x53_out_15,
   I1 => x26_out_15,
   I2 => x50_out_1,
   I3 => x50_out_22,
   I4 => x50_out_18,
   O => W_61_19_i_16_n_0
);
W_61_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x26_out_14,
   I1 => x50_out_17,
   I2 => x50_out_21,
   I3 => x50_out_0,
   I4 => x53_out_14,
   O => W_61_19_i_17_n_0
);
W_61_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x11_out_28,
   I1 => x11_out_3,
   I2 => x11_out_5,
   I3 => W_61_19_i_10_n_0,
   I4 => W_61_19_i_11_n_0,
   O => W_61_19_i_2_n_0
);
W_61_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x11_out_27,
   I1 => x11_out_2,
   I2 => x11_out_4,
   I3 => W_61_19_i_12_n_0,
   I4 => W_61_19_i_13_n_0,
   O => W_61_19_i_3_n_0
);
W_61_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x11_out_26,
   I1 => x11_out_1,
   I2 => x11_out_3,
   I3 => W_61_19_i_14_n_0,
   I4 => W_61_19_i_15_n_0,
   O => W_61_19_i_4_n_0
);
W_61_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x11_out_25,
   I1 => x11_out_0,
   I2 => x11_out_2,
   I3 => W_61_19_i_16_n_0,
   I4 => W_61_19_i_17_n_0,
   O => W_61_19_i_5_n_0
);
W_61_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_61_19_i_2_n_0,
   I1 => W_61_23_i_16_n_0,
   I2 => x11_out_29,
   I3 => x11_out_4,
   I4 => x11_out_6,
   I5 => W_61_23_i_17_n_0,
   O => W_61_19_i_6_n_0
);
W_61_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_61_19_i_3_n_0,
   I1 => W_61_19_i_10_n_0,
   I2 => x11_out_28,
   I3 => x11_out_3,
   I4 => x11_out_5,
   I5 => W_61_19_i_11_n_0,
   O => W_61_19_i_7_n_0
);
W_61_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_61_19_i_4_n_0,
   I1 => W_61_19_i_12_n_0,
   I2 => x11_out_27,
   I3 => x11_out_2,
   I4 => x11_out_4,
   I5 => W_61_19_i_13_n_0,
   O => W_61_19_i_8_n_0
);
W_61_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_61_19_i_5_n_0,
   I1 => W_61_19_i_14_n_0,
   I2 => x11_out_26,
   I3 => x11_out_1,
   I4 => x11_out_3,
   I5 => W_61_19_i_15_n_0,
   O => W_61_19_i_9_n_0
);
W_61_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x53_out_22,
   I1 => x26_out_22,
   I2 => x50_out_8,
   I3 => x50_out_29,
   I4 => x50_out_25,
   O => W_61_23_i_10_n_0
);
W_61_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x26_out_21,
   I1 => x50_out_24,
   I2 => x50_out_28,
   I3 => x50_out_7,
   I4 => x53_out_21,
   O => W_61_23_i_11_n_0
);
W_61_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x53_out_21,
   I1 => x26_out_21,
   I2 => x50_out_7,
   I3 => x50_out_28,
   I4 => x50_out_24,
   O => W_61_23_i_12_n_0
);
W_61_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x26_out_20,
   I1 => x50_out_23,
   I2 => x50_out_27,
   I3 => x50_out_6,
   I4 => x53_out_20,
   O => W_61_23_i_13_n_0
);
W_61_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x53_out_20,
   I1 => x26_out_20,
   I2 => x50_out_6,
   I3 => x50_out_27,
   I4 => x50_out_23,
   O => W_61_23_i_14_n_0
);
W_61_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x26_out_19,
   I1 => x50_out_22,
   I2 => x50_out_26,
   I3 => x50_out_5,
   I4 => x53_out_19,
   O => W_61_23_i_15_n_0
);
W_61_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x53_out_19,
   I1 => x26_out_19,
   I2 => x50_out_5,
   I3 => x50_out_26,
   I4 => x50_out_22,
   O => W_61_23_i_16_n_0
);
W_61_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x26_out_18,
   I1 => x50_out_21,
   I2 => x50_out_25,
   I3 => x50_out_4,
   I4 => x53_out_18,
   O => W_61_23_i_17_n_0
);
W_61_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x11_out_7,
   I1 => x11_out_9,
   I2 => W_61_23_i_10_n_0,
   I3 => W_61_23_i_11_n_0,
   O => W_61_23_i_2_n_0
);
W_61_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x11_out_31,
   I1 => x11_out_6,
   I2 => x11_out_8,
   I3 => W_61_23_i_12_n_0,
   I4 => W_61_23_i_13_n_0,
   O => W_61_23_i_3_n_0
);
W_61_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x11_out_30,
   I1 => x11_out_5,
   I2 => x11_out_7,
   I3 => W_61_23_i_14_n_0,
   I4 => W_61_23_i_15_n_0,
   O => W_61_23_i_4_n_0
);
W_61_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x11_out_29,
   I1 => x11_out_4,
   I2 => x11_out_6,
   I3 => W_61_23_i_16_n_0,
   I4 => W_61_23_i_17_n_0,
   O => W_61_23_i_5_n_0
);
W_61_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x11_out_8,
   I1 => x11_out_10,
   I2 => W_61_27_i_16_n_0,
   I3 => W_61_27_i_17_n_0,
   I4 => W_61_23_i_2_n_0,
   O => W_61_23_i_6_n_0
);
W_61_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x11_out_7,
   I1 => x11_out_9,
   I2 => W_61_23_i_10_n_0,
   I3 => W_61_23_i_11_n_0,
   I4 => W_61_23_i_3_n_0,
   O => W_61_23_i_7_n_0
);
W_61_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_61_23_i_4_n_0,
   I1 => W_61_23_i_12_n_0,
   I2 => x11_out_31,
   I3 => x11_out_6,
   I4 => x11_out_8,
   I5 => W_61_23_i_13_n_0,
   O => W_61_23_i_8_n_0
);
W_61_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_61_23_i_5_n_0,
   I1 => W_61_23_i_14_n_0,
   I2 => x11_out_30,
   I3 => x11_out_5,
   I4 => x11_out_7,
   I5 => W_61_23_i_15_n_0,
   O => W_61_23_i_9_n_0
);
W_61_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x53_out_26,
   I1 => x26_out_26,
   I2 => x50_out_12,
   I3 => x50_out_1,
   I4 => x50_out_29,
   O => W_61_27_i_10_n_0
);
W_61_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x26_out_25,
   I1 => x50_out_28,
   I2 => x50_out_0,
   I3 => x50_out_11,
   I4 => x53_out_25,
   O => W_61_27_i_11_n_0
);
W_61_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x53_out_25,
   I1 => x26_out_25,
   I2 => x50_out_11,
   I3 => x50_out_0,
   I4 => x50_out_28,
   O => W_61_27_i_12_n_0
);
W_61_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x26_out_24,
   I1 => x50_out_27,
   I2 => x50_out_31,
   I3 => x50_out_10,
   I4 => x53_out_24,
   O => W_61_27_i_13_n_0
);
W_61_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x53_out_24,
   I1 => x26_out_24,
   I2 => x50_out_10,
   I3 => x50_out_31,
   I4 => x50_out_27,
   O => W_61_27_i_14_n_0
);
W_61_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x26_out_23,
   I1 => x50_out_26,
   I2 => x50_out_30,
   I3 => x50_out_9,
   I4 => x53_out_23,
   O => W_61_27_i_15_n_0
);
W_61_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x53_out_23,
   I1 => x26_out_23,
   I2 => x50_out_9,
   I3 => x50_out_30,
   I4 => x50_out_26,
   O => W_61_27_i_16_n_0
);
W_61_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x26_out_22,
   I1 => x50_out_25,
   I2 => x50_out_29,
   I3 => x50_out_8,
   I4 => x53_out_22,
   O => W_61_27_i_17_n_0
);
W_61_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x11_out_11,
   I1 => x11_out_13,
   I2 => W_61_27_i_10_n_0,
   I3 => W_61_27_i_11_n_0,
   O => W_61_27_i_2_n_0
);
W_61_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x11_out_10,
   I1 => x11_out_12,
   I2 => W_61_27_i_12_n_0,
   I3 => W_61_27_i_13_n_0,
   O => W_61_27_i_3_n_0
);
W_61_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x11_out_9,
   I1 => x11_out_11,
   I2 => W_61_27_i_14_n_0,
   I3 => W_61_27_i_15_n_0,
   O => W_61_27_i_4_n_0
);
W_61_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x11_out_8,
   I1 => x11_out_10,
   I2 => W_61_27_i_16_n_0,
   I3 => W_61_27_i_17_n_0,
   O => W_61_27_i_5_n_0
);
W_61_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x11_out_12,
   I1 => x11_out_14,
   I2 => W_61_31_i_13_n_0,
   I3 => W_61_31_i_14_n_0,
   I4 => W_61_27_i_2_n_0,
   O => W_61_27_i_6_n_0
);
W_61_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x11_out_11,
   I1 => x11_out_13,
   I2 => W_61_27_i_10_n_0,
   I3 => W_61_27_i_11_n_0,
   I4 => W_61_27_i_3_n_0,
   O => W_61_27_i_7_n_0
);
W_61_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x11_out_10,
   I1 => x11_out_12,
   I2 => W_61_27_i_12_n_0,
   I3 => W_61_27_i_13_n_0,
   I4 => W_61_27_i_4_n_0,
   O => W_61_27_i_8_n_0
);
W_61_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x11_out_9,
   I1 => x11_out_11,
   I2 => W_61_27_i_14_n_0,
   I3 => W_61_27_i_15_n_0,
   I4 => W_61_27_i_5_n_0,
   O => W_61_27_i_9_n_0
);
W_61_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x26_out_28,
   I1 => x50_out_31,
   I2 => x50_out_3,
   I3 => x50_out_14,
   I4 => x53_out_28,
   O => W_61_31_i_10_n_0
);
W_61_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x53_out_28,
   I1 => x26_out_28,
   I2 => x50_out_14,
   I3 => x50_out_3,
   I4 => x50_out_31,
   O => W_61_31_i_11_n_0
);
W_61_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x26_out_27,
   I1 => x50_out_30,
   I2 => x50_out_2,
   I3 => x50_out_13,
   I4 => x53_out_27,
   O => W_61_31_i_12_n_0
);
W_61_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x53_out_27,
   I1 => x26_out_27,
   I2 => x50_out_13,
   I3 => x50_out_2,
   I4 => x50_out_30,
   O => W_61_31_i_13_n_0
);
W_61_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x26_out_26,
   I1 => x50_out_29,
   I2 => x50_out_1,
   I3 => x50_out_12,
   I4 => x53_out_26,
   O => W_61_31_i_14_n_0
);
W_61_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x26_out_29,
   I1 => x50_out_4,
   I2 => x50_out_15,
   I3 => x53_out_29,
   O => W_61_31_i_15_n_0
);
W_61_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x11_out_17,
   I1 => x11_out_15,
   O => SIGMA_LCASE_127_out_0_30
);
W_61_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => x50_out_6,
   I1 => x50_out_17,
   I2 => x26_out_31,
   I3 => x53_out_31,
   I4 => x11_out_16,
   I5 => x11_out_18,
   O => W_61_31_i_17_n_0
);
W_61_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x50_out_16,
   I1 => x50_out_5,
   O => SIGMA_LCASE_023_out_30
);
W_61_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x53_out_30,
   I1 => x26_out_30,
   I2 => x50_out_16,
   I3 => x50_out_5,
   O => W_61_31_i_19_n_0
);
W_61_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x11_out_14,
   I1 => x11_out_16,
   I2 => W_61_31_i_9_n_0,
   I3 => W_61_31_i_10_n_0,
   O => W_61_31_i_2_n_0
);
W_61_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x11_out_13,
   I1 => x11_out_15,
   I2 => W_61_31_i_11_n_0,
   I3 => W_61_31_i_12_n_0,
   O => W_61_31_i_3_n_0
);
W_61_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x11_out_12,
   I1 => x11_out_14,
   I2 => W_61_31_i_13_n_0,
   I3 => W_61_31_i_14_n_0,
   O => W_61_31_i_4_n_0
);
W_61_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_61_31_i_15_n_0,
   I1 => SIGMA_LCASE_127_out_0_30,
   I2 => W_61_31_i_17_n_0,
   I3 => x26_out_30,
   I4 => SIGMA_LCASE_023_out_30,
   I5 => x53_out_30,
   O => W_61_31_i_5_n_0
);
W_61_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_61_31_i_2_n_0,
   I1 => W_61_31_i_19_n_0,
   I2 => x11_out_15,
   I3 => x11_out_17,
   I4 => W_61_31_i_15_n_0,
   O => W_61_31_i_6_n_0
);
W_61_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x11_out_14,
   I1 => x11_out_16,
   I2 => W_61_31_i_9_n_0,
   I3 => W_61_31_i_10_n_0,
   I4 => W_61_31_i_3_n_0,
   O => W_61_31_i_7_n_0
);
W_61_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x11_out_13,
   I1 => x11_out_15,
   I2 => W_61_31_i_11_n_0,
   I3 => W_61_31_i_12_n_0,
   I4 => W_61_31_i_4_n_0,
   O => W_61_31_i_8_n_0
);
W_61_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x53_out_29,
   I1 => x26_out_29,
   I2 => x50_out_15,
   I3 => x50_out_4,
   O => W_61_31_i_9_n_0
);
W_61_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x53_out_2,
   I1 => x26_out_2,
   I2 => x50_out_20,
   I3 => x50_out_9,
   I4 => x50_out_5,
   O => W_61_3_i_10_n_0
);
W_61_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x26_out_1,
   I1 => x50_out_4,
   I2 => x50_out_8,
   I3 => x50_out_19,
   I4 => x53_out_1,
   O => W_61_3_i_11_n_0
);
W_61_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x50_out_19,
   I1 => x50_out_8,
   I2 => x50_out_4,
   O => SIGMA_LCASE_023_out_1
);
W_61_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x11_out_21,
   I1 => x11_out_19,
   I2 => x11_out_12,
   O => SIGMA_LCASE_127_out_0_2
);
W_61_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x11_out_20,
   I1 => x11_out_18,
   I2 => x11_out_11,
   O => SIGMA_LCASE_127_out_1
);
W_61_3_i_15 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x53_out_1,
   I1 => x26_out_1,
   I2 => x50_out_19,
   I3 => x50_out_8,
   I4 => x50_out_4,
   O => W_61_3_i_15_n_0
);
W_61_3_i_16 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x50_out_18,
   I1 => x50_out_7,
   I2 => x50_out_3,
   O => SIGMA_LCASE_023_out_0
);
W_61_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x11_out_12,
   I1 => x11_out_19,
   I2 => x11_out_21,
   I3 => W_61_3_i_10_n_0,
   I4 => W_61_3_i_11_n_0,
   O => W_61_3_i_2_n_0
);
W_61_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_61_3_i_11_n_0,
   I1 => x11_out_21,
   I2 => x11_out_19,
   I3 => x11_out_12,
   I4 => W_61_3_i_10_n_0,
   O => W_61_3_i_3_n_0
);
W_61_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_023_out_1,
   I1 => x26_out_1,
   I2 => x53_out_1,
   I3 => x11_out_11,
   I4 => x11_out_18,
   I5 => x11_out_20,
   O => W_61_3_i_4_n_0
);
W_61_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x53_out_0,
   I1 => x26_out_0,
   I2 => x50_out_18,
   I3 => x50_out_7,
   I4 => x50_out_3,
   O => W_61_3_i_5_n_0
);
W_61_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_61_3_i_2_n_0,
   I1 => W_61_7_i_16_n_0,
   I2 => x11_out_13,
   I3 => x11_out_20,
   I4 => x11_out_22,
   I5 => W_61_7_i_17_n_0,
   O => W_61_3_i_6_n_0
);
W_61_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_61_3_i_10_n_0,
   I1 => SIGMA_LCASE_127_out_0_2,
   I2 => x53_out_1,
   I3 => x26_out_1,
   I4 => SIGMA_LCASE_023_out_1,
   I5 => SIGMA_LCASE_127_out_1,
   O => W_61_3_i_7_n_0
);
W_61_3_i_8 : LUT5
  generic map(
   INIT => X"99969666"
  )
 port map (
   I0 => SIGMA_LCASE_127_out_1,
   I1 => W_61_3_i_15_n_0,
   I2 => x53_out_0,
   I3 => SIGMA_LCASE_023_out_0,
   I4 => x26_out_0,
   O => W_61_3_i_8_n_0
);
W_61_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_61_3_i_5_n_0,
   I1 => x11_out_10,
   I2 => x11_out_17,
   I3 => x11_out_19,
   O => W_61_3_i_9_n_0
);
W_61_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x53_out_6,
   I1 => x26_out_6,
   I2 => x50_out_24,
   I3 => x50_out_13,
   I4 => x50_out_9,
   O => W_61_7_i_10_n_0
);
W_61_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x26_out_5,
   I1 => x50_out_8,
   I2 => x50_out_12,
   I3 => x50_out_23,
   I4 => x53_out_5,
   O => W_61_7_i_11_n_0
);
W_61_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x53_out_5,
   I1 => x26_out_5,
   I2 => x50_out_23,
   I3 => x50_out_12,
   I4 => x50_out_8,
   O => W_61_7_i_12_n_0
);
W_61_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x26_out_4,
   I1 => x50_out_7,
   I2 => x50_out_11,
   I3 => x50_out_22,
   I4 => x53_out_4,
   O => W_61_7_i_13_n_0
);
W_61_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x53_out_4,
   I1 => x26_out_4,
   I2 => x50_out_22,
   I3 => x50_out_11,
   I4 => x50_out_7,
   O => W_61_7_i_14_n_0
);
W_61_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x26_out_3,
   I1 => x50_out_6,
   I2 => x50_out_10,
   I3 => x50_out_21,
   I4 => x53_out_3,
   O => W_61_7_i_15_n_0
);
W_61_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x53_out_3,
   I1 => x26_out_3,
   I2 => x50_out_21,
   I3 => x50_out_10,
   I4 => x50_out_6,
   O => W_61_7_i_16_n_0
);
W_61_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x26_out_2,
   I1 => x50_out_5,
   I2 => x50_out_9,
   I3 => x50_out_20,
   I4 => x53_out_2,
   O => W_61_7_i_17_n_0
);
W_61_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x11_out_16,
   I1 => x11_out_23,
   I2 => x11_out_25,
   I3 => W_61_7_i_10_n_0,
   I4 => W_61_7_i_11_n_0,
   O => W_61_7_i_2_n_0
);
W_61_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x11_out_15,
   I1 => x11_out_22,
   I2 => x11_out_24,
   I3 => W_61_7_i_12_n_0,
   I4 => W_61_7_i_13_n_0,
   O => W_61_7_i_3_n_0
);
W_61_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x11_out_14,
   I1 => x11_out_21,
   I2 => x11_out_23,
   I3 => W_61_7_i_14_n_0,
   I4 => W_61_7_i_15_n_0,
   O => W_61_7_i_4_n_0
);
W_61_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x11_out_13,
   I1 => x11_out_20,
   I2 => x11_out_22,
   I3 => W_61_7_i_16_n_0,
   I4 => W_61_7_i_17_n_0,
   O => W_61_7_i_5_n_0
);
W_61_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_61_7_i_2_n_0,
   I1 => W_61_11_i_16_n_0,
   I2 => x11_out_17,
   I3 => x11_out_24,
   I4 => x11_out_26,
   I5 => W_61_11_i_17_n_0,
   O => W_61_7_i_6_n_0
);
W_61_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_61_7_i_3_n_0,
   I1 => W_61_7_i_10_n_0,
   I2 => x11_out_16,
   I3 => x11_out_23,
   I4 => x11_out_25,
   I5 => W_61_7_i_11_n_0,
   O => W_61_7_i_7_n_0
);
W_61_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_61_7_i_4_n_0,
   I1 => W_61_7_i_12_n_0,
   I2 => x11_out_15,
   I3 => x11_out_22,
   I4 => x11_out_24,
   I5 => W_61_7_i_13_n_0,
   O => W_61_7_i_8_n_0
);
W_61_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_61_7_i_5_n_0,
   I1 => W_61_7_i_14_n_0,
   I2 => x11_out_14,
   I3 => x11_out_21,
   I4 => x11_out_23,
   I5 => W_61_7_i_15_n_0,
   O => W_61_7_i_9_n_0
);
W_62_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x50_out_10,
   I1 => x23_out_10,
   I2 => x47_out_28,
   I3 => x47_out_17,
   I4 => x47_out_13,
   O => W_62_11_i_10_n_0
);
W_62_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x23_out_9,
   I1 => x47_out_12,
   I2 => x47_out_16,
   I3 => x47_out_27,
   I4 => x50_out_9,
   O => W_62_11_i_11_n_0
);
W_62_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x50_out_9,
   I1 => x23_out_9,
   I2 => x47_out_27,
   I3 => x47_out_16,
   I4 => x47_out_12,
   O => W_62_11_i_12_n_0
);
W_62_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x23_out_8,
   I1 => x47_out_11,
   I2 => x47_out_15,
   I3 => x47_out_26,
   I4 => x50_out_8,
   O => W_62_11_i_13_n_0
);
W_62_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x50_out_8,
   I1 => x23_out_8,
   I2 => x47_out_26,
   I3 => x47_out_15,
   I4 => x47_out_11,
   O => W_62_11_i_14_n_0
);
W_62_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x23_out_7,
   I1 => x47_out_10,
   I2 => x47_out_14,
   I3 => x47_out_25,
   I4 => x50_out_7,
   O => W_62_11_i_15_n_0
);
W_62_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x50_out_7,
   I1 => x23_out_7,
   I2 => x47_out_25,
   I3 => x47_out_14,
   I4 => x47_out_10,
   O => W_62_11_i_16_n_0
);
W_62_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x23_out_6,
   I1 => x47_out_9,
   I2 => x47_out_13,
   I3 => x47_out_24,
   I4 => x50_out_6,
   O => W_62_11_i_17_n_0
);
W_62_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x8_out_20,
   I1 => x8_out_27,
   I2 => x8_out_29,
   I3 => W_62_11_i_10_n_0,
   I4 => W_62_11_i_11_n_0,
   O => W_62_11_i_2_n_0
);
W_62_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x8_out_19,
   I1 => x8_out_26,
   I2 => x8_out_28,
   I3 => W_62_11_i_12_n_0,
   I4 => W_62_11_i_13_n_0,
   O => W_62_11_i_3_n_0
);
W_62_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x8_out_18,
   I1 => x8_out_25,
   I2 => x8_out_27,
   I3 => W_62_11_i_14_n_0,
   I4 => W_62_11_i_15_n_0,
   O => W_62_11_i_4_n_0
);
W_62_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x8_out_17,
   I1 => x8_out_24,
   I2 => x8_out_26,
   I3 => W_62_11_i_16_n_0,
   I4 => W_62_11_i_17_n_0,
   O => W_62_11_i_5_n_0
);
W_62_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_62_11_i_2_n_0,
   I1 => W_62_15_i_16_n_0,
   I2 => x8_out_21,
   I3 => x8_out_28,
   I4 => x8_out_30,
   I5 => W_62_15_i_17_n_0,
   O => W_62_11_i_6_n_0
);
W_62_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_62_11_i_3_n_0,
   I1 => W_62_11_i_10_n_0,
   I2 => x8_out_20,
   I3 => x8_out_27,
   I4 => x8_out_29,
   I5 => W_62_11_i_11_n_0,
   O => W_62_11_i_7_n_0
);
W_62_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_62_11_i_4_n_0,
   I1 => W_62_11_i_12_n_0,
   I2 => x8_out_19,
   I3 => x8_out_26,
   I4 => x8_out_28,
   I5 => W_62_11_i_13_n_0,
   O => W_62_11_i_8_n_0
);
W_62_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_62_11_i_5_n_0,
   I1 => W_62_11_i_14_n_0,
   I2 => x8_out_18,
   I3 => x8_out_25,
   I4 => x8_out_27,
   I5 => W_62_11_i_15_n_0,
   O => W_62_11_i_9_n_0
);
W_62_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x50_out_14,
   I1 => x23_out_14,
   I2 => x47_out_0,
   I3 => x47_out_21,
   I4 => x47_out_17,
   O => W_62_15_i_10_n_0
);
W_62_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x23_out_13,
   I1 => x47_out_16,
   I2 => x47_out_20,
   I3 => x47_out_31,
   I4 => x50_out_13,
   O => W_62_15_i_11_n_0
);
W_62_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x50_out_13,
   I1 => x23_out_13,
   I2 => x47_out_31,
   I3 => x47_out_20,
   I4 => x47_out_16,
   O => W_62_15_i_12_n_0
);
W_62_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x23_out_12,
   I1 => x47_out_15,
   I2 => x47_out_19,
   I3 => x47_out_30,
   I4 => x50_out_12,
   O => W_62_15_i_13_n_0
);
W_62_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x50_out_12,
   I1 => x23_out_12,
   I2 => x47_out_30,
   I3 => x47_out_19,
   I4 => x47_out_15,
   O => W_62_15_i_14_n_0
);
W_62_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x23_out_11,
   I1 => x47_out_14,
   I2 => x47_out_18,
   I3 => x47_out_29,
   I4 => x50_out_11,
   O => W_62_15_i_15_n_0
);
W_62_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x50_out_11,
   I1 => x23_out_11,
   I2 => x47_out_29,
   I3 => x47_out_18,
   I4 => x47_out_14,
   O => W_62_15_i_16_n_0
);
W_62_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x23_out_10,
   I1 => x47_out_13,
   I2 => x47_out_17,
   I3 => x47_out_28,
   I4 => x50_out_10,
   O => W_62_15_i_17_n_0
);
W_62_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x8_out_24,
   I1 => x8_out_31,
   I2 => x8_out_1,
   I3 => W_62_15_i_10_n_0,
   I4 => W_62_15_i_11_n_0,
   O => W_62_15_i_2_n_0
);
W_62_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x8_out_23,
   I1 => x8_out_30,
   I2 => x8_out_0,
   I3 => W_62_15_i_12_n_0,
   I4 => W_62_15_i_13_n_0,
   O => W_62_15_i_3_n_0
);
W_62_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x8_out_22,
   I1 => x8_out_29,
   I2 => x8_out_31,
   I3 => W_62_15_i_14_n_0,
   I4 => W_62_15_i_15_n_0,
   O => W_62_15_i_4_n_0
);
W_62_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x8_out_21,
   I1 => x8_out_28,
   I2 => x8_out_30,
   I3 => W_62_15_i_16_n_0,
   I4 => W_62_15_i_17_n_0,
   O => W_62_15_i_5_n_0
);
W_62_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_62_15_i_2_n_0,
   I1 => W_62_19_i_16_n_0,
   I2 => x8_out_25,
   I3 => x8_out_0,
   I4 => x8_out_2,
   I5 => W_62_19_i_17_n_0,
   O => W_62_15_i_6_n_0
);
W_62_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_62_15_i_3_n_0,
   I1 => W_62_15_i_10_n_0,
   I2 => x8_out_24,
   I3 => x8_out_31,
   I4 => x8_out_1,
   I5 => W_62_15_i_11_n_0,
   O => W_62_15_i_7_n_0
);
W_62_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_62_15_i_4_n_0,
   I1 => W_62_15_i_12_n_0,
   I2 => x8_out_23,
   I3 => x8_out_30,
   I4 => x8_out_0,
   I5 => W_62_15_i_13_n_0,
   O => W_62_15_i_8_n_0
);
W_62_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_62_15_i_5_n_0,
   I1 => W_62_15_i_14_n_0,
   I2 => x8_out_22,
   I3 => x8_out_29,
   I4 => x8_out_31,
   I5 => W_62_15_i_15_n_0,
   O => W_62_15_i_9_n_0
);
W_62_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x50_out_18,
   I1 => x23_out_18,
   I2 => x47_out_4,
   I3 => x47_out_25,
   I4 => x47_out_21,
   O => W_62_19_i_10_n_0
);
W_62_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x23_out_17,
   I1 => x47_out_20,
   I2 => x47_out_24,
   I3 => x47_out_3,
   I4 => x50_out_17,
   O => W_62_19_i_11_n_0
);
W_62_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x50_out_17,
   I1 => x23_out_17,
   I2 => x47_out_3,
   I3 => x47_out_24,
   I4 => x47_out_20,
   O => W_62_19_i_12_n_0
);
W_62_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x23_out_16,
   I1 => x47_out_19,
   I2 => x47_out_23,
   I3 => x47_out_2,
   I4 => x50_out_16,
   O => W_62_19_i_13_n_0
);
W_62_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x50_out_16,
   I1 => x23_out_16,
   I2 => x47_out_2,
   I3 => x47_out_23,
   I4 => x47_out_19,
   O => W_62_19_i_14_n_0
);
W_62_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x23_out_15,
   I1 => x47_out_18,
   I2 => x47_out_22,
   I3 => x47_out_1,
   I4 => x50_out_15,
   O => W_62_19_i_15_n_0
);
W_62_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x50_out_15,
   I1 => x23_out_15,
   I2 => x47_out_1,
   I3 => x47_out_22,
   I4 => x47_out_18,
   O => W_62_19_i_16_n_0
);
W_62_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x23_out_14,
   I1 => x47_out_17,
   I2 => x47_out_21,
   I3 => x47_out_0,
   I4 => x50_out_14,
   O => W_62_19_i_17_n_0
);
W_62_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x8_out_28,
   I1 => x8_out_3,
   I2 => x8_out_5,
   I3 => W_62_19_i_10_n_0,
   I4 => W_62_19_i_11_n_0,
   O => W_62_19_i_2_n_0
);
W_62_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x8_out_27,
   I1 => x8_out_2,
   I2 => x8_out_4,
   I3 => W_62_19_i_12_n_0,
   I4 => W_62_19_i_13_n_0,
   O => W_62_19_i_3_n_0
);
W_62_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x8_out_26,
   I1 => x8_out_1,
   I2 => x8_out_3,
   I3 => W_62_19_i_14_n_0,
   I4 => W_62_19_i_15_n_0,
   O => W_62_19_i_4_n_0
);
W_62_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x8_out_25,
   I1 => x8_out_0,
   I2 => x8_out_2,
   I3 => W_62_19_i_16_n_0,
   I4 => W_62_19_i_17_n_0,
   O => W_62_19_i_5_n_0
);
W_62_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_62_19_i_2_n_0,
   I1 => W_62_23_i_16_n_0,
   I2 => x8_out_29,
   I3 => x8_out_4,
   I4 => x8_out_6,
   I5 => W_62_23_i_17_n_0,
   O => W_62_19_i_6_n_0
);
W_62_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_62_19_i_3_n_0,
   I1 => W_62_19_i_10_n_0,
   I2 => x8_out_28,
   I3 => x8_out_3,
   I4 => x8_out_5,
   I5 => W_62_19_i_11_n_0,
   O => W_62_19_i_7_n_0
);
W_62_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_62_19_i_4_n_0,
   I1 => W_62_19_i_12_n_0,
   I2 => x8_out_27,
   I3 => x8_out_2,
   I4 => x8_out_4,
   I5 => W_62_19_i_13_n_0,
   O => W_62_19_i_8_n_0
);
W_62_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_62_19_i_5_n_0,
   I1 => W_62_19_i_14_n_0,
   I2 => x8_out_26,
   I3 => x8_out_1,
   I4 => x8_out_3,
   I5 => W_62_19_i_15_n_0,
   O => W_62_19_i_9_n_0
);
W_62_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x50_out_22,
   I1 => x23_out_22,
   I2 => x47_out_8,
   I3 => x47_out_29,
   I4 => x47_out_25,
   O => W_62_23_i_10_n_0
);
W_62_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x23_out_21,
   I1 => x47_out_24,
   I2 => x47_out_28,
   I3 => x47_out_7,
   I4 => x50_out_21,
   O => W_62_23_i_11_n_0
);
W_62_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x50_out_21,
   I1 => x23_out_21,
   I2 => x47_out_7,
   I3 => x47_out_28,
   I4 => x47_out_24,
   O => W_62_23_i_12_n_0
);
W_62_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x23_out_20,
   I1 => x47_out_23,
   I2 => x47_out_27,
   I3 => x47_out_6,
   I4 => x50_out_20,
   O => W_62_23_i_13_n_0
);
W_62_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x50_out_20,
   I1 => x23_out_20,
   I2 => x47_out_6,
   I3 => x47_out_27,
   I4 => x47_out_23,
   O => W_62_23_i_14_n_0
);
W_62_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x23_out_19,
   I1 => x47_out_22,
   I2 => x47_out_26,
   I3 => x47_out_5,
   I4 => x50_out_19,
   O => W_62_23_i_15_n_0
);
W_62_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x50_out_19,
   I1 => x23_out_19,
   I2 => x47_out_5,
   I3 => x47_out_26,
   I4 => x47_out_22,
   O => W_62_23_i_16_n_0
);
W_62_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x23_out_18,
   I1 => x47_out_21,
   I2 => x47_out_25,
   I3 => x47_out_4,
   I4 => x50_out_18,
   O => W_62_23_i_17_n_0
);
W_62_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x8_out_7,
   I1 => x8_out_9,
   I2 => W_62_23_i_10_n_0,
   I3 => W_62_23_i_11_n_0,
   O => W_62_23_i_2_n_0
);
W_62_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x8_out_31,
   I1 => x8_out_6,
   I2 => x8_out_8,
   I3 => W_62_23_i_12_n_0,
   I4 => W_62_23_i_13_n_0,
   O => W_62_23_i_3_n_0
);
W_62_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x8_out_30,
   I1 => x8_out_5,
   I2 => x8_out_7,
   I3 => W_62_23_i_14_n_0,
   I4 => W_62_23_i_15_n_0,
   O => W_62_23_i_4_n_0
);
W_62_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x8_out_29,
   I1 => x8_out_4,
   I2 => x8_out_6,
   I3 => W_62_23_i_16_n_0,
   I4 => W_62_23_i_17_n_0,
   O => W_62_23_i_5_n_0
);
W_62_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x8_out_8,
   I1 => x8_out_10,
   I2 => W_62_27_i_16_n_0,
   I3 => W_62_27_i_17_n_0,
   I4 => W_62_23_i_2_n_0,
   O => W_62_23_i_6_n_0
);
W_62_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x8_out_7,
   I1 => x8_out_9,
   I2 => W_62_23_i_10_n_0,
   I3 => W_62_23_i_11_n_0,
   I4 => W_62_23_i_3_n_0,
   O => W_62_23_i_7_n_0
);
W_62_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_62_23_i_4_n_0,
   I1 => W_62_23_i_12_n_0,
   I2 => x8_out_31,
   I3 => x8_out_6,
   I4 => x8_out_8,
   I5 => W_62_23_i_13_n_0,
   O => W_62_23_i_8_n_0
);
W_62_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_62_23_i_5_n_0,
   I1 => W_62_23_i_14_n_0,
   I2 => x8_out_30,
   I3 => x8_out_5,
   I4 => x8_out_7,
   I5 => W_62_23_i_15_n_0,
   O => W_62_23_i_9_n_0
);
W_62_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x50_out_26,
   I1 => x23_out_26,
   I2 => x47_out_12,
   I3 => x47_out_1,
   I4 => x47_out_29,
   O => W_62_27_i_10_n_0
);
W_62_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x23_out_25,
   I1 => x47_out_28,
   I2 => x47_out_0,
   I3 => x47_out_11,
   I4 => x50_out_25,
   O => W_62_27_i_11_n_0
);
W_62_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x50_out_25,
   I1 => x23_out_25,
   I2 => x47_out_11,
   I3 => x47_out_0,
   I4 => x47_out_28,
   O => W_62_27_i_12_n_0
);
W_62_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x23_out_24,
   I1 => x47_out_27,
   I2 => x47_out_31,
   I3 => x47_out_10,
   I4 => x50_out_24,
   O => W_62_27_i_13_n_0
);
W_62_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x50_out_24,
   I1 => x23_out_24,
   I2 => x47_out_10,
   I3 => x47_out_31,
   I4 => x47_out_27,
   O => W_62_27_i_14_n_0
);
W_62_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x23_out_23,
   I1 => x47_out_26,
   I2 => x47_out_30,
   I3 => x47_out_9,
   I4 => x50_out_23,
   O => W_62_27_i_15_n_0
);
W_62_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x50_out_23,
   I1 => x23_out_23,
   I2 => x47_out_9,
   I3 => x47_out_30,
   I4 => x47_out_26,
   O => W_62_27_i_16_n_0
);
W_62_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x23_out_22,
   I1 => x47_out_25,
   I2 => x47_out_29,
   I3 => x47_out_8,
   I4 => x50_out_22,
   O => W_62_27_i_17_n_0
);
W_62_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x8_out_11,
   I1 => x8_out_13,
   I2 => W_62_27_i_10_n_0,
   I3 => W_62_27_i_11_n_0,
   O => W_62_27_i_2_n_0
);
W_62_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x8_out_10,
   I1 => x8_out_12,
   I2 => W_62_27_i_12_n_0,
   I3 => W_62_27_i_13_n_0,
   O => W_62_27_i_3_n_0
);
W_62_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x8_out_9,
   I1 => x8_out_11,
   I2 => W_62_27_i_14_n_0,
   I3 => W_62_27_i_15_n_0,
   O => W_62_27_i_4_n_0
);
W_62_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x8_out_8,
   I1 => x8_out_10,
   I2 => W_62_27_i_16_n_0,
   I3 => W_62_27_i_17_n_0,
   O => W_62_27_i_5_n_0
);
W_62_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x8_out_12,
   I1 => x8_out_14,
   I2 => W_62_31_i_13_n_0,
   I3 => W_62_31_i_14_n_0,
   I4 => W_62_27_i_2_n_0,
   O => W_62_27_i_6_n_0
);
W_62_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x8_out_11,
   I1 => x8_out_13,
   I2 => W_62_27_i_10_n_0,
   I3 => W_62_27_i_11_n_0,
   I4 => W_62_27_i_3_n_0,
   O => W_62_27_i_7_n_0
);
W_62_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x8_out_10,
   I1 => x8_out_12,
   I2 => W_62_27_i_12_n_0,
   I3 => W_62_27_i_13_n_0,
   I4 => W_62_27_i_4_n_0,
   O => W_62_27_i_8_n_0
);
W_62_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x8_out_9,
   I1 => x8_out_11,
   I2 => W_62_27_i_14_n_0,
   I3 => W_62_27_i_15_n_0,
   I4 => W_62_27_i_5_n_0,
   O => W_62_27_i_9_n_0
);
W_62_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x23_out_28,
   I1 => x47_out_31,
   I2 => x47_out_3,
   I3 => x47_out_14,
   I4 => x50_out_28,
   O => W_62_31_i_10_n_0
);
W_62_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x50_out_28,
   I1 => x23_out_28,
   I2 => x47_out_14,
   I3 => x47_out_3,
   I4 => x47_out_31,
   O => W_62_31_i_11_n_0
);
W_62_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x23_out_27,
   I1 => x47_out_30,
   I2 => x47_out_2,
   I3 => x47_out_13,
   I4 => x50_out_27,
   O => W_62_31_i_12_n_0
);
W_62_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x50_out_27,
   I1 => x23_out_27,
   I2 => x47_out_13,
   I3 => x47_out_2,
   I4 => x47_out_30,
   O => W_62_31_i_13_n_0
);
W_62_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x23_out_26,
   I1 => x47_out_29,
   I2 => x47_out_1,
   I3 => x47_out_12,
   I4 => x50_out_26,
   O => W_62_31_i_14_n_0
);
W_62_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x23_out_29,
   I1 => x47_out_4,
   I2 => x47_out_15,
   I3 => x50_out_29,
   O => W_62_31_i_15_n_0
);
W_62_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x8_out_17,
   I1 => x8_out_15,
   O => SIGMA_LCASE_119_out_0_30
);
W_62_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => x47_out_6,
   I1 => x47_out_17,
   I2 => x23_out_31,
   I3 => x50_out_31,
   I4 => x8_out_16,
   I5 => x8_out_18,
   O => W_62_31_i_17_n_0
);
W_62_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x47_out_16,
   I1 => x47_out_5,
   O => SIGMA_LCASE_015_out_30
);
W_62_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x50_out_30,
   I1 => x23_out_30,
   I2 => x47_out_16,
   I3 => x47_out_5,
   O => W_62_31_i_19_n_0
);
W_62_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x8_out_14,
   I1 => x8_out_16,
   I2 => W_62_31_i_9_n_0,
   I3 => W_62_31_i_10_n_0,
   O => W_62_31_i_2_n_0
);
W_62_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x8_out_13,
   I1 => x8_out_15,
   I2 => W_62_31_i_11_n_0,
   I3 => W_62_31_i_12_n_0,
   O => W_62_31_i_3_n_0
);
W_62_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x8_out_12,
   I1 => x8_out_14,
   I2 => W_62_31_i_13_n_0,
   I3 => W_62_31_i_14_n_0,
   O => W_62_31_i_4_n_0
);
W_62_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_62_31_i_15_n_0,
   I1 => SIGMA_LCASE_119_out_0_30,
   I2 => W_62_31_i_17_n_0,
   I3 => x23_out_30,
   I4 => SIGMA_LCASE_015_out_30,
   I5 => x50_out_30,
   O => W_62_31_i_5_n_0
);
W_62_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_62_31_i_2_n_0,
   I1 => W_62_31_i_19_n_0,
   I2 => x8_out_15,
   I3 => x8_out_17,
   I4 => W_62_31_i_15_n_0,
   O => W_62_31_i_6_n_0
);
W_62_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x8_out_14,
   I1 => x8_out_16,
   I2 => W_62_31_i_9_n_0,
   I3 => W_62_31_i_10_n_0,
   I4 => W_62_31_i_3_n_0,
   O => W_62_31_i_7_n_0
);
W_62_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x8_out_13,
   I1 => x8_out_15,
   I2 => W_62_31_i_11_n_0,
   I3 => W_62_31_i_12_n_0,
   I4 => W_62_31_i_4_n_0,
   O => W_62_31_i_8_n_0
);
W_62_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x50_out_29,
   I1 => x23_out_29,
   I2 => x47_out_15,
   I3 => x47_out_4,
   O => W_62_31_i_9_n_0
);
W_62_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x50_out_2,
   I1 => x23_out_2,
   I2 => x47_out_20,
   I3 => x47_out_9,
   I4 => x47_out_5,
   O => W_62_3_i_10_n_0
);
W_62_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x23_out_1,
   I1 => x47_out_4,
   I2 => x47_out_8,
   I3 => x47_out_19,
   I4 => x50_out_1,
   O => W_62_3_i_11_n_0
);
W_62_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x47_out_19,
   I1 => x47_out_8,
   I2 => x47_out_4,
   O => SIGMA_LCASE_015_out_1
);
W_62_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x8_out_21,
   I1 => x8_out_19,
   I2 => x8_out_12,
   O => SIGMA_LCASE_119_out_0_2
);
W_62_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x8_out_20,
   I1 => x8_out_18,
   I2 => x8_out_11,
   O => SIGMA_LCASE_119_out_1
);
W_62_3_i_15 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x50_out_1,
   I1 => x23_out_1,
   I2 => x47_out_19,
   I3 => x47_out_8,
   I4 => x47_out_4,
   O => W_62_3_i_15_n_0
);
W_62_3_i_16 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x47_out_18,
   I1 => x47_out_7,
   I2 => x47_out_3,
   O => SIGMA_LCASE_015_out_0
);
W_62_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x8_out_12,
   I1 => x8_out_19,
   I2 => x8_out_21,
   I3 => W_62_3_i_10_n_0,
   I4 => W_62_3_i_11_n_0,
   O => W_62_3_i_2_n_0
);
W_62_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_62_3_i_11_n_0,
   I1 => x8_out_21,
   I2 => x8_out_19,
   I3 => x8_out_12,
   I4 => W_62_3_i_10_n_0,
   O => W_62_3_i_3_n_0
);
W_62_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_015_out_1,
   I1 => x23_out_1,
   I2 => x50_out_1,
   I3 => x8_out_11,
   I4 => x8_out_18,
   I5 => x8_out_20,
   O => W_62_3_i_4_n_0
);
W_62_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x50_out_0,
   I1 => x23_out_0,
   I2 => x47_out_18,
   I3 => x47_out_7,
   I4 => x47_out_3,
   O => W_62_3_i_5_n_0
);
W_62_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_62_3_i_2_n_0,
   I1 => W_62_7_i_16_n_0,
   I2 => x8_out_13,
   I3 => x8_out_20,
   I4 => x8_out_22,
   I5 => W_62_7_i_17_n_0,
   O => W_62_3_i_6_n_0
);
W_62_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_62_3_i_10_n_0,
   I1 => SIGMA_LCASE_119_out_0_2,
   I2 => x50_out_1,
   I3 => x23_out_1,
   I4 => SIGMA_LCASE_015_out_1,
   I5 => SIGMA_LCASE_119_out_1,
   O => W_62_3_i_7_n_0
);
W_62_3_i_8 : LUT5
  generic map(
   INIT => X"99969666"
  )
 port map (
   I0 => SIGMA_LCASE_119_out_1,
   I1 => W_62_3_i_15_n_0,
   I2 => x50_out_0,
   I3 => SIGMA_LCASE_015_out_0,
   I4 => x23_out_0,
   O => W_62_3_i_8_n_0
);
W_62_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_62_3_i_5_n_0,
   I1 => x8_out_10,
   I2 => x8_out_17,
   I3 => x8_out_19,
   O => W_62_3_i_9_n_0
);
W_62_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x50_out_6,
   I1 => x23_out_6,
   I2 => x47_out_24,
   I3 => x47_out_13,
   I4 => x47_out_9,
   O => W_62_7_i_10_n_0
);
W_62_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x23_out_5,
   I1 => x47_out_8,
   I2 => x47_out_12,
   I3 => x47_out_23,
   I4 => x50_out_5,
   O => W_62_7_i_11_n_0
);
W_62_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x50_out_5,
   I1 => x23_out_5,
   I2 => x47_out_23,
   I3 => x47_out_12,
   I4 => x47_out_8,
   O => W_62_7_i_12_n_0
);
W_62_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x23_out_4,
   I1 => x47_out_7,
   I2 => x47_out_11,
   I3 => x47_out_22,
   I4 => x50_out_4,
   O => W_62_7_i_13_n_0
);
W_62_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x50_out_4,
   I1 => x23_out_4,
   I2 => x47_out_22,
   I3 => x47_out_11,
   I4 => x47_out_7,
   O => W_62_7_i_14_n_0
);
W_62_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x23_out_3,
   I1 => x47_out_6,
   I2 => x47_out_10,
   I3 => x47_out_21,
   I4 => x50_out_3,
   O => W_62_7_i_15_n_0
);
W_62_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x50_out_3,
   I1 => x23_out_3,
   I2 => x47_out_21,
   I3 => x47_out_10,
   I4 => x47_out_6,
   O => W_62_7_i_16_n_0
);
W_62_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x23_out_2,
   I1 => x47_out_5,
   I2 => x47_out_9,
   I3 => x47_out_20,
   I4 => x50_out_2,
   O => W_62_7_i_17_n_0
);
W_62_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x8_out_16,
   I1 => x8_out_23,
   I2 => x8_out_25,
   I3 => W_62_7_i_10_n_0,
   I4 => W_62_7_i_11_n_0,
   O => W_62_7_i_2_n_0
);
W_62_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x8_out_15,
   I1 => x8_out_22,
   I2 => x8_out_24,
   I3 => W_62_7_i_12_n_0,
   I4 => W_62_7_i_13_n_0,
   O => W_62_7_i_3_n_0
);
W_62_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x8_out_14,
   I1 => x8_out_21,
   I2 => x8_out_23,
   I3 => W_62_7_i_14_n_0,
   I4 => W_62_7_i_15_n_0,
   O => W_62_7_i_4_n_0
);
W_62_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x8_out_13,
   I1 => x8_out_20,
   I2 => x8_out_22,
   I3 => W_62_7_i_16_n_0,
   I4 => W_62_7_i_17_n_0,
   O => W_62_7_i_5_n_0
);
W_62_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_62_7_i_2_n_0,
   I1 => W_62_11_i_16_n_0,
   I2 => x8_out_17,
   I3 => x8_out_24,
   I4 => x8_out_26,
   I5 => W_62_11_i_17_n_0,
   O => W_62_7_i_6_n_0
);
W_62_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_62_7_i_3_n_0,
   I1 => W_62_7_i_10_n_0,
   I2 => x8_out_16,
   I3 => x8_out_23,
   I4 => x8_out_25,
   I5 => W_62_7_i_11_n_0,
   O => W_62_7_i_7_n_0
);
W_62_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_62_7_i_4_n_0,
   I1 => W_62_7_i_12_n_0,
   I2 => x8_out_15,
   I3 => x8_out_22,
   I4 => x8_out_24,
   I5 => W_62_7_i_13_n_0,
   O => W_62_7_i_8_n_0
);
W_62_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_62_7_i_5_n_0,
   I1 => W_62_7_i_14_n_0,
   I2 => x8_out_14,
   I3 => x8_out_21,
   I4 => x8_out_23,
   I5 => W_62_7_i_15_n_0,
   O => W_62_7_i_9_n_0
);
W_63_11_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x47_out_10,
   I1 => x20_out_10,
   I2 => x44_out_28,
   I3 => x44_out_17,
   I4 => x44_out_13,
   O => W_63_11_i_10_n_0
);
W_63_11_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x20_out_9,
   I1 => x44_out_12,
   I2 => x44_out_16,
   I3 => x44_out_27,
   I4 => x47_out_9,
   O => W_63_11_i_11_n_0
);
W_63_11_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x47_out_9,
   I1 => x20_out_9,
   I2 => x44_out_27,
   I3 => x44_out_16,
   I4 => x44_out_12,
   O => W_63_11_i_12_n_0
);
W_63_11_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x20_out_8,
   I1 => x44_out_11,
   I2 => x44_out_15,
   I3 => x44_out_26,
   I4 => x47_out_8,
   O => W_63_11_i_13_n_0
);
W_63_11_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x47_out_8,
   I1 => x20_out_8,
   I2 => x44_out_26,
   I3 => x44_out_15,
   I4 => x44_out_11,
   O => W_63_11_i_14_n_0
);
W_63_11_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x20_out_7,
   I1 => x44_out_10,
   I2 => x44_out_14,
   I3 => x44_out_25,
   I4 => x47_out_7,
   O => W_63_11_i_15_n_0
);
W_63_11_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x47_out_7,
   I1 => x20_out_7,
   I2 => x44_out_25,
   I3 => x44_out_14,
   I4 => x44_out_10,
   O => W_63_11_i_16_n_0
);
W_63_11_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x20_out_6,
   I1 => x44_out_9,
   I2 => x44_out_13,
   I3 => x44_out_24,
   I4 => x47_out_6,
   O => W_63_11_i_17_n_0
);
W_63_11_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x_20,
   I1 => x_27,
   I2 => x_29,
   I3 => W_63_11_i_10_n_0,
   I4 => W_63_11_i_11_n_0,
   O => W_63_11_i_2_n_0
);
W_63_11_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x_19,
   I1 => x_26,
   I2 => x_28,
   I3 => W_63_11_i_12_n_0,
   I4 => W_63_11_i_13_n_0,
   O => W_63_11_i_3_n_0
);
W_63_11_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x_18,
   I1 => x_25,
   I2 => x_27,
   I3 => W_63_11_i_14_n_0,
   I4 => W_63_11_i_15_n_0,
   O => W_63_11_i_4_n_0
);
W_63_11_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x_17,
   I1 => x_24,
   I2 => x_26,
   I3 => W_63_11_i_16_n_0,
   I4 => W_63_11_i_17_n_0,
   O => W_63_11_i_5_n_0
);
W_63_11_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_63_11_i_2_n_0,
   I1 => W_63_15_i_16_n_0,
   I2 => x_21,
   I3 => x_28,
   I4 => x_30,
   I5 => W_63_15_i_17_n_0,
   O => W_63_11_i_6_n_0
);
W_63_11_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_63_11_i_3_n_0,
   I1 => W_63_11_i_10_n_0,
   I2 => x_20,
   I3 => x_27,
   I4 => x_29,
   I5 => W_63_11_i_11_n_0,
   O => W_63_11_i_7_n_0
);
W_63_11_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_63_11_i_4_n_0,
   I1 => W_63_11_i_12_n_0,
   I2 => x_19,
   I3 => x_26,
   I4 => x_28,
   I5 => W_63_11_i_13_n_0,
   O => W_63_11_i_8_n_0
);
W_63_11_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_63_11_i_5_n_0,
   I1 => W_63_11_i_14_n_0,
   I2 => x_18,
   I3 => x_25,
   I4 => x_27,
   I5 => W_63_11_i_15_n_0,
   O => W_63_11_i_9_n_0
);
W_63_15_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x47_out_14,
   I1 => x20_out_14,
   I2 => x44_out_0,
   I3 => x44_out_21,
   I4 => x44_out_17,
   O => W_63_15_i_10_n_0
);
W_63_15_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x20_out_13,
   I1 => x44_out_16,
   I2 => x44_out_20,
   I3 => x44_out_31,
   I4 => x47_out_13,
   O => W_63_15_i_11_n_0
);
W_63_15_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x47_out_13,
   I1 => x20_out_13,
   I2 => x44_out_31,
   I3 => x44_out_20,
   I4 => x44_out_16,
   O => W_63_15_i_12_n_0
);
W_63_15_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x20_out_12,
   I1 => x44_out_15,
   I2 => x44_out_19,
   I3 => x44_out_30,
   I4 => x47_out_12,
   O => W_63_15_i_13_n_0
);
W_63_15_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x47_out_12,
   I1 => x20_out_12,
   I2 => x44_out_30,
   I3 => x44_out_19,
   I4 => x44_out_15,
   O => W_63_15_i_14_n_0
);
W_63_15_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x20_out_11,
   I1 => x44_out_14,
   I2 => x44_out_18,
   I3 => x44_out_29,
   I4 => x47_out_11,
   O => W_63_15_i_15_n_0
);
W_63_15_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x47_out_11,
   I1 => x20_out_11,
   I2 => x44_out_29,
   I3 => x44_out_18,
   I4 => x44_out_14,
   O => W_63_15_i_16_n_0
);
W_63_15_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x20_out_10,
   I1 => x44_out_13,
   I2 => x44_out_17,
   I3 => x44_out_28,
   I4 => x47_out_10,
   O => W_63_15_i_17_n_0
);
W_63_15_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x_24,
   I1 => x_31,
   I2 => x_1,
   I3 => W_63_15_i_10_n_0,
   I4 => W_63_15_i_11_n_0,
   O => W_63_15_i_2_n_0
);
W_63_15_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x_23,
   I1 => x_30,
   I2 => x_0,
   I3 => W_63_15_i_12_n_0,
   I4 => W_63_15_i_13_n_0,
   O => W_63_15_i_3_n_0
);
W_63_15_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x_22,
   I1 => x_29,
   I2 => x_31,
   I3 => W_63_15_i_14_n_0,
   I4 => W_63_15_i_15_n_0,
   O => W_63_15_i_4_n_0
);
W_63_15_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x_21,
   I1 => x_28,
   I2 => x_30,
   I3 => W_63_15_i_16_n_0,
   I4 => W_63_15_i_17_n_0,
   O => W_63_15_i_5_n_0
);
W_63_15_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_63_15_i_2_n_0,
   I1 => W_63_19_i_16_n_0,
   I2 => x_25,
   I3 => x_0,
   I4 => x_2,
   I5 => W_63_19_i_17_n_0,
   O => W_63_15_i_6_n_0
);
W_63_15_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_63_15_i_3_n_0,
   I1 => W_63_15_i_10_n_0,
   I2 => x_24,
   I3 => x_31,
   I4 => x_1,
   I5 => W_63_15_i_11_n_0,
   O => W_63_15_i_7_n_0
);
W_63_15_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_63_15_i_4_n_0,
   I1 => W_63_15_i_12_n_0,
   I2 => x_23,
   I3 => x_30,
   I4 => x_0,
   I5 => W_63_15_i_13_n_0,
   O => W_63_15_i_8_n_0
);
W_63_15_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_63_15_i_5_n_0,
   I1 => W_63_15_i_14_n_0,
   I2 => x_22,
   I3 => x_29,
   I4 => x_31,
   I5 => W_63_15_i_15_n_0,
   O => W_63_15_i_9_n_0
);
W_63_19_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x47_out_18,
   I1 => x20_out_18,
   I2 => x44_out_4,
   I3 => x44_out_25,
   I4 => x44_out_21,
   O => W_63_19_i_10_n_0
);
W_63_19_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x20_out_17,
   I1 => x44_out_20,
   I2 => x44_out_24,
   I3 => x44_out_3,
   I4 => x47_out_17,
   O => W_63_19_i_11_n_0
);
W_63_19_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x47_out_17,
   I1 => x20_out_17,
   I2 => x44_out_3,
   I3 => x44_out_24,
   I4 => x44_out_20,
   O => W_63_19_i_12_n_0
);
W_63_19_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x20_out_16,
   I1 => x44_out_19,
   I2 => x44_out_23,
   I3 => x44_out_2,
   I4 => x47_out_16,
   O => W_63_19_i_13_n_0
);
W_63_19_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x47_out_16,
   I1 => x20_out_16,
   I2 => x44_out_2,
   I3 => x44_out_23,
   I4 => x44_out_19,
   O => W_63_19_i_14_n_0
);
W_63_19_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x20_out_15,
   I1 => x44_out_18,
   I2 => x44_out_22,
   I3 => x44_out_1,
   I4 => x47_out_15,
   O => W_63_19_i_15_n_0
);
W_63_19_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x47_out_15,
   I1 => x20_out_15,
   I2 => x44_out_1,
   I3 => x44_out_22,
   I4 => x44_out_18,
   O => W_63_19_i_16_n_0
);
W_63_19_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x20_out_14,
   I1 => x44_out_17,
   I2 => x44_out_21,
   I3 => x44_out_0,
   I4 => x47_out_14,
   O => W_63_19_i_17_n_0
);
W_63_19_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x_28,
   I1 => x_3,
   I2 => x_5,
   I3 => W_63_19_i_10_n_0,
   I4 => W_63_19_i_11_n_0,
   O => W_63_19_i_2_n_0
);
W_63_19_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x_27,
   I1 => x_2,
   I2 => x_4,
   I3 => W_63_19_i_12_n_0,
   I4 => W_63_19_i_13_n_0,
   O => W_63_19_i_3_n_0
);
W_63_19_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x_26,
   I1 => x_1,
   I2 => x_3,
   I3 => W_63_19_i_14_n_0,
   I4 => W_63_19_i_15_n_0,
   O => W_63_19_i_4_n_0
);
W_63_19_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x_25,
   I1 => x_0,
   I2 => x_2,
   I3 => W_63_19_i_16_n_0,
   I4 => W_63_19_i_17_n_0,
   O => W_63_19_i_5_n_0
);
W_63_19_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_63_19_i_2_n_0,
   I1 => W_63_23_i_16_n_0,
   I2 => x_29,
   I3 => x_4,
   I4 => x_6,
   I5 => W_63_23_i_17_n_0,
   O => W_63_19_i_6_n_0
);
W_63_19_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_63_19_i_3_n_0,
   I1 => W_63_19_i_10_n_0,
   I2 => x_28,
   I3 => x_3,
   I4 => x_5,
   I5 => W_63_19_i_11_n_0,
   O => W_63_19_i_7_n_0
);
W_63_19_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_63_19_i_4_n_0,
   I1 => W_63_19_i_12_n_0,
   I2 => x_27,
   I3 => x_2,
   I4 => x_4,
   I5 => W_63_19_i_13_n_0,
   O => W_63_19_i_8_n_0
);
W_63_19_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_63_19_i_5_n_0,
   I1 => W_63_19_i_14_n_0,
   I2 => x_26,
   I3 => x_1,
   I4 => x_3,
   I5 => W_63_19_i_15_n_0,
   O => W_63_19_i_9_n_0
);
W_63_23_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x47_out_22,
   I1 => x20_out_22,
   I2 => x44_out_8,
   I3 => x44_out_29,
   I4 => x44_out_25,
   O => W_63_23_i_10_n_0
);
W_63_23_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x20_out_21,
   I1 => x44_out_24,
   I2 => x44_out_28,
   I3 => x44_out_7,
   I4 => x47_out_21,
   O => W_63_23_i_11_n_0
);
W_63_23_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x47_out_21,
   I1 => x20_out_21,
   I2 => x44_out_7,
   I3 => x44_out_28,
   I4 => x44_out_24,
   O => W_63_23_i_12_n_0
);
W_63_23_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x20_out_20,
   I1 => x44_out_23,
   I2 => x44_out_27,
   I3 => x44_out_6,
   I4 => x47_out_20,
   O => W_63_23_i_13_n_0
);
W_63_23_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x47_out_20,
   I1 => x20_out_20,
   I2 => x44_out_6,
   I3 => x44_out_27,
   I4 => x44_out_23,
   O => W_63_23_i_14_n_0
);
W_63_23_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x20_out_19,
   I1 => x44_out_22,
   I2 => x44_out_26,
   I3 => x44_out_5,
   I4 => x47_out_19,
   O => W_63_23_i_15_n_0
);
W_63_23_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x47_out_19,
   I1 => x20_out_19,
   I2 => x44_out_5,
   I3 => x44_out_26,
   I4 => x44_out_22,
   O => W_63_23_i_16_n_0
);
W_63_23_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x20_out_18,
   I1 => x44_out_21,
   I2 => x44_out_25,
   I3 => x44_out_4,
   I4 => x47_out_18,
   O => W_63_23_i_17_n_0
);
W_63_23_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x_7,
   I1 => x_9,
   I2 => W_63_23_i_10_n_0,
   I3 => W_63_23_i_11_n_0,
   O => W_63_23_i_2_n_0
);
W_63_23_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x_31,
   I1 => x_6,
   I2 => x_8,
   I3 => W_63_23_i_12_n_0,
   I4 => W_63_23_i_13_n_0,
   O => W_63_23_i_3_n_0
);
W_63_23_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x_30,
   I1 => x_5,
   I2 => x_7,
   I3 => W_63_23_i_14_n_0,
   I4 => W_63_23_i_15_n_0,
   O => W_63_23_i_4_n_0
);
W_63_23_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x_29,
   I1 => x_4,
   I2 => x_6,
   I3 => W_63_23_i_16_n_0,
   I4 => W_63_23_i_17_n_0,
   O => W_63_23_i_5_n_0
);
W_63_23_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x_8,
   I1 => x_10,
   I2 => W_63_27_i_16_n_0,
   I3 => W_63_27_i_17_n_0,
   I4 => W_63_23_i_2_n_0,
   O => W_63_23_i_6_n_0
);
W_63_23_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x_7,
   I1 => x_9,
   I2 => W_63_23_i_10_n_0,
   I3 => W_63_23_i_11_n_0,
   I4 => W_63_23_i_3_n_0,
   O => W_63_23_i_7_n_0
);
W_63_23_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_63_23_i_4_n_0,
   I1 => W_63_23_i_12_n_0,
   I2 => x_31,
   I3 => x_6,
   I4 => x_8,
   I5 => W_63_23_i_13_n_0,
   O => W_63_23_i_8_n_0
);
W_63_23_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_63_23_i_5_n_0,
   I1 => W_63_23_i_14_n_0,
   I2 => x_30,
   I3 => x_5,
   I4 => x_7,
   I5 => W_63_23_i_15_n_0,
   O => W_63_23_i_9_n_0
);
W_63_27_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x47_out_26,
   I1 => x20_out_26,
   I2 => x44_out_12,
   I3 => x44_out_1,
   I4 => x44_out_29,
   O => W_63_27_i_10_n_0
);
W_63_27_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x20_out_25,
   I1 => x44_out_28,
   I2 => x44_out_0,
   I3 => x44_out_11,
   I4 => x47_out_25,
   O => W_63_27_i_11_n_0
);
W_63_27_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x47_out_25,
   I1 => x20_out_25,
   I2 => x44_out_11,
   I3 => x44_out_0,
   I4 => x44_out_28,
   O => W_63_27_i_12_n_0
);
W_63_27_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x20_out_24,
   I1 => x44_out_27,
   I2 => x44_out_31,
   I3 => x44_out_10,
   I4 => x47_out_24,
   O => W_63_27_i_13_n_0
);
W_63_27_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x47_out_24,
   I1 => x20_out_24,
   I2 => x44_out_10,
   I3 => x44_out_31,
   I4 => x44_out_27,
   O => W_63_27_i_14_n_0
);
W_63_27_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x20_out_23,
   I1 => x44_out_26,
   I2 => x44_out_30,
   I3 => x44_out_9,
   I4 => x47_out_23,
   O => W_63_27_i_15_n_0
);
W_63_27_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x47_out_23,
   I1 => x20_out_23,
   I2 => x44_out_9,
   I3 => x44_out_30,
   I4 => x44_out_26,
   O => W_63_27_i_16_n_0
);
W_63_27_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x20_out_22,
   I1 => x44_out_25,
   I2 => x44_out_29,
   I3 => x44_out_8,
   I4 => x47_out_22,
   O => W_63_27_i_17_n_0
);
W_63_27_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x_11,
   I1 => x_13,
   I2 => W_63_27_i_10_n_0,
   I3 => W_63_27_i_11_n_0,
   O => W_63_27_i_2_n_0
);
W_63_27_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x_10,
   I1 => x_12,
   I2 => W_63_27_i_12_n_0,
   I3 => W_63_27_i_13_n_0,
   O => W_63_27_i_3_n_0
);
W_63_27_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x_9,
   I1 => x_11,
   I2 => W_63_27_i_14_n_0,
   I3 => W_63_27_i_15_n_0,
   O => W_63_27_i_4_n_0
);
W_63_27_i_5 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x_8,
   I1 => x_10,
   I2 => W_63_27_i_16_n_0,
   I3 => W_63_27_i_17_n_0,
   O => W_63_27_i_5_n_0
);
W_63_27_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x_12,
   I1 => x_14,
   I2 => W_63_31_i_13_n_0,
   I3 => W_63_31_i_14_n_0,
   I4 => W_63_27_i_2_n_0,
   O => W_63_27_i_6_n_0
);
W_63_27_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x_11,
   I1 => x_13,
   I2 => W_63_27_i_10_n_0,
   I3 => W_63_27_i_11_n_0,
   I4 => W_63_27_i_3_n_0,
   O => W_63_27_i_7_n_0
);
W_63_27_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x_10,
   I1 => x_12,
   I2 => W_63_27_i_12_n_0,
   I3 => W_63_27_i_13_n_0,
   I4 => W_63_27_i_4_n_0,
   O => W_63_27_i_8_n_0
);
W_63_27_i_9 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x_9,
   I1 => x_11,
   I2 => W_63_27_i_14_n_0,
   I3 => W_63_27_i_15_n_0,
   I4 => W_63_27_i_5_n_0,
   O => W_63_27_i_9_n_0
);
W_63_31_i_10 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x20_out_28,
   I1 => x44_out_31,
   I2 => x44_out_3,
   I3 => x44_out_14,
   I4 => x47_out_28,
   O => W_63_31_i_10_n_0
);
W_63_31_i_11 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x47_out_28,
   I1 => x20_out_28,
   I2 => x44_out_14,
   I3 => x44_out_3,
   I4 => x44_out_31,
   O => W_63_31_i_11_n_0
);
W_63_31_i_12 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x20_out_27,
   I1 => x44_out_30,
   I2 => x44_out_2,
   I3 => x44_out_13,
   I4 => x47_out_27,
   O => W_63_31_i_12_n_0
);
W_63_31_i_13 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x47_out_27,
   I1 => x20_out_27,
   I2 => x44_out_13,
   I3 => x44_out_2,
   I4 => x44_out_30,
   O => W_63_31_i_13_n_0
);
W_63_31_i_14 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x20_out_26,
   I1 => x44_out_29,
   I2 => x44_out_1,
   I3 => x44_out_12,
   I4 => x47_out_26,
   O => W_63_31_i_14_n_0
);
W_63_31_i_15 : LUT4
  generic map(
   INIT => X"be28"
  )
 port map (
   I0 => x20_out_29,
   I1 => x44_out_4,
   I2 => x44_out_15,
   I3 => x47_out_29,
   O => W_63_31_i_15_n_0
);
W_63_31_i_16 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x_17,
   I1 => x_15,
   O => SIGMA_LCASE_1_0_30
);
W_63_31_i_17 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => x44_out_6,
   I1 => x44_out_17,
   I2 => x20_out_31,
   I3 => x47_out_31,
   I4 => x_16,
   I5 => x_18,
   O => W_63_31_i_17_n_0
);
W_63_31_i_18 : LUT2
  generic map(
   INIT => X"6"
  )
 port map (
   I0 => x44_out_16,
   I1 => x44_out_5,
   O => SIGMA_LCASE_0_30
);
W_63_31_i_19 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x47_out_30,
   I1 => x20_out_30,
   I2 => x44_out_16,
   I3 => x44_out_5,
   O => W_63_31_i_19_n_0
);
W_63_31_i_2 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x_14,
   I1 => x_16,
   I2 => W_63_31_i_9_n_0,
   I3 => W_63_31_i_10_n_0,
   O => W_63_31_i_2_n_0
);
W_63_31_i_3 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x_13,
   I1 => x_15,
   I2 => W_63_31_i_11_n_0,
   I3 => W_63_31_i_12_n_0,
   O => W_63_31_i_3_n_0
);
W_63_31_i_4 : LUT4
  generic map(
   INIT => X"f660"
  )
 port map (
   I0 => x_12,
   I1 => x_14,
   I2 => W_63_31_i_13_n_0,
   I3 => W_63_31_i_14_n_0,
   O => W_63_31_i_4_n_0
);
W_63_31_i_5 : LUT6
  generic map(
   INIT => X"e187871e871e1e78"
  )
 port map (
   I0 => W_63_31_i_15_n_0,
   I1 => SIGMA_LCASE_1_0_30,
   I2 => W_63_31_i_17_n_0,
   I3 => x20_out_30,
   I4 => SIGMA_LCASE_0_30,
   I5 => x47_out_30,
   O => W_63_31_i_5_n_0
);
W_63_31_i_6 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_63_31_i_2_n_0,
   I1 => W_63_31_i_19_n_0,
   I2 => x_15,
   I3 => x_17,
   I4 => W_63_31_i_15_n_0,
   O => W_63_31_i_6_n_0
);
W_63_31_i_7 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x_14,
   I1 => x_16,
   I2 => W_63_31_i_9_n_0,
   I3 => W_63_31_i_10_n_0,
   I4 => W_63_31_i_3_n_0,
   O => W_63_31_i_7_n_0
);
W_63_31_i_8 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x_13,
   I1 => x_15,
   I2 => W_63_31_i_11_n_0,
   I3 => W_63_31_i_12_n_0,
   I4 => W_63_31_i_4_n_0,
   O => W_63_31_i_8_n_0
);
W_63_31_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => x47_out_29,
   I1 => x20_out_29,
   I2 => x44_out_15,
   I3 => x44_out_4,
   O => W_63_31_i_9_n_0
);
W_63_3_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x47_out_2,
   I1 => x20_out_2,
   I2 => x44_out_20,
   I3 => x44_out_9,
   I4 => x44_out_5,
   O => W_63_3_i_10_n_0
);
W_63_3_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x20_out_1,
   I1 => x44_out_4,
   I2 => x44_out_8,
   I3 => x44_out_19,
   I4 => x47_out_1,
   O => W_63_3_i_11_n_0
);
W_63_3_i_12 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x44_out_19,
   I1 => x44_out_8,
   I2 => x44_out_4,
   O => SIGMA_LCASE_0_1
);
W_63_3_i_13 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x_21,
   I1 => x_19,
   I2 => x_12,
   O => SIGMA_LCASE_1_0_2
);
W_63_3_i_14 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x_20,
   I1 => x_18,
   I2 => x_11,
   O => SIGMA_LCASE_1_1
);
W_63_3_i_15 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x47_out_1,
   I1 => x20_out_1,
   I2 => x44_out_19,
   I3 => x44_out_8,
   I4 => x44_out_4,
   O => W_63_3_i_15_n_0
);
W_63_3_i_16 : LUT3
  generic map(
   INIT => X"96"
  )
 port map (
   I0 => x44_out_18,
   I1 => x44_out_7,
   I2 => x44_out_3,
   O => SIGMA_LCASE_0_0
);
W_63_3_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x_12,
   I1 => x_19,
   I2 => x_21,
   I3 => W_63_3_i_10_n_0,
   I4 => W_63_3_i_11_n_0,
   O => W_63_3_i_2_n_0
);
W_63_3_i_3 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => W_63_3_i_11_n_0,
   I1 => x_21,
   I2 => x_19,
   I3 => x_12,
   I4 => W_63_3_i_10_n_0,
   O => W_63_3_i_3_n_0
);
W_63_3_i_4 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => SIGMA_LCASE_0_1,
   I1 => x20_out_1,
   I2 => x47_out_1,
   I3 => x_11,
   I4 => x_18,
   I5 => x_20,
   O => W_63_3_i_4_n_0
);
W_63_3_i_5 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x47_out_0,
   I1 => x20_out_0,
   I2 => x44_out_18,
   I3 => x44_out_7,
   I4 => x44_out_3,
   O => W_63_3_i_5_n_0
);
W_63_3_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_63_3_i_2_n_0,
   I1 => W_63_7_i_16_n_0,
   I2 => x_13,
   I3 => x_20,
   I4 => x_22,
   I5 => W_63_7_i_17_n_0,
   O => W_63_3_i_6_n_0
);
W_63_3_i_7 : LUT6
  generic map(
   INIT => X"6999999699969666"
  )
 port map (
   I0 => W_63_3_i_10_n_0,
   I1 => SIGMA_LCASE_1_0_2,
   I2 => x47_out_1,
   I3 => x20_out_1,
   I4 => SIGMA_LCASE_0_1,
   I5 => SIGMA_LCASE_1_1,
   O => W_63_3_i_7_n_0
);
W_63_3_i_8 : LUT5
  generic map(
   INIT => X"99969666"
  )
 port map (
   I0 => SIGMA_LCASE_1_1,
   I1 => W_63_3_i_15_n_0,
   I2 => x47_out_0,
   I3 => SIGMA_LCASE_0_0,
   I4 => x20_out_0,
   O => W_63_3_i_8_n_0
);
W_63_3_i_9 : LUT4
  generic map(
   INIT => X"6996"
  )
 port map (
   I0 => W_63_3_i_5_n_0,
   I1 => x_10,
   I2 => x_17,
   I3 => x_19,
   O => W_63_3_i_9_n_0
);
W_63_7_i_10 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x47_out_6,
   I1 => x20_out_6,
   I2 => x44_out_24,
   I3 => x44_out_13,
   I4 => x44_out_9,
   O => W_63_7_i_10_n_0
);
W_63_7_i_11 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x20_out_5,
   I1 => x44_out_8,
   I2 => x44_out_12,
   I3 => x44_out_23,
   I4 => x47_out_5,
   O => W_63_7_i_11_n_0
);
W_63_7_i_12 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x47_out_5,
   I1 => x20_out_5,
   I2 => x44_out_23,
   I3 => x44_out_12,
   I4 => x44_out_8,
   O => W_63_7_i_12_n_0
);
W_63_7_i_13 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x20_out_4,
   I1 => x44_out_7,
   I2 => x44_out_11,
   I3 => x44_out_22,
   I4 => x47_out_4,
   O => W_63_7_i_13_n_0
);
W_63_7_i_14 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x47_out_4,
   I1 => x20_out_4,
   I2 => x44_out_22,
   I3 => x44_out_11,
   I4 => x44_out_7,
   O => W_63_7_i_14_n_0
);
W_63_7_i_15 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x20_out_3,
   I1 => x44_out_6,
   I2 => x44_out_10,
   I3 => x44_out_21,
   I4 => x47_out_3,
   O => W_63_7_i_15_n_0
);
W_63_7_i_16 : LUT5
  generic map(
   INIT => X"96696996"
  )
 port map (
   I0 => x47_out_3,
   I1 => x20_out_3,
   I2 => x44_out_21,
   I3 => x44_out_10,
   I4 => x44_out_6,
   O => W_63_7_i_16_n_0
);
W_63_7_i_17 : LUT5
  generic map(
   INIT => X"ebbe8228"
  )
 port map (
   I0 => x20_out_2,
   I1 => x44_out_5,
   I2 => x44_out_9,
   I3 => x44_out_20,
   I4 => x47_out_2,
   O => W_63_7_i_17_n_0
);
W_63_7_i_2 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x_16,
   I1 => x_23,
   I2 => x_25,
   I3 => W_63_7_i_10_n_0,
   I4 => W_63_7_i_11_n_0,
   O => W_63_7_i_2_n_0
);
W_63_7_i_3 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x_15,
   I1 => x_22,
   I2 => x_24,
   I3 => W_63_7_i_12_n_0,
   I4 => W_63_7_i_13_n_0,
   O => W_63_7_i_3_n_0
);
W_63_7_i_4 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x_14,
   I1 => x_21,
   I2 => x_23,
   I3 => W_63_7_i_14_n_0,
   I4 => W_63_7_i_15_n_0,
   O => W_63_7_i_4_n_0
);
W_63_7_i_5 : LUT5
  generic map(
   INIT => X"ff969600"
  )
 port map (
   I0 => x_13,
   I1 => x_20,
   I2 => x_22,
   I3 => W_63_7_i_16_n_0,
   I4 => W_63_7_i_17_n_0,
   O => W_63_7_i_5_n_0
);
W_63_7_i_6 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_63_7_i_2_n_0,
   I1 => W_63_11_i_16_n_0,
   I2 => x_17,
   I3 => x_24,
   I4 => x_26,
   I5 => W_63_11_i_17_n_0,
   O => W_63_7_i_6_n_0
);
W_63_7_i_7 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_63_7_i_3_n_0,
   I1 => W_63_7_i_10_n_0,
   I2 => x_16,
   I3 => x_23,
   I4 => x_25,
   I5 => W_63_7_i_11_n_0,
   O => W_63_7_i_7_n_0
);
W_63_7_i_8 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_63_7_i_4_n_0,
   I1 => W_63_7_i_12_n_0,
   I2 => x_15,
   I3 => x_22,
   I4 => x_24,
   I5 => W_63_7_i_13_n_0,
   O => W_63_7_i_8_n_0
);
W_63_7_i_9 : LUT6
  generic map(
   INIT => X"6996966996696996"
  )
 port map (
   I0 => W_63_7_i_5_n_0,
   I1 => W_63_7_i_14_n_0,
   I2 => x_14,
   I3 => x_21,
   I4 => x_23,
   I5 => W_63_7_i_15_n_0,
   O => W_63_7_i_9_n_0
);
W_reg_0_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_0_0,
   R => '0',
   Q => W_reg_0_0
);
W_reg_0_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_0_10,
   R => '0',
   Q => W_reg_0_10
);
W_reg_0_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_0_11,
   R => '0',
   Q => W_reg_0_11
);
W_reg_0_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_0_12,
   R => '0',
   Q => W_reg_0_12
);
W_reg_0_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_0_13,
   R => '0',
   Q => W_reg_0_13
);
W_reg_0_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_0_14,
   R => '0',
   Q => W_reg_0_14
);
W_reg_0_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_0_15,
   R => '0',
   Q => W_reg_0_15
);
W_reg_0_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_0_16,
   R => '0',
   Q => W_reg_0_16
);
W_reg_0_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_0_17,
   R => '0',
   Q => W_reg_0_17
);
W_reg_0_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_0_18,
   R => '0',
   Q => W_reg_0_18
);
W_reg_0_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_0_19,
   R => '0',
   Q => W_reg_0_19
);
W_reg_0_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_0_1,
   R => '0',
   Q => W_reg_0_1
);
W_reg_0_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_0_20,
   R => '0',
   Q => W_reg_0_20
);
W_reg_0_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_0_21,
   R => '0',
   Q => W_reg_0_21
);
W_reg_0_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_0_22,
   R => '0',
   Q => W_reg_0_22
);
W_reg_0_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_0_23,
   R => '0',
   Q => W_reg_0_23
);
W_reg_0_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_0_24,
   R => '0',
   Q => W_reg_0_24
);
W_reg_0_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_0_25,
   R => '0',
   Q => W_reg_0_25
);
W_reg_0_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_0_26,
   R => '0',
   Q => W_reg_0_26
);
W_reg_0_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_0_27,
   R => '0',
   Q => W_reg_0_27
);
W_reg_0_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_0_28,
   R => '0',
   Q => W_reg_0_28
);
W_reg_0_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_0_29,
   R => '0',
   Q => W_reg_0_29
);
W_reg_0_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_0_2,
   R => '0',
   Q => W_reg_0_2
);
W_reg_0_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_0_30,
   R => '0',
   Q => W_reg_0_30
);
W_reg_0_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_0_31,
   R => '0',
   Q => W_reg_0_31
);
W_reg_0_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_0_3,
   R => '0',
   Q => W_reg_0_3
);
W_reg_0_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_0_4,
   R => '0',
   Q => W_reg_0_4
);
W_reg_0_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_0_5,
   R => '0',
   Q => W_reg_0_5
);
W_reg_0_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_0_6,
   R => '0',
   Q => W_reg_0_6
);
W_reg_0_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_0_7,
   R => '0',
   Q => W_reg_0_7
);
W_reg_0_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_0_8,
   R => '0',
   Q => W_reg_0_8
);
W_reg_0_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_0_9,
   R => '0',
   Q => W_reg_0_9
);
W_reg_10_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_10_0,
   R => '0',
   Q => W_reg_10_0
);
W_reg_10_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_10_10,
   R => '0',
   Q => W_reg_10_10
);
W_reg_10_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_10_11,
   R => '0',
   Q => W_reg_10_11
);
W_reg_10_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_10_12,
   R => '0',
   Q => W_reg_10_12
);
W_reg_10_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_10_13,
   R => '0',
   Q => W_reg_10_13
);
W_reg_10_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_10_14,
   R => '0',
   Q => W_reg_10_14
);
W_reg_10_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_10_15,
   R => '0',
   Q => W_reg_10_15
);
W_reg_10_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_10_16,
   R => '0',
   Q => W_reg_10_16
);
W_reg_10_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_10_17,
   R => '0',
   Q => W_reg_10_17
);
W_reg_10_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_10_18,
   R => '0',
   Q => W_reg_10_18
);
W_reg_10_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_10_19,
   R => '0',
   Q => W_reg_10_19
);
W_reg_10_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_10_1,
   R => '0',
   Q => W_reg_10_1
);
W_reg_10_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_10_20,
   R => '0',
   Q => W_reg_10_20
);
W_reg_10_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_10_21,
   R => '0',
   Q => W_reg_10_21
);
W_reg_10_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_10_22,
   R => '0',
   Q => W_reg_10_22
);
W_reg_10_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_10_23,
   R => '0',
   Q => W_reg_10_23
);
W_reg_10_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_10_24,
   R => '0',
   Q => W_reg_10_24
);
W_reg_10_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_10_25,
   R => '0',
   Q => W_reg_10_25
);
W_reg_10_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_10_26,
   R => '0',
   Q => W_reg_10_26
);
W_reg_10_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_10_27,
   R => '0',
   Q => W_reg_10_27
);
W_reg_10_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_10_28,
   R => '0',
   Q => W_reg_10_28
);
W_reg_10_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_10_29,
   R => '0',
   Q => W_reg_10_29
);
W_reg_10_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_10_2,
   R => '0',
   Q => W_reg_10_2
);
W_reg_10_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_10_30,
   R => '0',
   Q => W_reg_10_30
);
W_reg_10_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_10_31,
   R => '0',
   Q => W_reg_10_31
);
W_reg_10_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_10_3,
   R => '0',
   Q => W_reg_10_3
);
W_reg_10_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_10_4,
   R => '0',
   Q => W_reg_10_4
);
W_reg_10_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_10_5,
   R => '0',
   Q => W_reg_10_5
);
W_reg_10_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_10_6,
   R => '0',
   Q => W_reg_10_6
);
W_reg_10_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_10_7,
   R => '0',
   Q => W_reg_10_7
);
W_reg_10_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_10_8,
   R => '0',
   Q => W_reg_10_8
);
W_reg_10_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_10_9,
   R => '0',
   Q => W_reg_10_9
);
W_reg_11_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_11_0,
   R => '0',
   Q => W_reg_11_0
);
W_reg_11_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_11_10,
   R => '0',
   Q => W_reg_11_10
);
W_reg_11_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_11_11,
   R => '0',
   Q => W_reg_11_11
);
W_reg_11_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_11_12,
   R => '0',
   Q => W_reg_11_12
);
W_reg_11_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_11_13,
   R => '0',
   Q => W_reg_11_13
);
W_reg_11_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_11_14,
   R => '0',
   Q => W_reg_11_14
);
W_reg_11_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_11_15,
   R => '0',
   Q => W_reg_11_15
);
W_reg_11_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_11_16,
   R => '0',
   Q => W_reg_11_16
);
W_reg_11_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_11_17,
   R => '0',
   Q => W_reg_11_17
);
W_reg_11_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_11_18,
   R => '0',
   Q => W_reg_11_18
);
W_reg_11_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_11_19,
   R => '0',
   Q => W_reg_11_19
);
W_reg_11_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_11_1,
   R => '0',
   Q => W_reg_11_1
);
W_reg_11_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_11_20,
   R => '0',
   Q => W_reg_11_20
);
W_reg_11_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_11_21,
   R => '0',
   Q => W_reg_11_21
);
W_reg_11_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_11_22,
   R => '0',
   Q => W_reg_11_22
);
W_reg_11_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_11_23,
   R => '0',
   Q => W_reg_11_23
);
W_reg_11_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_11_24,
   R => '0',
   Q => W_reg_11_24
);
W_reg_11_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_11_25,
   R => '0',
   Q => W_reg_11_25
);
W_reg_11_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_11_26,
   R => '0',
   Q => W_reg_11_26
);
W_reg_11_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_11_27,
   R => '0',
   Q => W_reg_11_27
);
W_reg_11_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_11_28,
   R => '0',
   Q => W_reg_11_28
);
W_reg_11_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_11_29,
   R => '0',
   Q => W_reg_11_29
);
W_reg_11_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_11_2,
   R => '0',
   Q => W_reg_11_2
);
W_reg_11_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_11_30,
   R => '0',
   Q => W_reg_11_30
);
W_reg_11_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_11_31,
   R => '0',
   Q => W_reg_11_31
);
W_reg_11_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_11_3,
   R => '0',
   Q => W_reg_11_3
);
W_reg_11_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_11_4,
   R => '0',
   Q => W_reg_11_4
);
W_reg_11_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_11_5,
   R => '0',
   Q => W_reg_11_5
);
W_reg_11_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_11_6,
   R => '0',
   Q => W_reg_11_6
);
W_reg_11_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_11_7,
   R => '0',
   Q => W_reg_11_7
);
W_reg_11_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_11_8,
   R => '0',
   Q => W_reg_11_8
);
W_reg_11_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_11_9,
   R => '0',
   Q => W_reg_11_9
);
W_reg_12_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_12_0,
   R => '0',
   Q => W_reg_12_0
);
W_reg_12_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_12_10,
   R => '0',
   Q => W_reg_12_10
);
W_reg_12_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_12_11,
   R => '0',
   Q => W_reg_12_11
);
W_reg_12_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_12_12,
   R => '0',
   Q => W_reg_12_12
);
W_reg_12_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_12_13,
   R => '0',
   Q => W_reg_12_13
);
W_reg_12_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_12_14,
   R => '0',
   Q => W_reg_12_14
);
W_reg_12_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_12_15,
   R => '0',
   Q => W_reg_12_15
);
W_reg_12_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_12_16,
   R => '0',
   Q => W_reg_12_16
);
W_reg_12_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_12_17,
   R => '0',
   Q => W_reg_12_17
);
W_reg_12_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_12_18,
   R => '0',
   Q => W_reg_12_18
);
W_reg_12_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_12_19,
   R => '0',
   Q => W_reg_12_19
);
W_reg_12_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_12_1,
   R => '0',
   Q => W_reg_12_1
);
W_reg_12_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_12_20,
   R => '0',
   Q => W_reg_12_20
);
W_reg_12_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_12_21,
   R => '0',
   Q => W_reg_12_21
);
W_reg_12_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_12_22,
   R => '0',
   Q => W_reg_12_22
);
W_reg_12_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_12_23,
   R => '0',
   Q => W_reg_12_23
);
W_reg_12_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_12_24,
   R => '0',
   Q => W_reg_12_24
);
W_reg_12_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_12_25,
   R => '0',
   Q => W_reg_12_25
);
W_reg_12_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_12_26,
   R => '0',
   Q => W_reg_12_26
);
W_reg_12_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_12_27,
   R => '0',
   Q => W_reg_12_27
);
W_reg_12_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_12_28,
   R => '0',
   Q => W_reg_12_28
);
W_reg_12_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_12_29,
   R => '0',
   Q => W_reg_12_29
);
W_reg_12_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_12_2,
   R => '0',
   Q => W_reg_12_2
);
W_reg_12_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_12_30,
   R => '0',
   Q => W_reg_12_30
);
W_reg_12_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_12_31,
   R => '0',
   Q => W_reg_12_31
);
W_reg_12_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_12_3,
   R => '0',
   Q => W_reg_12_3
);
W_reg_12_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_12_4,
   R => '0',
   Q => W_reg_12_4
);
W_reg_12_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_12_5,
   R => '0',
   Q => W_reg_12_5
);
W_reg_12_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_12_6,
   R => '0',
   Q => W_reg_12_6
);
W_reg_12_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_12_7,
   R => '0',
   Q => W_reg_12_7
);
W_reg_12_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_12_8,
   R => '0',
   Q => W_reg_12_8
);
W_reg_12_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_12_9,
   R => '0',
   Q => W_reg_12_9
);
W_reg_13_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_13_0,
   R => '0',
   Q => W_reg_13_0
);
W_reg_13_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_13_10,
   R => '0',
   Q => W_reg_13_10
);
W_reg_13_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_13_11,
   R => '0',
   Q => W_reg_13_11
);
W_reg_13_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_13_12,
   R => '0',
   Q => W_reg_13_12
);
W_reg_13_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_13_13,
   R => '0',
   Q => W_reg_13_13
);
W_reg_13_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_13_14,
   R => '0',
   Q => W_reg_13_14
);
W_reg_13_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_13_15,
   R => '0',
   Q => W_reg_13_15
);
W_reg_13_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_13_16,
   R => '0',
   Q => W_reg_13_16
);
W_reg_13_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_13_17,
   R => '0',
   Q => W_reg_13_17
);
W_reg_13_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_13_18,
   R => '0',
   Q => W_reg_13_18
);
W_reg_13_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_13_19,
   R => '0',
   Q => W_reg_13_19
);
W_reg_13_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_13_1,
   R => '0',
   Q => W_reg_13_1
);
W_reg_13_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_13_20,
   R => '0',
   Q => W_reg_13_20
);
W_reg_13_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_13_21,
   R => '0',
   Q => W_reg_13_21
);
W_reg_13_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_13_22,
   R => '0',
   Q => W_reg_13_22
);
W_reg_13_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_13_23,
   R => '0',
   Q => W_reg_13_23
);
W_reg_13_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_13_24,
   R => '0',
   Q => W_reg_13_24
);
W_reg_13_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_13_25,
   R => '0',
   Q => W_reg_13_25
);
W_reg_13_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_13_26,
   R => '0',
   Q => W_reg_13_26
);
W_reg_13_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_13_27,
   R => '0',
   Q => W_reg_13_27
);
W_reg_13_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_13_28,
   R => '0',
   Q => W_reg_13_28
);
W_reg_13_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_13_29,
   R => '0',
   Q => W_reg_13_29
);
W_reg_13_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_13_2,
   R => '0',
   Q => W_reg_13_2
);
W_reg_13_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_13_30,
   R => '0',
   Q => W_reg_13_30
);
W_reg_13_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_13_31,
   R => '0',
   Q => W_reg_13_31
);
W_reg_13_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_13_3,
   R => '0',
   Q => W_reg_13_3
);
W_reg_13_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_13_4,
   R => '0',
   Q => W_reg_13_4
);
W_reg_13_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_13_5,
   R => '0',
   Q => W_reg_13_5
);
W_reg_13_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_13_6,
   R => '0',
   Q => W_reg_13_6
);
W_reg_13_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_13_7,
   R => '0',
   Q => W_reg_13_7
);
W_reg_13_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_13_8,
   R => '0',
   Q => W_reg_13_8
);
W_reg_13_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_13_9,
   R => '0',
   Q => W_reg_13_9
);
W_reg_14_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_14_0,
   R => '0',
   Q => W_reg_14_0
);
W_reg_14_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_14_10,
   R => '0',
   Q => W_reg_14_10
);
W_reg_14_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_14_11,
   R => '0',
   Q => W_reg_14_11
);
W_reg_14_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_14_12,
   R => '0',
   Q => W_reg_14_12
);
W_reg_14_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_14_13,
   R => '0',
   Q => W_reg_14_13
);
W_reg_14_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_14_14,
   R => '0',
   Q => W_reg_14_14
);
W_reg_14_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_14_15,
   R => '0',
   Q => W_reg_14_15
);
W_reg_14_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_14_16,
   R => '0',
   Q => W_reg_14_16
);
W_reg_14_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_14_17,
   R => '0',
   Q => W_reg_14_17
);
W_reg_14_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_14_18,
   R => '0',
   Q => W_reg_14_18
);
W_reg_14_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_14_19,
   R => '0',
   Q => W_reg_14_19
);
W_reg_14_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_14_1,
   R => '0',
   Q => W_reg_14_1
);
W_reg_14_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_14_20,
   R => '0',
   Q => W_reg_14_20
);
W_reg_14_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_14_21,
   R => '0',
   Q => W_reg_14_21
);
W_reg_14_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_14_22,
   R => '0',
   Q => W_reg_14_22
);
W_reg_14_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_14_23,
   R => '0',
   Q => W_reg_14_23
);
W_reg_14_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_14_24,
   R => '0',
   Q => W_reg_14_24
);
W_reg_14_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_14_25,
   R => '0',
   Q => W_reg_14_25
);
W_reg_14_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_14_26,
   R => '0',
   Q => W_reg_14_26
);
W_reg_14_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_14_27,
   R => '0',
   Q => W_reg_14_27
);
W_reg_14_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_14_28,
   R => '0',
   Q => W_reg_14_28
);
W_reg_14_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_14_29,
   R => '0',
   Q => W_reg_14_29
);
W_reg_14_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_14_2,
   R => '0',
   Q => W_reg_14_2
);
W_reg_14_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_14_30,
   R => '0',
   Q => W_reg_14_30
);
W_reg_14_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_14_31,
   R => '0',
   Q => W_reg_14_31
);
W_reg_14_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_14_3,
   R => '0',
   Q => W_reg_14_3
);
W_reg_14_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_14_4,
   R => '0',
   Q => W_reg_14_4
);
W_reg_14_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_14_5,
   R => '0',
   Q => W_reg_14_5
);
W_reg_14_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_14_6,
   R => '0',
   Q => W_reg_14_6
);
W_reg_14_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_14_7,
   R => '0',
   Q => W_reg_14_7
);
W_reg_14_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_14_8,
   R => '0',
   Q => W_reg_14_8
);
W_reg_14_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_14_9,
   R => '0',
   Q => W_reg_14_9
);
W_reg_15_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_15_0,
   R => '0',
   Q => W_reg_15_0
);
W_reg_15_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_15_10,
   R => '0',
   Q => W_reg_15_10
);
W_reg_15_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_15_11,
   R => '0',
   Q => W_reg_15_11
);
W_reg_15_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_15_12,
   R => '0',
   Q => W_reg_15_12
);
W_reg_15_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_15_13,
   R => '0',
   Q => W_reg_15_13
);
W_reg_15_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_15_14,
   R => '0',
   Q => W_reg_15_14
);
W_reg_15_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_15_15,
   R => '0',
   Q => W_reg_15_15
);
W_reg_15_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_15_16,
   R => '0',
   Q => W_reg_15_16
);
W_reg_15_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_15_17,
   R => '0',
   Q => W_reg_15_17
);
W_reg_15_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_15_18,
   R => '0',
   Q => W_reg_15_18
);
W_reg_15_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_15_19,
   R => '0',
   Q => W_reg_15_19
);
W_reg_15_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_15_1,
   R => '0',
   Q => W_reg_15_1
);
W_reg_15_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_15_20,
   R => '0',
   Q => W_reg_15_20
);
W_reg_15_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_15_21,
   R => '0',
   Q => W_reg_15_21
);
W_reg_15_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_15_22,
   R => '0',
   Q => W_reg_15_22
);
W_reg_15_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_15_23,
   R => '0',
   Q => W_reg_15_23
);
W_reg_15_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_15_24,
   R => '0',
   Q => W_reg_15_24
);
W_reg_15_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_15_25,
   R => '0',
   Q => W_reg_15_25
);
W_reg_15_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_15_26,
   R => '0',
   Q => W_reg_15_26
);
W_reg_15_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_15_27,
   R => '0',
   Q => W_reg_15_27
);
W_reg_15_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_15_28,
   R => '0',
   Q => W_reg_15_28
);
W_reg_15_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_15_29,
   R => '0',
   Q => W_reg_15_29
);
W_reg_15_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_15_2,
   R => '0',
   Q => W_reg_15_2
);
W_reg_15_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_15_30,
   R => '0',
   Q => W_reg_15_30
);
W_reg_15_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_15_31,
   R => '0',
   Q => W_reg_15_31
);
W_reg_15_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_15_3,
   R => '0',
   Q => W_reg_15_3
);
W_reg_15_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_15_4,
   R => '0',
   Q => W_reg_15_4
);
W_reg_15_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_15_5,
   R => '0',
   Q => W_reg_15_5
);
W_reg_15_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_15_6,
   R => '0',
   Q => W_reg_15_6
);
W_reg_15_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_15_7,
   R => '0',
   Q => W_reg_15_7
);
W_reg_15_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_15_8,
   R => '0',
   Q => W_reg_15_8
);
W_reg_15_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_15_9,
   R => '0',
   Q => W_reg_15_9
);
W_reg_16_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x117_out_0,
   R => '0',
   Q => W_reg_16_0
);
W_reg_16_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x117_out_10,
   R => '0',
   Q => W_reg_16_10
);
W_reg_16_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x117_out_11,
   R => '0',
   Q => W_reg_16_11
);
W_reg_16_11_i_1 : CARRY4
 port map (
   CI => W_reg_16_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_16_11_i_5_n_0,
   DI(1) => W_16_11_i_4_n_0,
   DI(2) => W_16_11_i_3_n_0,
   DI(3) => W_16_11_i_2_n_0,
   S(0) => W_16_11_i_9_n_0,
   S(1) => W_16_11_i_8_n_0,
   S(2) => W_16_11_i_7_n_0,
   S(3) => W_16_11_i_6_n_0,
   CO(0) => W_reg_16_11_i_1_n_3,
   CO(1) => W_reg_16_11_i_1_n_2,
   CO(2) => W_reg_16_11_i_1_n_1,
   CO(3) => W_reg_16_11_i_1_n_0,
   O(0) => x117_out_8,
   O(1) => x117_out_9,
   O(2) => x117_out_10,
   O(3) => x117_out_11
);
W_reg_16_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x117_out_12,
   R => '0',
   Q => W_reg_16_12
);
W_reg_16_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x117_out_13,
   R => '0',
   Q => W_reg_16_13
);
W_reg_16_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x117_out_14,
   R => '0',
   Q => W_reg_16_14
);
W_reg_16_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x117_out_15,
   R => '0',
   Q => W_reg_16_15
);
W_reg_16_15_i_1 : CARRY4
 port map (
   CI => W_reg_16_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_16_15_i_5_n_0,
   DI(1) => W_16_15_i_4_n_0,
   DI(2) => W_16_15_i_3_n_0,
   DI(3) => W_16_15_i_2_n_0,
   S(0) => W_16_15_i_9_n_0,
   S(1) => W_16_15_i_8_n_0,
   S(2) => W_16_15_i_7_n_0,
   S(3) => W_16_15_i_6_n_0,
   CO(0) => W_reg_16_15_i_1_n_3,
   CO(1) => W_reg_16_15_i_1_n_2,
   CO(2) => W_reg_16_15_i_1_n_1,
   CO(3) => W_reg_16_15_i_1_n_0,
   O(0) => x117_out_12,
   O(1) => x117_out_13,
   O(2) => x117_out_14,
   O(3) => x117_out_15
);
W_reg_16_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x117_out_16,
   R => '0',
   Q => W_reg_16_16
);
W_reg_16_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x117_out_17,
   R => '0',
   Q => W_reg_16_17
);
W_reg_16_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x117_out_18,
   R => '0',
   Q => W_reg_16_18
);
W_reg_16_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x117_out_19,
   R => '0',
   Q => W_reg_16_19
);
W_reg_16_19_i_1 : CARRY4
 port map (
   CI => W_reg_16_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_16_19_i_5_n_0,
   DI(1) => W_16_19_i_4_n_0,
   DI(2) => W_16_19_i_3_n_0,
   DI(3) => W_16_19_i_2_n_0,
   S(0) => W_16_19_i_9_n_0,
   S(1) => W_16_19_i_8_n_0,
   S(2) => W_16_19_i_7_n_0,
   S(3) => W_16_19_i_6_n_0,
   CO(0) => W_reg_16_19_i_1_n_3,
   CO(1) => W_reg_16_19_i_1_n_2,
   CO(2) => W_reg_16_19_i_1_n_1,
   CO(3) => W_reg_16_19_i_1_n_0,
   O(0) => x117_out_16,
   O(1) => x117_out_17,
   O(2) => x117_out_18,
   O(3) => x117_out_19
);
W_reg_16_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x117_out_1,
   R => '0',
   Q => W_reg_16_1
);
W_reg_16_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x117_out_20,
   R => '0',
   Q => W_reg_16_20
);
W_reg_16_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x117_out_21,
   R => '0',
   Q => W_reg_16_21
);
W_reg_16_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x117_out_22,
   R => '0',
   Q => W_reg_16_22
);
W_reg_16_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x117_out_23,
   R => '0',
   Q => W_reg_16_23
);
W_reg_16_23_i_1 : CARRY4
 port map (
   CI => W_reg_16_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_16_23_i_5_n_0,
   DI(1) => W_16_23_i_4_n_0,
   DI(2) => W_16_23_i_3_n_0,
   DI(3) => W_16_23_i_2_n_0,
   S(0) => W_16_23_i_9_n_0,
   S(1) => W_16_23_i_8_n_0,
   S(2) => W_16_23_i_7_n_0,
   S(3) => W_16_23_i_6_n_0,
   CO(0) => W_reg_16_23_i_1_n_3,
   CO(1) => W_reg_16_23_i_1_n_2,
   CO(2) => W_reg_16_23_i_1_n_1,
   CO(3) => W_reg_16_23_i_1_n_0,
   O(0) => x117_out_20,
   O(1) => x117_out_21,
   O(2) => x117_out_22,
   O(3) => x117_out_23
);
W_reg_16_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x117_out_24,
   R => '0',
   Q => W_reg_16_24
);
W_reg_16_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x117_out_25,
   R => '0',
   Q => W_reg_16_25
);
W_reg_16_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x117_out_26,
   R => '0',
   Q => W_reg_16_26
);
W_reg_16_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x117_out_27,
   R => '0',
   Q => W_reg_16_27
);
W_reg_16_27_i_1 : CARRY4
 port map (
   CI => W_reg_16_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_16_27_i_5_n_0,
   DI(1) => W_16_27_i_4_n_0,
   DI(2) => W_16_27_i_3_n_0,
   DI(3) => W_16_27_i_2_n_0,
   S(0) => W_16_27_i_9_n_0,
   S(1) => W_16_27_i_8_n_0,
   S(2) => W_16_27_i_7_n_0,
   S(3) => W_16_27_i_6_n_0,
   CO(0) => W_reg_16_27_i_1_n_3,
   CO(1) => W_reg_16_27_i_1_n_2,
   CO(2) => W_reg_16_27_i_1_n_1,
   CO(3) => W_reg_16_27_i_1_n_0,
   O(0) => x117_out_24,
   O(1) => x117_out_25,
   O(2) => x117_out_26,
   O(3) => x117_out_27
);
W_reg_16_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x117_out_28,
   R => '0',
   Q => W_reg_16_28
);
W_reg_16_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x117_out_29,
   R => '0',
   Q => W_reg_16_29
);
W_reg_16_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x117_out_2,
   R => '0',
   Q => W_reg_16_2
);
W_reg_16_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x117_out_30,
   R => '0',
   Q => W_reg_16_30
);
W_reg_16_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x117_out_31,
   R => '0',
   Q => W_reg_16_31
);
W_reg_16_31_i_2 : CARRY4
 port map (
   CI => W_reg_16_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_16_31_i_5_n_0,
   DI(1) => W_16_31_i_4_n_0,
   DI(2) => W_16_31_i_3_n_0,
   DI(3) => '0',
   S(0) => W_16_31_i_9_n_0,
   S(1) => W_16_31_i_8_n_0,
   S(2) => W_16_31_i_7_n_0,
   S(3) => W_16_31_i_6_n_0,
   CO(0) => W_reg_16_31_i_2_n_3,
   CO(1) => W_reg_16_31_i_2_n_2,
   CO(2) => W_reg_16_31_i_2_n_1,
   CO(3) => NLW_W_reg_16_31_i_2_CO_UNCONNECTED_3,
   O(0) => x117_out_28,
   O(1) => x117_out_29,
   O(2) => x117_out_30,
   O(3) => x117_out_31
);
W_reg_16_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x117_out_3,
   R => '0',
   Q => W_reg_16_3
);
W_reg_16_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_16_3_i_5_n_0,
   DI(1) => W_16_3_i_4_n_0,
   DI(2) => W_16_3_i_3_n_0,
   DI(3) => W_16_3_i_2_n_0,
   S(0) => W_16_3_i_9_n_0,
   S(1) => W_16_3_i_8_n_0,
   S(2) => W_16_3_i_7_n_0,
   S(3) => W_16_3_i_6_n_0,
   CO(0) => W_reg_16_3_i_1_n_3,
   CO(1) => W_reg_16_3_i_1_n_2,
   CO(2) => W_reg_16_3_i_1_n_1,
   CO(3) => W_reg_16_3_i_1_n_0,
   O(0) => x117_out_0,
   O(1) => x117_out_1,
   O(2) => x117_out_2,
   O(3) => x117_out_3
);
W_reg_16_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x117_out_4,
   R => '0',
   Q => W_reg_16_4
);
W_reg_16_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x117_out_5,
   R => '0',
   Q => W_reg_16_5
);
W_reg_16_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x117_out_6,
   R => '0',
   Q => W_reg_16_6
);
W_reg_16_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x117_out_7,
   R => '0',
   Q => W_reg_16_7
);
W_reg_16_7_i_1 : CARRY4
 port map (
   CI => W_reg_16_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_16_7_i_5_n_0,
   DI(1) => W_16_7_i_4_n_0,
   DI(2) => W_16_7_i_3_n_0,
   DI(3) => W_16_7_i_2_n_0,
   S(0) => W_16_7_i_9_n_0,
   S(1) => W_16_7_i_8_n_0,
   S(2) => W_16_7_i_7_n_0,
   S(3) => W_16_7_i_6_n_0,
   CO(0) => W_reg_16_7_i_1_n_3,
   CO(1) => W_reg_16_7_i_1_n_2,
   CO(2) => W_reg_16_7_i_1_n_1,
   CO(3) => W_reg_16_7_i_1_n_0,
   O(0) => x117_out_4,
   O(1) => x117_out_5,
   O(2) => x117_out_6,
   O(3) => x117_out_7
);
W_reg_16_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x117_out_8,
   R => '0',
   Q => W_reg_16_8
);
W_reg_16_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x117_out_9,
   R => '0',
   Q => W_reg_16_9
);
W_reg_17_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x116_out_0,
   R => '0',
   Q => W_reg_17_0
);
W_reg_17_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x116_out_10,
   R => '0',
   Q => W_reg_17_10
);
W_reg_17_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x116_out_11,
   R => '0',
   Q => W_reg_17_11
);
W_reg_17_11_i_1 : CARRY4
 port map (
   CI => W_reg_17_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_17_11_i_5_n_0,
   DI(1) => W_17_11_i_4_n_0,
   DI(2) => W_17_11_i_3_n_0,
   DI(3) => W_17_11_i_2_n_0,
   S(0) => W_17_11_i_9_n_0,
   S(1) => W_17_11_i_8_n_0,
   S(2) => W_17_11_i_7_n_0,
   S(3) => W_17_11_i_6_n_0,
   CO(0) => W_reg_17_11_i_1_n_3,
   CO(1) => W_reg_17_11_i_1_n_2,
   CO(2) => W_reg_17_11_i_1_n_1,
   CO(3) => W_reg_17_11_i_1_n_0,
   O(0) => x116_out_8,
   O(1) => x116_out_9,
   O(2) => x116_out_10,
   O(3) => x116_out_11
);
W_reg_17_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x116_out_12,
   R => '0',
   Q => W_reg_17_12
);
W_reg_17_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x116_out_13,
   R => '0',
   Q => W_reg_17_13
);
W_reg_17_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x116_out_14,
   R => '0',
   Q => W_reg_17_14
);
W_reg_17_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x116_out_15,
   R => '0',
   Q => W_reg_17_15
);
W_reg_17_15_i_1 : CARRY4
 port map (
   CI => W_reg_17_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_17_15_i_5_n_0,
   DI(1) => W_17_15_i_4_n_0,
   DI(2) => W_17_15_i_3_n_0,
   DI(3) => W_17_15_i_2_n_0,
   S(0) => W_17_15_i_9_n_0,
   S(1) => W_17_15_i_8_n_0,
   S(2) => W_17_15_i_7_n_0,
   S(3) => W_17_15_i_6_n_0,
   CO(0) => W_reg_17_15_i_1_n_3,
   CO(1) => W_reg_17_15_i_1_n_2,
   CO(2) => W_reg_17_15_i_1_n_1,
   CO(3) => W_reg_17_15_i_1_n_0,
   O(0) => x116_out_12,
   O(1) => x116_out_13,
   O(2) => x116_out_14,
   O(3) => x116_out_15
);
W_reg_17_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x116_out_16,
   R => '0',
   Q => W_reg_17_16
);
W_reg_17_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x116_out_17,
   R => '0',
   Q => W_reg_17_17
);
W_reg_17_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x116_out_18,
   R => '0',
   Q => W_reg_17_18
);
W_reg_17_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x116_out_19,
   R => '0',
   Q => W_reg_17_19
);
W_reg_17_19_i_1 : CARRY4
 port map (
   CI => W_reg_17_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_17_19_i_5_n_0,
   DI(1) => W_17_19_i_4_n_0,
   DI(2) => W_17_19_i_3_n_0,
   DI(3) => W_17_19_i_2_n_0,
   S(0) => W_17_19_i_9_n_0,
   S(1) => W_17_19_i_8_n_0,
   S(2) => W_17_19_i_7_n_0,
   S(3) => W_17_19_i_6_n_0,
   CO(0) => W_reg_17_19_i_1_n_3,
   CO(1) => W_reg_17_19_i_1_n_2,
   CO(2) => W_reg_17_19_i_1_n_1,
   CO(3) => W_reg_17_19_i_1_n_0,
   O(0) => x116_out_16,
   O(1) => x116_out_17,
   O(2) => x116_out_18,
   O(3) => x116_out_19
);
W_reg_17_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x116_out_1,
   R => '0',
   Q => W_reg_17_1
);
W_reg_17_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x116_out_20,
   R => '0',
   Q => W_reg_17_20
);
W_reg_17_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x116_out_21,
   R => '0',
   Q => W_reg_17_21
);
W_reg_17_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x116_out_22,
   R => '0',
   Q => W_reg_17_22
);
W_reg_17_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x116_out_23,
   R => '0',
   Q => W_reg_17_23
);
W_reg_17_23_i_1 : CARRY4
 port map (
   CI => W_reg_17_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_17_23_i_5_n_0,
   DI(1) => W_17_23_i_4_n_0,
   DI(2) => W_17_23_i_3_n_0,
   DI(3) => W_17_23_i_2_n_0,
   S(0) => W_17_23_i_9_n_0,
   S(1) => W_17_23_i_8_n_0,
   S(2) => W_17_23_i_7_n_0,
   S(3) => W_17_23_i_6_n_0,
   CO(0) => W_reg_17_23_i_1_n_3,
   CO(1) => W_reg_17_23_i_1_n_2,
   CO(2) => W_reg_17_23_i_1_n_1,
   CO(3) => W_reg_17_23_i_1_n_0,
   O(0) => x116_out_20,
   O(1) => x116_out_21,
   O(2) => x116_out_22,
   O(3) => x116_out_23
);
W_reg_17_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x116_out_24,
   R => '0',
   Q => W_reg_17_24
);
W_reg_17_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x116_out_25,
   R => '0',
   Q => W_reg_17_25
);
W_reg_17_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x116_out_26,
   R => '0',
   Q => W_reg_17_26
);
W_reg_17_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x116_out_27,
   R => '0',
   Q => W_reg_17_27
);
W_reg_17_27_i_1 : CARRY4
 port map (
   CI => W_reg_17_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_17_27_i_5_n_0,
   DI(1) => W_17_27_i_4_n_0,
   DI(2) => W_17_27_i_3_n_0,
   DI(3) => W_17_27_i_2_n_0,
   S(0) => W_17_27_i_9_n_0,
   S(1) => W_17_27_i_8_n_0,
   S(2) => W_17_27_i_7_n_0,
   S(3) => W_17_27_i_6_n_0,
   CO(0) => W_reg_17_27_i_1_n_3,
   CO(1) => W_reg_17_27_i_1_n_2,
   CO(2) => W_reg_17_27_i_1_n_1,
   CO(3) => W_reg_17_27_i_1_n_0,
   O(0) => x116_out_24,
   O(1) => x116_out_25,
   O(2) => x116_out_26,
   O(3) => x116_out_27
);
W_reg_17_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x116_out_28,
   R => '0',
   Q => W_reg_17_28
);
W_reg_17_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x116_out_29,
   R => '0',
   Q => W_reg_17_29
);
W_reg_17_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x116_out_2,
   R => '0',
   Q => W_reg_17_2
);
W_reg_17_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x116_out_30,
   R => '0',
   Q => W_reg_17_30
);
W_reg_17_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x116_out_31,
   R => '0',
   Q => W_reg_17_31
);
W_reg_17_31_i_1 : CARRY4
 port map (
   CI => W_reg_17_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_17_31_i_4_n_0,
   DI(1) => W_17_31_i_3_n_0,
   DI(2) => W_17_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_17_31_i_8_n_0,
   S(1) => W_17_31_i_7_n_0,
   S(2) => W_17_31_i_6_n_0,
   S(3) => W_17_31_i_5_n_0,
   CO(0) => W_reg_17_31_i_1_n_3,
   CO(1) => W_reg_17_31_i_1_n_2,
   CO(2) => W_reg_17_31_i_1_n_1,
   CO(3) => NLW_W_reg_17_31_i_1_CO_UNCONNECTED_3,
   O(0) => x116_out_28,
   O(1) => x116_out_29,
   O(2) => x116_out_30,
   O(3) => x116_out_31
);
W_reg_17_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x116_out_3,
   R => '0',
   Q => W_reg_17_3
);
W_reg_17_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_17_3_i_5_n_0,
   DI(1) => W_17_3_i_4_n_0,
   DI(2) => W_17_3_i_3_n_0,
   DI(3) => W_17_3_i_2_n_0,
   S(0) => W_17_3_i_9_n_0,
   S(1) => W_17_3_i_8_n_0,
   S(2) => W_17_3_i_7_n_0,
   S(3) => W_17_3_i_6_n_0,
   CO(0) => W_reg_17_3_i_1_n_3,
   CO(1) => W_reg_17_3_i_1_n_2,
   CO(2) => W_reg_17_3_i_1_n_1,
   CO(3) => W_reg_17_3_i_1_n_0,
   O(0) => x116_out_0,
   O(1) => x116_out_1,
   O(2) => x116_out_2,
   O(3) => x116_out_3
);
W_reg_17_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x116_out_4,
   R => '0',
   Q => W_reg_17_4
);
W_reg_17_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x116_out_5,
   R => '0',
   Q => W_reg_17_5
);
W_reg_17_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x116_out_6,
   R => '0',
   Q => W_reg_17_6
);
W_reg_17_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x116_out_7,
   R => '0',
   Q => W_reg_17_7
);
W_reg_17_7_i_1 : CARRY4
 port map (
   CI => W_reg_17_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_17_7_i_5_n_0,
   DI(1) => W_17_7_i_4_n_0,
   DI(2) => W_17_7_i_3_n_0,
   DI(3) => W_17_7_i_2_n_0,
   S(0) => W_17_7_i_9_n_0,
   S(1) => W_17_7_i_8_n_0,
   S(2) => W_17_7_i_7_n_0,
   S(3) => W_17_7_i_6_n_0,
   CO(0) => W_reg_17_7_i_1_n_3,
   CO(1) => W_reg_17_7_i_1_n_2,
   CO(2) => W_reg_17_7_i_1_n_1,
   CO(3) => W_reg_17_7_i_1_n_0,
   O(0) => x116_out_4,
   O(1) => x116_out_5,
   O(2) => x116_out_6,
   O(3) => x116_out_7
);
W_reg_17_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x116_out_8,
   R => '0',
   Q => W_reg_17_8
);
W_reg_17_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x116_out_9,
   R => '0',
   Q => W_reg_17_9
);
W_reg_18_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x115_out_0,
   R => '0',
   Q => W_reg_18_0
);
W_reg_18_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x115_out_10,
   R => '0',
   Q => W_reg_18_10
);
W_reg_18_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x115_out_11,
   R => '0',
   Q => W_reg_18_11
);
W_reg_18_11_i_1 : CARRY4
 port map (
   CI => W_reg_18_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_18_11_i_5_n_0,
   DI(1) => W_18_11_i_4_n_0,
   DI(2) => W_18_11_i_3_n_0,
   DI(3) => W_18_11_i_2_n_0,
   S(0) => W_18_11_i_9_n_0,
   S(1) => W_18_11_i_8_n_0,
   S(2) => W_18_11_i_7_n_0,
   S(3) => W_18_11_i_6_n_0,
   CO(0) => W_reg_18_11_i_1_n_3,
   CO(1) => W_reg_18_11_i_1_n_2,
   CO(2) => W_reg_18_11_i_1_n_1,
   CO(3) => W_reg_18_11_i_1_n_0,
   O(0) => x115_out_8,
   O(1) => x115_out_9,
   O(2) => x115_out_10,
   O(3) => x115_out_11
);
W_reg_18_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x115_out_12,
   R => '0',
   Q => W_reg_18_12
);
W_reg_18_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x115_out_13,
   R => '0',
   Q => W_reg_18_13
);
W_reg_18_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x115_out_14,
   R => '0',
   Q => W_reg_18_14
);
W_reg_18_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x115_out_15,
   R => '0',
   Q => W_reg_18_15
);
W_reg_18_15_i_1 : CARRY4
 port map (
   CI => W_reg_18_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_18_15_i_5_n_0,
   DI(1) => W_18_15_i_4_n_0,
   DI(2) => W_18_15_i_3_n_0,
   DI(3) => W_18_15_i_2_n_0,
   S(0) => W_18_15_i_9_n_0,
   S(1) => W_18_15_i_8_n_0,
   S(2) => W_18_15_i_7_n_0,
   S(3) => W_18_15_i_6_n_0,
   CO(0) => W_reg_18_15_i_1_n_3,
   CO(1) => W_reg_18_15_i_1_n_2,
   CO(2) => W_reg_18_15_i_1_n_1,
   CO(3) => W_reg_18_15_i_1_n_0,
   O(0) => x115_out_12,
   O(1) => x115_out_13,
   O(2) => x115_out_14,
   O(3) => x115_out_15
);
W_reg_18_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x115_out_16,
   R => '0',
   Q => W_reg_18_16
);
W_reg_18_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x115_out_17,
   R => '0',
   Q => W_reg_18_17
);
W_reg_18_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x115_out_18,
   R => '0',
   Q => W_reg_18_18
);
W_reg_18_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x115_out_19,
   R => '0',
   Q => W_reg_18_19
);
W_reg_18_19_i_1 : CARRY4
 port map (
   CI => W_reg_18_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_18_19_i_5_n_0,
   DI(1) => W_18_19_i_4_n_0,
   DI(2) => W_18_19_i_3_n_0,
   DI(3) => W_18_19_i_2_n_0,
   S(0) => W_18_19_i_9_n_0,
   S(1) => W_18_19_i_8_n_0,
   S(2) => W_18_19_i_7_n_0,
   S(3) => W_18_19_i_6_n_0,
   CO(0) => W_reg_18_19_i_1_n_3,
   CO(1) => W_reg_18_19_i_1_n_2,
   CO(2) => W_reg_18_19_i_1_n_1,
   CO(3) => W_reg_18_19_i_1_n_0,
   O(0) => x115_out_16,
   O(1) => x115_out_17,
   O(2) => x115_out_18,
   O(3) => x115_out_19
);
W_reg_18_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x115_out_1,
   R => '0',
   Q => W_reg_18_1
);
W_reg_18_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x115_out_20,
   R => '0',
   Q => W_reg_18_20
);
W_reg_18_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x115_out_21,
   R => '0',
   Q => W_reg_18_21
);
W_reg_18_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x115_out_22,
   R => '0',
   Q => W_reg_18_22
);
W_reg_18_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x115_out_23,
   R => '0',
   Q => W_reg_18_23
);
W_reg_18_23_i_1 : CARRY4
 port map (
   CI => W_reg_18_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_18_23_i_5_n_0,
   DI(1) => W_18_23_i_4_n_0,
   DI(2) => W_18_23_i_3_n_0,
   DI(3) => W_18_23_i_2_n_0,
   S(0) => W_18_23_i_9_n_0,
   S(1) => W_18_23_i_8_n_0,
   S(2) => W_18_23_i_7_n_0,
   S(3) => W_18_23_i_6_n_0,
   CO(0) => W_reg_18_23_i_1_n_3,
   CO(1) => W_reg_18_23_i_1_n_2,
   CO(2) => W_reg_18_23_i_1_n_1,
   CO(3) => W_reg_18_23_i_1_n_0,
   O(0) => x115_out_20,
   O(1) => x115_out_21,
   O(2) => x115_out_22,
   O(3) => x115_out_23
);
W_reg_18_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x115_out_24,
   R => '0',
   Q => W_reg_18_24
);
W_reg_18_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x115_out_25,
   R => '0',
   Q => W_reg_18_25
);
W_reg_18_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x115_out_26,
   R => '0',
   Q => W_reg_18_26
);
W_reg_18_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x115_out_27,
   R => '0',
   Q => W_reg_18_27
);
W_reg_18_27_i_1 : CARRY4
 port map (
   CI => W_reg_18_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_18_27_i_5_n_0,
   DI(1) => W_18_27_i_4_n_0,
   DI(2) => W_18_27_i_3_n_0,
   DI(3) => W_18_27_i_2_n_0,
   S(0) => W_18_27_i_9_n_0,
   S(1) => W_18_27_i_8_n_0,
   S(2) => W_18_27_i_7_n_0,
   S(3) => W_18_27_i_6_n_0,
   CO(0) => W_reg_18_27_i_1_n_3,
   CO(1) => W_reg_18_27_i_1_n_2,
   CO(2) => W_reg_18_27_i_1_n_1,
   CO(3) => W_reg_18_27_i_1_n_0,
   O(0) => x115_out_24,
   O(1) => x115_out_25,
   O(2) => x115_out_26,
   O(3) => x115_out_27
);
W_reg_18_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x115_out_28,
   R => '0',
   Q => W_reg_18_28
);
W_reg_18_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x115_out_29,
   R => '0',
   Q => W_reg_18_29
);
W_reg_18_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x115_out_2,
   R => '0',
   Q => W_reg_18_2
);
W_reg_18_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x115_out_30,
   R => '0',
   Q => W_reg_18_30
);
W_reg_18_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x115_out_31,
   R => '0',
   Q => W_reg_18_31
);
W_reg_18_31_i_1 : CARRY4
 port map (
   CI => W_reg_18_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_18_31_i_4_n_0,
   DI(1) => W_18_31_i_3_n_0,
   DI(2) => W_18_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_18_31_i_8_n_0,
   S(1) => W_18_31_i_7_n_0,
   S(2) => W_18_31_i_6_n_0,
   S(3) => W_18_31_i_5_n_0,
   CO(0) => W_reg_18_31_i_1_n_3,
   CO(1) => W_reg_18_31_i_1_n_2,
   CO(2) => W_reg_18_31_i_1_n_1,
   CO(3) => NLW_W_reg_18_31_i_1_CO_UNCONNECTED_3,
   O(0) => x115_out_28,
   O(1) => x115_out_29,
   O(2) => x115_out_30,
   O(3) => x115_out_31
);
W_reg_18_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x115_out_3,
   R => '0',
   Q => W_reg_18_3
);
W_reg_18_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_18_3_i_5_n_0,
   DI(1) => W_18_3_i_4_n_0,
   DI(2) => W_18_3_i_3_n_0,
   DI(3) => W_18_3_i_2_n_0,
   S(0) => W_18_3_i_9_n_0,
   S(1) => W_18_3_i_8_n_0,
   S(2) => W_18_3_i_7_n_0,
   S(3) => W_18_3_i_6_n_0,
   CO(0) => W_reg_18_3_i_1_n_3,
   CO(1) => W_reg_18_3_i_1_n_2,
   CO(2) => W_reg_18_3_i_1_n_1,
   CO(3) => W_reg_18_3_i_1_n_0,
   O(0) => x115_out_0,
   O(1) => x115_out_1,
   O(2) => x115_out_2,
   O(3) => x115_out_3
);
W_reg_18_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x115_out_4,
   R => '0',
   Q => W_reg_18_4
);
W_reg_18_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x115_out_5,
   R => '0',
   Q => W_reg_18_5
);
W_reg_18_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x115_out_6,
   R => '0',
   Q => W_reg_18_6
);
W_reg_18_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x115_out_7,
   R => '0',
   Q => W_reg_18_7
);
W_reg_18_7_i_1 : CARRY4
 port map (
   CI => W_reg_18_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_18_7_i_5_n_0,
   DI(1) => W_18_7_i_4_n_0,
   DI(2) => W_18_7_i_3_n_0,
   DI(3) => W_18_7_i_2_n_0,
   S(0) => W_18_7_i_9_n_0,
   S(1) => W_18_7_i_8_n_0,
   S(2) => W_18_7_i_7_n_0,
   S(3) => W_18_7_i_6_n_0,
   CO(0) => W_reg_18_7_i_1_n_3,
   CO(1) => W_reg_18_7_i_1_n_2,
   CO(2) => W_reg_18_7_i_1_n_1,
   CO(3) => W_reg_18_7_i_1_n_0,
   O(0) => x115_out_4,
   O(1) => x115_out_5,
   O(2) => x115_out_6,
   O(3) => x115_out_7
);
W_reg_18_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x115_out_8,
   R => '0',
   Q => W_reg_18_8
);
W_reg_18_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x115_out_9,
   R => '0',
   Q => W_reg_18_9
);
W_reg_19_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x114_out_0,
   R => '0',
   Q => W_reg_19_0
);
W_reg_19_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x114_out_10,
   R => '0',
   Q => W_reg_19_10
);
W_reg_19_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x114_out_11,
   R => '0',
   Q => W_reg_19_11
);
W_reg_19_11_i_1 : CARRY4
 port map (
   CI => W_reg_19_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_19_11_i_5_n_0,
   DI(1) => W_19_11_i_4_n_0,
   DI(2) => W_19_11_i_3_n_0,
   DI(3) => W_19_11_i_2_n_0,
   S(0) => W_19_11_i_9_n_0,
   S(1) => W_19_11_i_8_n_0,
   S(2) => W_19_11_i_7_n_0,
   S(3) => W_19_11_i_6_n_0,
   CO(0) => W_reg_19_11_i_1_n_3,
   CO(1) => W_reg_19_11_i_1_n_2,
   CO(2) => W_reg_19_11_i_1_n_1,
   CO(3) => W_reg_19_11_i_1_n_0,
   O(0) => x114_out_8,
   O(1) => x114_out_9,
   O(2) => x114_out_10,
   O(3) => x114_out_11
);
W_reg_19_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x114_out_12,
   R => '0',
   Q => W_reg_19_12
);
W_reg_19_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x114_out_13,
   R => '0',
   Q => W_reg_19_13
);
W_reg_19_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x114_out_14,
   R => '0',
   Q => W_reg_19_14
);
W_reg_19_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x114_out_15,
   R => '0',
   Q => W_reg_19_15
);
W_reg_19_15_i_1 : CARRY4
 port map (
   CI => W_reg_19_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_19_15_i_5_n_0,
   DI(1) => W_19_15_i_4_n_0,
   DI(2) => W_19_15_i_3_n_0,
   DI(3) => W_19_15_i_2_n_0,
   S(0) => W_19_15_i_9_n_0,
   S(1) => W_19_15_i_8_n_0,
   S(2) => W_19_15_i_7_n_0,
   S(3) => W_19_15_i_6_n_0,
   CO(0) => W_reg_19_15_i_1_n_3,
   CO(1) => W_reg_19_15_i_1_n_2,
   CO(2) => W_reg_19_15_i_1_n_1,
   CO(3) => W_reg_19_15_i_1_n_0,
   O(0) => x114_out_12,
   O(1) => x114_out_13,
   O(2) => x114_out_14,
   O(3) => x114_out_15
);
W_reg_19_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x114_out_16,
   R => '0',
   Q => W_reg_19_16
);
W_reg_19_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x114_out_17,
   R => '0',
   Q => W_reg_19_17
);
W_reg_19_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x114_out_18,
   R => '0',
   Q => W_reg_19_18
);
W_reg_19_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x114_out_19,
   R => '0',
   Q => W_reg_19_19
);
W_reg_19_19_i_1 : CARRY4
 port map (
   CI => W_reg_19_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_19_19_i_5_n_0,
   DI(1) => W_19_19_i_4_n_0,
   DI(2) => W_19_19_i_3_n_0,
   DI(3) => W_19_19_i_2_n_0,
   S(0) => W_19_19_i_9_n_0,
   S(1) => W_19_19_i_8_n_0,
   S(2) => W_19_19_i_7_n_0,
   S(3) => W_19_19_i_6_n_0,
   CO(0) => W_reg_19_19_i_1_n_3,
   CO(1) => W_reg_19_19_i_1_n_2,
   CO(2) => W_reg_19_19_i_1_n_1,
   CO(3) => W_reg_19_19_i_1_n_0,
   O(0) => x114_out_16,
   O(1) => x114_out_17,
   O(2) => x114_out_18,
   O(3) => x114_out_19
);
W_reg_19_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x114_out_1,
   R => '0',
   Q => W_reg_19_1
);
W_reg_19_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x114_out_20,
   R => '0',
   Q => W_reg_19_20
);
W_reg_19_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x114_out_21,
   R => '0',
   Q => W_reg_19_21
);
W_reg_19_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x114_out_22,
   R => '0',
   Q => W_reg_19_22
);
W_reg_19_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x114_out_23,
   R => '0',
   Q => W_reg_19_23
);
W_reg_19_23_i_1 : CARRY4
 port map (
   CI => W_reg_19_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_19_23_i_5_n_0,
   DI(1) => W_19_23_i_4_n_0,
   DI(2) => W_19_23_i_3_n_0,
   DI(3) => W_19_23_i_2_n_0,
   S(0) => W_19_23_i_9_n_0,
   S(1) => W_19_23_i_8_n_0,
   S(2) => W_19_23_i_7_n_0,
   S(3) => W_19_23_i_6_n_0,
   CO(0) => W_reg_19_23_i_1_n_3,
   CO(1) => W_reg_19_23_i_1_n_2,
   CO(2) => W_reg_19_23_i_1_n_1,
   CO(3) => W_reg_19_23_i_1_n_0,
   O(0) => x114_out_20,
   O(1) => x114_out_21,
   O(2) => x114_out_22,
   O(3) => x114_out_23
);
W_reg_19_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x114_out_24,
   R => '0',
   Q => W_reg_19_24
);
W_reg_19_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x114_out_25,
   R => '0',
   Q => W_reg_19_25
);
W_reg_19_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x114_out_26,
   R => '0',
   Q => W_reg_19_26
);
W_reg_19_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x114_out_27,
   R => '0',
   Q => W_reg_19_27
);
W_reg_19_27_i_1 : CARRY4
 port map (
   CI => W_reg_19_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_19_27_i_5_n_0,
   DI(1) => W_19_27_i_4_n_0,
   DI(2) => W_19_27_i_3_n_0,
   DI(3) => W_19_27_i_2_n_0,
   S(0) => W_19_27_i_9_n_0,
   S(1) => W_19_27_i_8_n_0,
   S(2) => W_19_27_i_7_n_0,
   S(3) => W_19_27_i_6_n_0,
   CO(0) => W_reg_19_27_i_1_n_3,
   CO(1) => W_reg_19_27_i_1_n_2,
   CO(2) => W_reg_19_27_i_1_n_1,
   CO(3) => W_reg_19_27_i_1_n_0,
   O(0) => x114_out_24,
   O(1) => x114_out_25,
   O(2) => x114_out_26,
   O(3) => x114_out_27
);
W_reg_19_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x114_out_28,
   R => '0',
   Q => W_reg_19_28
);
W_reg_19_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x114_out_29,
   R => '0',
   Q => W_reg_19_29
);
W_reg_19_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x114_out_2,
   R => '0',
   Q => W_reg_19_2
);
W_reg_19_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x114_out_30,
   R => '0',
   Q => W_reg_19_30
);
W_reg_19_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x114_out_31,
   R => '0',
   Q => W_reg_19_31
);
W_reg_19_31_i_1 : CARRY4
 port map (
   CI => W_reg_19_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_19_31_i_4_n_0,
   DI(1) => W_19_31_i_3_n_0,
   DI(2) => W_19_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_19_31_i_8_n_0,
   S(1) => W_19_31_i_7_n_0,
   S(2) => W_19_31_i_6_n_0,
   S(3) => W_19_31_i_5_n_0,
   CO(0) => W_reg_19_31_i_1_n_3,
   CO(1) => W_reg_19_31_i_1_n_2,
   CO(2) => W_reg_19_31_i_1_n_1,
   CO(3) => NLW_W_reg_19_31_i_1_CO_UNCONNECTED_3,
   O(0) => x114_out_28,
   O(1) => x114_out_29,
   O(2) => x114_out_30,
   O(3) => x114_out_31
);
W_reg_19_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x114_out_3,
   R => '0',
   Q => W_reg_19_3
);
W_reg_19_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_19_3_i_5_n_0,
   DI(1) => W_19_3_i_4_n_0,
   DI(2) => W_19_3_i_3_n_0,
   DI(3) => W_19_3_i_2_n_0,
   S(0) => W_19_3_i_9_n_0,
   S(1) => W_19_3_i_8_n_0,
   S(2) => W_19_3_i_7_n_0,
   S(3) => W_19_3_i_6_n_0,
   CO(0) => W_reg_19_3_i_1_n_3,
   CO(1) => W_reg_19_3_i_1_n_2,
   CO(2) => W_reg_19_3_i_1_n_1,
   CO(3) => W_reg_19_3_i_1_n_0,
   O(0) => x114_out_0,
   O(1) => x114_out_1,
   O(2) => x114_out_2,
   O(3) => x114_out_3
);
W_reg_19_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x114_out_4,
   R => '0',
   Q => W_reg_19_4
);
W_reg_19_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x114_out_5,
   R => '0',
   Q => W_reg_19_5
);
W_reg_19_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x114_out_6,
   R => '0',
   Q => W_reg_19_6
);
W_reg_19_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x114_out_7,
   R => '0',
   Q => W_reg_19_7
);
W_reg_19_7_i_1 : CARRY4
 port map (
   CI => W_reg_19_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_19_7_i_5_n_0,
   DI(1) => W_19_7_i_4_n_0,
   DI(2) => W_19_7_i_3_n_0,
   DI(3) => W_19_7_i_2_n_0,
   S(0) => W_19_7_i_9_n_0,
   S(1) => W_19_7_i_8_n_0,
   S(2) => W_19_7_i_7_n_0,
   S(3) => W_19_7_i_6_n_0,
   CO(0) => W_reg_19_7_i_1_n_3,
   CO(1) => W_reg_19_7_i_1_n_2,
   CO(2) => W_reg_19_7_i_1_n_1,
   CO(3) => W_reg_19_7_i_1_n_0,
   O(0) => x114_out_4,
   O(1) => x114_out_5,
   O(2) => x114_out_6,
   O(3) => x114_out_7
);
W_reg_19_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x114_out_8,
   R => '0',
   Q => W_reg_19_8
);
W_reg_19_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x114_out_9,
   R => '0',
   Q => W_reg_19_9
);
W_reg_1_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_1_0,
   R => '0',
   Q => W_reg_1_0
);
W_reg_1_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_1_10,
   R => '0',
   Q => W_reg_1_10
);
W_reg_1_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_1_11,
   R => '0',
   Q => W_reg_1_11
);
W_reg_1_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_1_12,
   R => '0',
   Q => W_reg_1_12
);
W_reg_1_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_1_13,
   R => '0',
   Q => W_reg_1_13
);
W_reg_1_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_1_14,
   R => '0',
   Q => W_reg_1_14
);
W_reg_1_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_1_15,
   R => '0',
   Q => W_reg_1_15
);
W_reg_1_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_1_16,
   R => '0',
   Q => W_reg_1_16
);
W_reg_1_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_1_17,
   R => '0',
   Q => W_reg_1_17
);
W_reg_1_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_1_18,
   R => '0',
   Q => W_reg_1_18
);
W_reg_1_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_1_19,
   R => '0',
   Q => W_reg_1_19
);
W_reg_1_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_1_1,
   R => '0',
   Q => W_reg_1_1
);
W_reg_1_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_1_20,
   R => '0',
   Q => W_reg_1_20
);
W_reg_1_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_1_21,
   R => '0',
   Q => W_reg_1_21
);
W_reg_1_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_1_22,
   R => '0',
   Q => W_reg_1_22
);
W_reg_1_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_1_23,
   R => '0',
   Q => W_reg_1_23
);
W_reg_1_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_1_24,
   R => '0',
   Q => W_reg_1_24
);
W_reg_1_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_1_25,
   R => '0',
   Q => W_reg_1_25
);
W_reg_1_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_1_26,
   R => '0',
   Q => W_reg_1_26
);
W_reg_1_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_1_27,
   R => '0',
   Q => W_reg_1_27
);
W_reg_1_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_1_28,
   R => '0',
   Q => W_reg_1_28
);
W_reg_1_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_1_29,
   R => '0',
   Q => W_reg_1_29
);
W_reg_1_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_1_2,
   R => '0',
   Q => W_reg_1_2
);
W_reg_1_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_1_30,
   R => '0',
   Q => W_reg_1_30
);
W_reg_1_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_1_31,
   R => '0',
   Q => W_reg_1_31
);
W_reg_1_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_1_3,
   R => '0',
   Q => W_reg_1_3
);
W_reg_1_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_1_4,
   R => '0',
   Q => W_reg_1_4
);
W_reg_1_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_1_5,
   R => '0',
   Q => W_reg_1_5
);
W_reg_1_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_1_6,
   R => '0',
   Q => W_reg_1_6
);
W_reg_1_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_1_7,
   R => '0',
   Q => W_reg_1_7
);
W_reg_1_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_1_8,
   R => '0',
   Q => W_reg_1_8
);
W_reg_1_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_1_9,
   R => '0',
   Q => W_reg_1_9
);
W_reg_20_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x113_out_0,
   R => '0',
   Q => W_reg_20_0
);
W_reg_20_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x113_out_10,
   R => '0',
   Q => W_reg_20_10
);
W_reg_20_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x113_out_11,
   R => '0',
   Q => W_reg_20_11
);
W_reg_20_11_i_1 : CARRY4
 port map (
   CI => W_reg_20_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_20_11_i_5_n_0,
   DI(1) => W_20_11_i_4_n_0,
   DI(2) => W_20_11_i_3_n_0,
   DI(3) => W_20_11_i_2_n_0,
   S(0) => W_20_11_i_9_n_0,
   S(1) => W_20_11_i_8_n_0,
   S(2) => W_20_11_i_7_n_0,
   S(3) => W_20_11_i_6_n_0,
   CO(0) => W_reg_20_11_i_1_n_3,
   CO(1) => W_reg_20_11_i_1_n_2,
   CO(2) => W_reg_20_11_i_1_n_1,
   CO(3) => W_reg_20_11_i_1_n_0,
   O(0) => x113_out_8,
   O(1) => x113_out_9,
   O(2) => x113_out_10,
   O(3) => x113_out_11
);
W_reg_20_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x113_out_12,
   R => '0',
   Q => W_reg_20_12
);
W_reg_20_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x113_out_13,
   R => '0',
   Q => W_reg_20_13
);
W_reg_20_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x113_out_14,
   R => '0',
   Q => W_reg_20_14
);
W_reg_20_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x113_out_15,
   R => '0',
   Q => W_reg_20_15
);
W_reg_20_15_i_1 : CARRY4
 port map (
   CI => W_reg_20_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_20_15_i_5_n_0,
   DI(1) => W_20_15_i_4_n_0,
   DI(2) => W_20_15_i_3_n_0,
   DI(3) => W_20_15_i_2_n_0,
   S(0) => W_20_15_i_9_n_0,
   S(1) => W_20_15_i_8_n_0,
   S(2) => W_20_15_i_7_n_0,
   S(3) => W_20_15_i_6_n_0,
   CO(0) => W_reg_20_15_i_1_n_3,
   CO(1) => W_reg_20_15_i_1_n_2,
   CO(2) => W_reg_20_15_i_1_n_1,
   CO(3) => W_reg_20_15_i_1_n_0,
   O(0) => x113_out_12,
   O(1) => x113_out_13,
   O(2) => x113_out_14,
   O(3) => x113_out_15
);
W_reg_20_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x113_out_16,
   R => '0',
   Q => W_reg_20_16
);
W_reg_20_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x113_out_17,
   R => '0',
   Q => W_reg_20_17
);
W_reg_20_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x113_out_18,
   R => '0',
   Q => W_reg_20_18
);
W_reg_20_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x113_out_19,
   R => '0',
   Q => W_reg_20_19
);
W_reg_20_19_i_1 : CARRY4
 port map (
   CI => W_reg_20_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_20_19_i_5_n_0,
   DI(1) => W_20_19_i_4_n_0,
   DI(2) => W_20_19_i_3_n_0,
   DI(3) => W_20_19_i_2_n_0,
   S(0) => W_20_19_i_9_n_0,
   S(1) => W_20_19_i_8_n_0,
   S(2) => W_20_19_i_7_n_0,
   S(3) => W_20_19_i_6_n_0,
   CO(0) => W_reg_20_19_i_1_n_3,
   CO(1) => W_reg_20_19_i_1_n_2,
   CO(2) => W_reg_20_19_i_1_n_1,
   CO(3) => W_reg_20_19_i_1_n_0,
   O(0) => x113_out_16,
   O(1) => x113_out_17,
   O(2) => x113_out_18,
   O(3) => x113_out_19
);
W_reg_20_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x113_out_1,
   R => '0',
   Q => W_reg_20_1
);
W_reg_20_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x113_out_20,
   R => '0',
   Q => W_reg_20_20
);
W_reg_20_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x113_out_21,
   R => '0',
   Q => W_reg_20_21
);
W_reg_20_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x113_out_22,
   R => '0',
   Q => W_reg_20_22
);
W_reg_20_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x113_out_23,
   R => '0',
   Q => W_reg_20_23
);
W_reg_20_23_i_1 : CARRY4
 port map (
   CI => W_reg_20_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_20_23_i_5_n_0,
   DI(1) => W_20_23_i_4_n_0,
   DI(2) => W_20_23_i_3_n_0,
   DI(3) => W_20_23_i_2_n_0,
   S(0) => W_20_23_i_9_n_0,
   S(1) => W_20_23_i_8_n_0,
   S(2) => W_20_23_i_7_n_0,
   S(3) => W_20_23_i_6_n_0,
   CO(0) => W_reg_20_23_i_1_n_3,
   CO(1) => W_reg_20_23_i_1_n_2,
   CO(2) => W_reg_20_23_i_1_n_1,
   CO(3) => W_reg_20_23_i_1_n_0,
   O(0) => x113_out_20,
   O(1) => x113_out_21,
   O(2) => x113_out_22,
   O(3) => x113_out_23
);
W_reg_20_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x113_out_24,
   R => '0',
   Q => W_reg_20_24
);
W_reg_20_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x113_out_25,
   R => '0',
   Q => W_reg_20_25
);
W_reg_20_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x113_out_26,
   R => '0',
   Q => W_reg_20_26
);
W_reg_20_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x113_out_27,
   R => '0',
   Q => W_reg_20_27
);
W_reg_20_27_i_1 : CARRY4
 port map (
   CI => W_reg_20_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_20_27_i_5_n_0,
   DI(1) => W_20_27_i_4_n_0,
   DI(2) => W_20_27_i_3_n_0,
   DI(3) => W_20_27_i_2_n_0,
   S(0) => W_20_27_i_9_n_0,
   S(1) => W_20_27_i_8_n_0,
   S(2) => W_20_27_i_7_n_0,
   S(3) => W_20_27_i_6_n_0,
   CO(0) => W_reg_20_27_i_1_n_3,
   CO(1) => W_reg_20_27_i_1_n_2,
   CO(2) => W_reg_20_27_i_1_n_1,
   CO(3) => W_reg_20_27_i_1_n_0,
   O(0) => x113_out_24,
   O(1) => x113_out_25,
   O(2) => x113_out_26,
   O(3) => x113_out_27
);
W_reg_20_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x113_out_28,
   R => '0',
   Q => W_reg_20_28
);
W_reg_20_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x113_out_29,
   R => '0',
   Q => W_reg_20_29
);
W_reg_20_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x113_out_2,
   R => '0',
   Q => W_reg_20_2
);
W_reg_20_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x113_out_30,
   R => '0',
   Q => W_reg_20_30
);
W_reg_20_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x113_out_31,
   R => '0',
   Q => W_reg_20_31
);
W_reg_20_31_i_1 : CARRY4
 port map (
   CI => W_reg_20_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_20_31_i_4_n_0,
   DI(1) => W_20_31_i_3_n_0,
   DI(2) => W_20_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_20_31_i_8_n_0,
   S(1) => W_20_31_i_7_n_0,
   S(2) => W_20_31_i_6_n_0,
   S(3) => W_20_31_i_5_n_0,
   CO(0) => W_reg_20_31_i_1_n_3,
   CO(1) => W_reg_20_31_i_1_n_2,
   CO(2) => W_reg_20_31_i_1_n_1,
   CO(3) => NLW_W_reg_20_31_i_1_CO_UNCONNECTED_3,
   O(0) => x113_out_28,
   O(1) => x113_out_29,
   O(2) => x113_out_30,
   O(3) => x113_out_31
);
W_reg_20_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x113_out_3,
   R => '0',
   Q => W_reg_20_3
);
W_reg_20_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_20_3_i_5_n_0,
   DI(1) => W_20_3_i_4_n_0,
   DI(2) => W_20_3_i_3_n_0,
   DI(3) => W_20_3_i_2_n_0,
   S(0) => W_20_3_i_9_n_0,
   S(1) => W_20_3_i_8_n_0,
   S(2) => W_20_3_i_7_n_0,
   S(3) => W_20_3_i_6_n_0,
   CO(0) => W_reg_20_3_i_1_n_3,
   CO(1) => W_reg_20_3_i_1_n_2,
   CO(2) => W_reg_20_3_i_1_n_1,
   CO(3) => W_reg_20_3_i_1_n_0,
   O(0) => x113_out_0,
   O(1) => x113_out_1,
   O(2) => x113_out_2,
   O(3) => x113_out_3
);
W_reg_20_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x113_out_4,
   R => '0',
   Q => W_reg_20_4
);
W_reg_20_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x113_out_5,
   R => '0',
   Q => W_reg_20_5
);
W_reg_20_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x113_out_6,
   R => '0',
   Q => W_reg_20_6
);
W_reg_20_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x113_out_7,
   R => '0',
   Q => W_reg_20_7
);
W_reg_20_7_i_1 : CARRY4
 port map (
   CI => W_reg_20_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_20_7_i_5_n_0,
   DI(1) => W_20_7_i_4_n_0,
   DI(2) => W_20_7_i_3_n_0,
   DI(3) => W_20_7_i_2_n_0,
   S(0) => W_20_7_i_9_n_0,
   S(1) => W_20_7_i_8_n_0,
   S(2) => W_20_7_i_7_n_0,
   S(3) => W_20_7_i_6_n_0,
   CO(0) => W_reg_20_7_i_1_n_3,
   CO(1) => W_reg_20_7_i_1_n_2,
   CO(2) => W_reg_20_7_i_1_n_1,
   CO(3) => W_reg_20_7_i_1_n_0,
   O(0) => x113_out_4,
   O(1) => x113_out_5,
   O(2) => x113_out_6,
   O(3) => x113_out_7
);
W_reg_20_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x113_out_8,
   R => '0',
   Q => W_reg_20_8
);
W_reg_20_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x113_out_9,
   R => '0',
   Q => W_reg_20_9
);
W_reg_21_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x112_out_0,
   R => '0',
   Q => W_reg_21_0
);
W_reg_21_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x112_out_10,
   R => '0',
   Q => W_reg_21_10
);
W_reg_21_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x112_out_11,
   R => '0',
   Q => W_reg_21_11
);
W_reg_21_11_i_1 : CARRY4
 port map (
   CI => W_reg_21_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_21_11_i_5_n_0,
   DI(1) => W_21_11_i_4_n_0,
   DI(2) => W_21_11_i_3_n_0,
   DI(3) => W_21_11_i_2_n_0,
   S(0) => W_21_11_i_9_n_0,
   S(1) => W_21_11_i_8_n_0,
   S(2) => W_21_11_i_7_n_0,
   S(3) => W_21_11_i_6_n_0,
   CO(0) => W_reg_21_11_i_1_n_3,
   CO(1) => W_reg_21_11_i_1_n_2,
   CO(2) => W_reg_21_11_i_1_n_1,
   CO(3) => W_reg_21_11_i_1_n_0,
   O(0) => x112_out_8,
   O(1) => x112_out_9,
   O(2) => x112_out_10,
   O(3) => x112_out_11
);
W_reg_21_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x112_out_12,
   R => '0',
   Q => W_reg_21_12
);
W_reg_21_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x112_out_13,
   R => '0',
   Q => W_reg_21_13
);
W_reg_21_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x112_out_14,
   R => '0',
   Q => W_reg_21_14
);
W_reg_21_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x112_out_15,
   R => '0',
   Q => W_reg_21_15
);
W_reg_21_15_i_1 : CARRY4
 port map (
   CI => W_reg_21_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_21_15_i_5_n_0,
   DI(1) => W_21_15_i_4_n_0,
   DI(2) => W_21_15_i_3_n_0,
   DI(3) => W_21_15_i_2_n_0,
   S(0) => W_21_15_i_9_n_0,
   S(1) => W_21_15_i_8_n_0,
   S(2) => W_21_15_i_7_n_0,
   S(3) => W_21_15_i_6_n_0,
   CO(0) => W_reg_21_15_i_1_n_3,
   CO(1) => W_reg_21_15_i_1_n_2,
   CO(2) => W_reg_21_15_i_1_n_1,
   CO(3) => W_reg_21_15_i_1_n_0,
   O(0) => x112_out_12,
   O(1) => x112_out_13,
   O(2) => x112_out_14,
   O(3) => x112_out_15
);
W_reg_21_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x112_out_16,
   R => '0',
   Q => W_reg_21_16
);
W_reg_21_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x112_out_17,
   R => '0',
   Q => W_reg_21_17
);
W_reg_21_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x112_out_18,
   R => '0',
   Q => W_reg_21_18
);
W_reg_21_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x112_out_19,
   R => '0',
   Q => W_reg_21_19
);
W_reg_21_19_i_1 : CARRY4
 port map (
   CI => W_reg_21_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_21_19_i_5_n_0,
   DI(1) => W_21_19_i_4_n_0,
   DI(2) => W_21_19_i_3_n_0,
   DI(3) => W_21_19_i_2_n_0,
   S(0) => W_21_19_i_9_n_0,
   S(1) => W_21_19_i_8_n_0,
   S(2) => W_21_19_i_7_n_0,
   S(3) => W_21_19_i_6_n_0,
   CO(0) => W_reg_21_19_i_1_n_3,
   CO(1) => W_reg_21_19_i_1_n_2,
   CO(2) => W_reg_21_19_i_1_n_1,
   CO(3) => W_reg_21_19_i_1_n_0,
   O(0) => x112_out_16,
   O(1) => x112_out_17,
   O(2) => x112_out_18,
   O(3) => x112_out_19
);
W_reg_21_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x112_out_1,
   R => '0',
   Q => W_reg_21_1
);
W_reg_21_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x112_out_20,
   R => '0',
   Q => W_reg_21_20
);
W_reg_21_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x112_out_21,
   R => '0',
   Q => W_reg_21_21
);
W_reg_21_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x112_out_22,
   R => '0',
   Q => W_reg_21_22
);
W_reg_21_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x112_out_23,
   R => '0',
   Q => W_reg_21_23
);
W_reg_21_23_i_1 : CARRY4
 port map (
   CI => W_reg_21_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_21_23_i_5_n_0,
   DI(1) => W_21_23_i_4_n_0,
   DI(2) => W_21_23_i_3_n_0,
   DI(3) => W_21_23_i_2_n_0,
   S(0) => W_21_23_i_9_n_0,
   S(1) => W_21_23_i_8_n_0,
   S(2) => W_21_23_i_7_n_0,
   S(3) => W_21_23_i_6_n_0,
   CO(0) => W_reg_21_23_i_1_n_3,
   CO(1) => W_reg_21_23_i_1_n_2,
   CO(2) => W_reg_21_23_i_1_n_1,
   CO(3) => W_reg_21_23_i_1_n_0,
   O(0) => x112_out_20,
   O(1) => x112_out_21,
   O(2) => x112_out_22,
   O(3) => x112_out_23
);
W_reg_21_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x112_out_24,
   R => '0',
   Q => W_reg_21_24
);
W_reg_21_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x112_out_25,
   R => '0',
   Q => W_reg_21_25
);
W_reg_21_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x112_out_26,
   R => '0',
   Q => W_reg_21_26
);
W_reg_21_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x112_out_27,
   R => '0',
   Q => W_reg_21_27
);
W_reg_21_27_i_1 : CARRY4
 port map (
   CI => W_reg_21_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_21_27_i_5_n_0,
   DI(1) => W_21_27_i_4_n_0,
   DI(2) => W_21_27_i_3_n_0,
   DI(3) => W_21_27_i_2_n_0,
   S(0) => W_21_27_i_9_n_0,
   S(1) => W_21_27_i_8_n_0,
   S(2) => W_21_27_i_7_n_0,
   S(3) => W_21_27_i_6_n_0,
   CO(0) => W_reg_21_27_i_1_n_3,
   CO(1) => W_reg_21_27_i_1_n_2,
   CO(2) => W_reg_21_27_i_1_n_1,
   CO(3) => W_reg_21_27_i_1_n_0,
   O(0) => x112_out_24,
   O(1) => x112_out_25,
   O(2) => x112_out_26,
   O(3) => x112_out_27
);
W_reg_21_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x112_out_28,
   R => '0',
   Q => W_reg_21_28
);
W_reg_21_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x112_out_29,
   R => '0',
   Q => W_reg_21_29
);
W_reg_21_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x112_out_2,
   R => '0',
   Q => W_reg_21_2
);
W_reg_21_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x112_out_30,
   R => '0',
   Q => W_reg_21_30
);
W_reg_21_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x112_out_31,
   R => '0',
   Q => W_reg_21_31
);
W_reg_21_31_i_1 : CARRY4
 port map (
   CI => W_reg_21_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_21_31_i_4_n_0,
   DI(1) => W_21_31_i_3_n_0,
   DI(2) => W_21_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_21_31_i_8_n_0,
   S(1) => W_21_31_i_7_n_0,
   S(2) => W_21_31_i_6_n_0,
   S(3) => W_21_31_i_5_n_0,
   CO(0) => W_reg_21_31_i_1_n_3,
   CO(1) => W_reg_21_31_i_1_n_2,
   CO(2) => W_reg_21_31_i_1_n_1,
   CO(3) => NLW_W_reg_21_31_i_1_CO_UNCONNECTED_3,
   O(0) => x112_out_28,
   O(1) => x112_out_29,
   O(2) => x112_out_30,
   O(3) => x112_out_31
);
W_reg_21_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x112_out_3,
   R => '0',
   Q => W_reg_21_3
);
W_reg_21_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_21_3_i_5_n_0,
   DI(1) => W_21_3_i_4_n_0,
   DI(2) => W_21_3_i_3_n_0,
   DI(3) => W_21_3_i_2_n_0,
   S(0) => W_21_3_i_9_n_0,
   S(1) => W_21_3_i_8_n_0,
   S(2) => W_21_3_i_7_n_0,
   S(3) => W_21_3_i_6_n_0,
   CO(0) => W_reg_21_3_i_1_n_3,
   CO(1) => W_reg_21_3_i_1_n_2,
   CO(2) => W_reg_21_3_i_1_n_1,
   CO(3) => W_reg_21_3_i_1_n_0,
   O(0) => x112_out_0,
   O(1) => x112_out_1,
   O(2) => x112_out_2,
   O(3) => x112_out_3
);
W_reg_21_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x112_out_4,
   R => '0',
   Q => W_reg_21_4
);
W_reg_21_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x112_out_5,
   R => '0',
   Q => W_reg_21_5
);
W_reg_21_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x112_out_6,
   R => '0',
   Q => W_reg_21_6
);
W_reg_21_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x112_out_7,
   R => '0',
   Q => W_reg_21_7
);
W_reg_21_7_i_1 : CARRY4
 port map (
   CI => W_reg_21_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_21_7_i_5_n_0,
   DI(1) => W_21_7_i_4_n_0,
   DI(2) => W_21_7_i_3_n_0,
   DI(3) => W_21_7_i_2_n_0,
   S(0) => W_21_7_i_9_n_0,
   S(1) => W_21_7_i_8_n_0,
   S(2) => W_21_7_i_7_n_0,
   S(3) => W_21_7_i_6_n_0,
   CO(0) => W_reg_21_7_i_1_n_3,
   CO(1) => W_reg_21_7_i_1_n_2,
   CO(2) => W_reg_21_7_i_1_n_1,
   CO(3) => W_reg_21_7_i_1_n_0,
   O(0) => x112_out_4,
   O(1) => x112_out_5,
   O(2) => x112_out_6,
   O(3) => x112_out_7
);
W_reg_21_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x112_out_8,
   R => '0',
   Q => W_reg_21_8
);
W_reg_21_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x112_out_9,
   R => '0',
   Q => W_reg_21_9
);
W_reg_22_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x111_out_0,
   R => '0',
   Q => W_reg_22_0
);
W_reg_22_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x111_out_10,
   R => '0',
   Q => W_reg_22_10
);
W_reg_22_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x111_out_11,
   R => '0',
   Q => W_reg_22_11
);
W_reg_22_11_i_1 : CARRY4
 port map (
   CI => W_reg_22_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_22_11_i_5_n_0,
   DI(1) => W_22_11_i_4_n_0,
   DI(2) => W_22_11_i_3_n_0,
   DI(3) => W_22_11_i_2_n_0,
   S(0) => W_22_11_i_9_n_0,
   S(1) => W_22_11_i_8_n_0,
   S(2) => W_22_11_i_7_n_0,
   S(3) => W_22_11_i_6_n_0,
   CO(0) => W_reg_22_11_i_1_n_3,
   CO(1) => W_reg_22_11_i_1_n_2,
   CO(2) => W_reg_22_11_i_1_n_1,
   CO(3) => W_reg_22_11_i_1_n_0,
   O(0) => x111_out_8,
   O(1) => x111_out_9,
   O(2) => x111_out_10,
   O(3) => x111_out_11
);
W_reg_22_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x111_out_12,
   R => '0',
   Q => W_reg_22_12
);
W_reg_22_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x111_out_13,
   R => '0',
   Q => W_reg_22_13
);
W_reg_22_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x111_out_14,
   R => '0',
   Q => W_reg_22_14
);
W_reg_22_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x111_out_15,
   R => '0',
   Q => W_reg_22_15
);
W_reg_22_15_i_1 : CARRY4
 port map (
   CI => W_reg_22_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_22_15_i_5_n_0,
   DI(1) => W_22_15_i_4_n_0,
   DI(2) => W_22_15_i_3_n_0,
   DI(3) => W_22_15_i_2_n_0,
   S(0) => W_22_15_i_9_n_0,
   S(1) => W_22_15_i_8_n_0,
   S(2) => W_22_15_i_7_n_0,
   S(3) => W_22_15_i_6_n_0,
   CO(0) => W_reg_22_15_i_1_n_3,
   CO(1) => W_reg_22_15_i_1_n_2,
   CO(2) => W_reg_22_15_i_1_n_1,
   CO(3) => W_reg_22_15_i_1_n_0,
   O(0) => x111_out_12,
   O(1) => x111_out_13,
   O(2) => x111_out_14,
   O(3) => x111_out_15
);
W_reg_22_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x111_out_16,
   R => '0',
   Q => W_reg_22_16
);
W_reg_22_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x111_out_17,
   R => '0',
   Q => W_reg_22_17
);
W_reg_22_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x111_out_18,
   R => '0',
   Q => W_reg_22_18
);
W_reg_22_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x111_out_19,
   R => '0',
   Q => W_reg_22_19
);
W_reg_22_19_i_1 : CARRY4
 port map (
   CI => W_reg_22_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_22_19_i_5_n_0,
   DI(1) => W_22_19_i_4_n_0,
   DI(2) => W_22_19_i_3_n_0,
   DI(3) => W_22_19_i_2_n_0,
   S(0) => W_22_19_i_9_n_0,
   S(1) => W_22_19_i_8_n_0,
   S(2) => W_22_19_i_7_n_0,
   S(3) => W_22_19_i_6_n_0,
   CO(0) => W_reg_22_19_i_1_n_3,
   CO(1) => W_reg_22_19_i_1_n_2,
   CO(2) => W_reg_22_19_i_1_n_1,
   CO(3) => W_reg_22_19_i_1_n_0,
   O(0) => x111_out_16,
   O(1) => x111_out_17,
   O(2) => x111_out_18,
   O(3) => x111_out_19
);
W_reg_22_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x111_out_1,
   R => '0',
   Q => W_reg_22_1
);
W_reg_22_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x111_out_20,
   R => '0',
   Q => W_reg_22_20
);
W_reg_22_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x111_out_21,
   R => '0',
   Q => W_reg_22_21
);
W_reg_22_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x111_out_22,
   R => '0',
   Q => W_reg_22_22
);
W_reg_22_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x111_out_23,
   R => '0',
   Q => W_reg_22_23
);
W_reg_22_23_i_1 : CARRY4
 port map (
   CI => W_reg_22_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_22_23_i_5_n_0,
   DI(1) => W_22_23_i_4_n_0,
   DI(2) => W_22_23_i_3_n_0,
   DI(3) => W_22_23_i_2_n_0,
   S(0) => W_22_23_i_9_n_0,
   S(1) => W_22_23_i_8_n_0,
   S(2) => W_22_23_i_7_n_0,
   S(3) => W_22_23_i_6_n_0,
   CO(0) => W_reg_22_23_i_1_n_3,
   CO(1) => W_reg_22_23_i_1_n_2,
   CO(2) => W_reg_22_23_i_1_n_1,
   CO(3) => W_reg_22_23_i_1_n_0,
   O(0) => x111_out_20,
   O(1) => x111_out_21,
   O(2) => x111_out_22,
   O(3) => x111_out_23
);
W_reg_22_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x111_out_24,
   R => '0',
   Q => W_reg_22_24
);
W_reg_22_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x111_out_25,
   R => '0',
   Q => W_reg_22_25
);
W_reg_22_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x111_out_26,
   R => '0',
   Q => W_reg_22_26
);
W_reg_22_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x111_out_27,
   R => '0',
   Q => W_reg_22_27
);
W_reg_22_27_i_1 : CARRY4
 port map (
   CI => W_reg_22_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_22_27_i_5_n_0,
   DI(1) => W_22_27_i_4_n_0,
   DI(2) => W_22_27_i_3_n_0,
   DI(3) => W_22_27_i_2_n_0,
   S(0) => W_22_27_i_9_n_0,
   S(1) => W_22_27_i_8_n_0,
   S(2) => W_22_27_i_7_n_0,
   S(3) => W_22_27_i_6_n_0,
   CO(0) => W_reg_22_27_i_1_n_3,
   CO(1) => W_reg_22_27_i_1_n_2,
   CO(2) => W_reg_22_27_i_1_n_1,
   CO(3) => W_reg_22_27_i_1_n_0,
   O(0) => x111_out_24,
   O(1) => x111_out_25,
   O(2) => x111_out_26,
   O(3) => x111_out_27
);
W_reg_22_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x111_out_28,
   R => '0',
   Q => W_reg_22_28
);
W_reg_22_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x111_out_29,
   R => '0',
   Q => W_reg_22_29
);
W_reg_22_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x111_out_2,
   R => '0',
   Q => W_reg_22_2
);
W_reg_22_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x111_out_30,
   R => '0',
   Q => W_reg_22_30
);
W_reg_22_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x111_out_31,
   R => '0',
   Q => W_reg_22_31
);
W_reg_22_31_i_1 : CARRY4
 port map (
   CI => W_reg_22_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_22_31_i_4_n_0,
   DI(1) => W_22_31_i_3_n_0,
   DI(2) => W_22_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_22_31_i_8_n_0,
   S(1) => W_22_31_i_7_n_0,
   S(2) => W_22_31_i_6_n_0,
   S(3) => W_22_31_i_5_n_0,
   CO(0) => W_reg_22_31_i_1_n_3,
   CO(1) => W_reg_22_31_i_1_n_2,
   CO(2) => W_reg_22_31_i_1_n_1,
   CO(3) => NLW_W_reg_22_31_i_1_CO_UNCONNECTED_3,
   O(0) => x111_out_28,
   O(1) => x111_out_29,
   O(2) => x111_out_30,
   O(3) => x111_out_31
);
W_reg_22_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x111_out_3,
   R => '0',
   Q => W_reg_22_3
);
W_reg_22_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_22_3_i_5_n_0,
   DI(1) => W_22_3_i_4_n_0,
   DI(2) => W_22_3_i_3_n_0,
   DI(3) => W_22_3_i_2_n_0,
   S(0) => W_22_3_i_9_n_0,
   S(1) => W_22_3_i_8_n_0,
   S(2) => W_22_3_i_7_n_0,
   S(3) => W_22_3_i_6_n_0,
   CO(0) => W_reg_22_3_i_1_n_3,
   CO(1) => W_reg_22_3_i_1_n_2,
   CO(2) => W_reg_22_3_i_1_n_1,
   CO(3) => W_reg_22_3_i_1_n_0,
   O(0) => x111_out_0,
   O(1) => x111_out_1,
   O(2) => x111_out_2,
   O(3) => x111_out_3
);
W_reg_22_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x111_out_4,
   R => '0',
   Q => W_reg_22_4
);
W_reg_22_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x111_out_5,
   R => '0',
   Q => W_reg_22_5
);
W_reg_22_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x111_out_6,
   R => '0',
   Q => W_reg_22_6
);
W_reg_22_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x111_out_7,
   R => '0',
   Q => W_reg_22_7
);
W_reg_22_7_i_1 : CARRY4
 port map (
   CI => W_reg_22_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_22_7_i_5_n_0,
   DI(1) => W_22_7_i_4_n_0,
   DI(2) => W_22_7_i_3_n_0,
   DI(3) => W_22_7_i_2_n_0,
   S(0) => W_22_7_i_9_n_0,
   S(1) => W_22_7_i_8_n_0,
   S(2) => W_22_7_i_7_n_0,
   S(3) => W_22_7_i_6_n_0,
   CO(0) => W_reg_22_7_i_1_n_3,
   CO(1) => W_reg_22_7_i_1_n_2,
   CO(2) => W_reg_22_7_i_1_n_1,
   CO(3) => W_reg_22_7_i_1_n_0,
   O(0) => x111_out_4,
   O(1) => x111_out_5,
   O(2) => x111_out_6,
   O(3) => x111_out_7
);
W_reg_22_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x111_out_8,
   R => '0',
   Q => W_reg_22_8
);
W_reg_22_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x111_out_9,
   R => '0',
   Q => W_reg_22_9
);
W_reg_23_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x110_out_0,
   R => '0',
   Q => W_reg_23_0
);
W_reg_23_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x110_out_10,
   R => '0',
   Q => W_reg_23_10
);
W_reg_23_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x110_out_11,
   R => '0',
   Q => W_reg_23_11
);
W_reg_23_11_i_1 : CARRY4
 port map (
   CI => W_reg_23_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_23_11_i_5_n_0,
   DI(1) => W_23_11_i_4_n_0,
   DI(2) => W_23_11_i_3_n_0,
   DI(3) => W_23_11_i_2_n_0,
   S(0) => W_23_11_i_9_n_0,
   S(1) => W_23_11_i_8_n_0,
   S(2) => W_23_11_i_7_n_0,
   S(3) => W_23_11_i_6_n_0,
   CO(0) => W_reg_23_11_i_1_n_3,
   CO(1) => W_reg_23_11_i_1_n_2,
   CO(2) => W_reg_23_11_i_1_n_1,
   CO(3) => W_reg_23_11_i_1_n_0,
   O(0) => x110_out_8,
   O(1) => x110_out_9,
   O(2) => x110_out_10,
   O(3) => x110_out_11
);
W_reg_23_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x110_out_12,
   R => '0',
   Q => W_reg_23_12
);
W_reg_23_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x110_out_13,
   R => '0',
   Q => W_reg_23_13
);
W_reg_23_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x110_out_14,
   R => '0',
   Q => W_reg_23_14
);
W_reg_23_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x110_out_15,
   R => '0',
   Q => W_reg_23_15
);
W_reg_23_15_i_1 : CARRY4
 port map (
   CI => W_reg_23_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_23_15_i_5_n_0,
   DI(1) => W_23_15_i_4_n_0,
   DI(2) => W_23_15_i_3_n_0,
   DI(3) => W_23_15_i_2_n_0,
   S(0) => W_23_15_i_9_n_0,
   S(1) => W_23_15_i_8_n_0,
   S(2) => W_23_15_i_7_n_0,
   S(3) => W_23_15_i_6_n_0,
   CO(0) => W_reg_23_15_i_1_n_3,
   CO(1) => W_reg_23_15_i_1_n_2,
   CO(2) => W_reg_23_15_i_1_n_1,
   CO(3) => W_reg_23_15_i_1_n_0,
   O(0) => x110_out_12,
   O(1) => x110_out_13,
   O(2) => x110_out_14,
   O(3) => x110_out_15
);
W_reg_23_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x110_out_16,
   R => '0',
   Q => W_reg_23_16
);
W_reg_23_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x110_out_17,
   R => '0',
   Q => W_reg_23_17
);
W_reg_23_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x110_out_18,
   R => '0',
   Q => W_reg_23_18
);
W_reg_23_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x110_out_19,
   R => '0',
   Q => W_reg_23_19
);
W_reg_23_19_i_1 : CARRY4
 port map (
   CI => W_reg_23_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_23_19_i_5_n_0,
   DI(1) => W_23_19_i_4_n_0,
   DI(2) => W_23_19_i_3_n_0,
   DI(3) => W_23_19_i_2_n_0,
   S(0) => W_23_19_i_9_n_0,
   S(1) => W_23_19_i_8_n_0,
   S(2) => W_23_19_i_7_n_0,
   S(3) => W_23_19_i_6_n_0,
   CO(0) => W_reg_23_19_i_1_n_3,
   CO(1) => W_reg_23_19_i_1_n_2,
   CO(2) => W_reg_23_19_i_1_n_1,
   CO(3) => W_reg_23_19_i_1_n_0,
   O(0) => x110_out_16,
   O(1) => x110_out_17,
   O(2) => x110_out_18,
   O(3) => x110_out_19
);
W_reg_23_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x110_out_1,
   R => '0',
   Q => W_reg_23_1
);
W_reg_23_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x110_out_20,
   R => '0',
   Q => W_reg_23_20
);
W_reg_23_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x110_out_21,
   R => '0',
   Q => W_reg_23_21
);
W_reg_23_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x110_out_22,
   R => '0',
   Q => W_reg_23_22
);
W_reg_23_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x110_out_23,
   R => '0',
   Q => W_reg_23_23
);
W_reg_23_23_i_1 : CARRY4
 port map (
   CI => W_reg_23_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_23_23_i_5_n_0,
   DI(1) => W_23_23_i_4_n_0,
   DI(2) => W_23_23_i_3_n_0,
   DI(3) => W_23_23_i_2_n_0,
   S(0) => W_23_23_i_9_n_0,
   S(1) => W_23_23_i_8_n_0,
   S(2) => W_23_23_i_7_n_0,
   S(3) => W_23_23_i_6_n_0,
   CO(0) => W_reg_23_23_i_1_n_3,
   CO(1) => W_reg_23_23_i_1_n_2,
   CO(2) => W_reg_23_23_i_1_n_1,
   CO(3) => W_reg_23_23_i_1_n_0,
   O(0) => x110_out_20,
   O(1) => x110_out_21,
   O(2) => x110_out_22,
   O(3) => x110_out_23
);
W_reg_23_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x110_out_24,
   R => '0',
   Q => W_reg_23_24
);
W_reg_23_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x110_out_25,
   R => '0',
   Q => W_reg_23_25
);
W_reg_23_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x110_out_26,
   R => '0',
   Q => W_reg_23_26
);
W_reg_23_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x110_out_27,
   R => '0',
   Q => W_reg_23_27
);
W_reg_23_27_i_1 : CARRY4
 port map (
   CI => W_reg_23_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_23_27_i_5_n_0,
   DI(1) => W_23_27_i_4_n_0,
   DI(2) => W_23_27_i_3_n_0,
   DI(3) => W_23_27_i_2_n_0,
   S(0) => W_23_27_i_9_n_0,
   S(1) => W_23_27_i_8_n_0,
   S(2) => W_23_27_i_7_n_0,
   S(3) => W_23_27_i_6_n_0,
   CO(0) => W_reg_23_27_i_1_n_3,
   CO(1) => W_reg_23_27_i_1_n_2,
   CO(2) => W_reg_23_27_i_1_n_1,
   CO(3) => W_reg_23_27_i_1_n_0,
   O(0) => x110_out_24,
   O(1) => x110_out_25,
   O(2) => x110_out_26,
   O(3) => x110_out_27
);
W_reg_23_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x110_out_28,
   R => '0',
   Q => W_reg_23_28
);
W_reg_23_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x110_out_29,
   R => '0',
   Q => W_reg_23_29
);
W_reg_23_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x110_out_2,
   R => '0',
   Q => W_reg_23_2
);
W_reg_23_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x110_out_30,
   R => '0',
   Q => W_reg_23_30
);
W_reg_23_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x110_out_31,
   R => '0',
   Q => W_reg_23_31
);
W_reg_23_31_i_1 : CARRY4
 port map (
   CI => W_reg_23_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_23_31_i_4_n_0,
   DI(1) => W_23_31_i_3_n_0,
   DI(2) => W_23_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_23_31_i_8_n_0,
   S(1) => W_23_31_i_7_n_0,
   S(2) => W_23_31_i_6_n_0,
   S(3) => W_23_31_i_5_n_0,
   CO(0) => W_reg_23_31_i_1_n_3,
   CO(1) => W_reg_23_31_i_1_n_2,
   CO(2) => W_reg_23_31_i_1_n_1,
   CO(3) => NLW_W_reg_23_31_i_1_CO_UNCONNECTED_3,
   O(0) => x110_out_28,
   O(1) => x110_out_29,
   O(2) => x110_out_30,
   O(3) => x110_out_31
);
W_reg_23_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x110_out_3,
   R => '0',
   Q => W_reg_23_3
);
W_reg_23_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_23_3_i_5_n_0,
   DI(1) => W_23_3_i_4_n_0,
   DI(2) => W_23_3_i_3_n_0,
   DI(3) => W_23_3_i_2_n_0,
   S(0) => W_23_3_i_9_n_0,
   S(1) => W_23_3_i_8_n_0,
   S(2) => W_23_3_i_7_n_0,
   S(3) => W_23_3_i_6_n_0,
   CO(0) => W_reg_23_3_i_1_n_3,
   CO(1) => W_reg_23_3_i_1_n_2,
   CO(2) => W_reg_23_3_i_1_n_1,
   CO(3) => W_reg_23_3_i_1_n_0,
   O(0) => x110_out_0,
   O(1) => x110_out_1,
   O(2) => x110_out_2,
   O(3) => x110_out_3
);
W_reg_23_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x110_out_4,
   R => '0',
   Q => W_reg_23_4
);
W_reg_23_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x110_out_5,
   R => '0',
   Q => W_reg_23_5
);
W_reg_23_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x110_out_6,
   R => '0',
   Q => W_reg_23_6
);
W_reg_23_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x110_out_7,
   R => '0',
   Q => W_reg_23_7
);
W_reg_23_7_i_1 : CARRY4
 port map (
   CI => W_reg_23_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_23_7_i_5_n_0,
   DI(1) => W_23_7_i_4_n_0,
   DI(2) => W_23_7_i_3_n_0,
   DI(3) => W_23_7_i_2_n_0,
   S(0) => W_23_7_i_9_n_0,
   S(1) => W_23_7_i_8_n_0,
   S(2) => W_23_7_i_7_n_0,
   S(3) => W_23_7_i_6_n_0,
   CO(0) => W_reg_23_7_i_1_n_3,
   CO(1) => W_reg_23_7_i_1_n_2,
   CO(2) => W_reg_23_7_i_1_n_1,
   CO(3) => W_reg_23_7_i_1_n_0,
   O(0) => x110_out_4,
   O(1) => x110_out_5,
   O(2) => x110_out_6,
   O(3) => x110_out_7
);
W_reg_23_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x110_out_8,
   R => '0',
   Q => W_reg_23_8
);
W_reg_23_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x110_out_9,
   R => '0',
   Q => W_reg_23_9
);
W_reg_24_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x108_out_0,
   R => '0',
   Q => W_reg_24_0
);
W_reg_24_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x108_out_10,
   R => '0',
   Q => W_reg_24_10
);
W_reg_24_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x108_out_11,
   R => '0',
   Q => W_reg_24_11
);
W_reg_24_11_i_1 : CARRY4
 port map (
   CI => W_reg_24_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_24_11_i_5_n_0,
   DI(1) => W_24_11_i_4_n_0,
   DI(2) => W_24_11_i_3_n_0,
   DI(3) => W_24_11_i_2_n_0,
   S(0) => W_24_11_i_9_n_0,
   S(1) => W_24_11_i_8_n_0,
   S(2) => W_24_11_i_7_n_0,
   S(3) => W_24_11_i_6_n_0,
   CO(0) => W_reg_24_11_i_1_n_3,
   CO(1) => W_reg_24_11_i_1_n_2,
   CO(2) => W_reg_24_11_i_1_n_1,
   CO(3) => W_reg_24_11_i_1_n_0,
   O(0) => x108_out_8,
   O(1) => x108_out_9,
   O(2) => x108_out_10,
   O(3) => x108_out_11
);
W_reg_24_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x108_out_12,
   R => '0',
   Q => W_reg_24_12
);
W_reg_24_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x108_out_13,
   R => '0',
   Q => W_reg_24_13
);
W_reg_24_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x108_out_14,
   R => '0',
   Q => W_reg_24_14
);
W_reg_24_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x108_out_15,
   R => '0',
   Q => W_reg_24_15
);
W_reg_24_15_i_1 : CARRY4
 port map (
   CI => W_reg_24_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_24_15_i_5_n_0,
   DI(1) => W_24_15_i_4_n_0,
   DI(2) => W_24_15_i_3_n_0,
   DI(3) => W_24_15_i_2_n_0,
   S(0) => W_24_15_i_9_n_0,
   S(1) => W_24_15_i_8_n_0,
   S(2) => W_24_15_i_7_n_0,
   S(3) => W_24_15_i_6_n_0,
   CO(0) => W_reg_24_15_i_1_n_3,
   CO(1) => W_reg_24_15_i_1_n_2,
   CO(2) => W_reg_24_15_i_1_n_1,
   CO(3) => W_reg_24_15_i_1_n_0,
   O(0) => x108_out_12,
   O(1) => x108_out_13,
   O(2) => x108_out_14,
   O(3) => x108_out_15
);
W_reg_24_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x108_out_16,
   R => '0',
   Q => W_reg_24_16
);
W_reg_24_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x108_out_17,
   R => '0',
   Q => W_reg_24_17
);
W_reg_24_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x108_out_18,
   R => '0',
   Q => W_reg_24_18
);
W_reg_24_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x108_out_19,
   R => '0',
   Q => W_reg_24_19
);
W_reg_24_19_i_1 : CARRY4
 port map (
   CI => W_reg_24_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_24_19_i_5_n_0,
   DI(1) => W_24_19_i_4_n_0,
   DI(2) => W_24_19_i_3_n_0,
   DI(3) => W_24_19_i_2_n_0,
   S(0) => W_24_19_i_9_n_0,
   S(1) => W_24_19_i_8_n_0,
   S(2) => W_24_19_i_7_n_0,
   S(3) => W_24_19_i_6_n_0,
   CO(0) => W_reg_24_19_i_1_n_3,
   CO(1) => W_reg_24_19_i_1_n_2,
   CO(2) => W_reg_24_19_i_1_n_1,
   CO(3) => W_reg_24_19_i_1_n_0,
   O(0) => x108_out_16,
   O(1) => x108_out_17,
   O(2) => x108_out_18,
   O(3) => x108_out_19
);
W_reg_24_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x108_out_1,
   R => '0',
   Q => W_reg_24_1
);
W_reg_24_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x108_out_20,
   R => '0',
   Q => W_reg_24_20
);
W_reg_24_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x108_out_21,
   R => '0',
   Q => W_reg_24_21
);
W_reg_24_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x108_out_22,
   R => '0',
   Q => W_reg_24_22
);
W_reg_24_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x108_out_23,
   R => '0',
   Q => W_reg_24_23
);
W_reg_24_23_i_1 : CARRY4
 port map (
   CI => W_reg_24_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_24_23_i_5_n_0,
   DI(1) => W_24_23_i_4_n_0,
   DI(2) => W_24_23_i_3_n_0,
   DI(3) => W_24_23_i_2_n_0,
   S(0) => W_24_23_i_9_n_0,
   S(1) => W_24_23_i_8_n_0,
   S(2) => W_24_23_i_7_n_0,
   S(3) => W_24_23_i_6_n_0,
   CO(0) => W_reg_24_23_i_1_n_3,
   CO(1) => W_reg_24_23_i_1_n_2,
   CO(2) => W_reg_24_23_i_1_n_1,
   CO(3) => W_reg_24_23_i_1_n_0,
   O(0) => x108_out_20,
   O(1) => x108_out_21,
   O(2) => x108_out_22,
   O(3) => x108_out_23
);
W_reg_24_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x108_out_24,
   R => '0',
   Q => W_reg_24_24
);
W_reg_24_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x108_out_25,
   R => '0',
   Q => W_reg_24_25
);
W_reg_24_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x108_out_26,
   R => '0',
   Q => W_reg_24_26
);
W_reg_24_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x108_out_27,
   R => '0',
   Q => W_reg_24_27
);
W_reg_24_27_i_1 : CARRY4
 port map (
   CI => W_reg_24_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_24_27_i_5_n_0,
   DI(1) => W_24_27_i_4_n_0,
   DI(2) => W_24_27_i_3_n_0,
   DI(3) => W_24_27_i_2_n_0,
   S(0) => W_24_27_i_9_n_0,
   S(1) => W_24_27_i_8_n_0,
   S(2) => W_24_27_i_7_n_0,
   S(3) => W_24_27_i_6_n_0,
   CO(0) => W_reg_24_27_i_1_n_3,
   CO(1) => W_reg_24_27_i_1_n_2,
   CO(2) => W_reg_24_27_i_1_n_1,
   CO(3) => W_reg_24_27_i_1_n_0,
   O(0) => x108_out_24,
   O(1) => x108_out_25,
   O(2) => x108_out_26,
   O(3) => x108_out_27
);
W_reg_24_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x108_out_28,
   R => '0',
   Q => W_reg_24_28
);
W_reg_24_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x108_out_29,
   R => '0',
   Q => W_reg_24_29
);
W_reg_24_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x108_out_2,
   R => '0',
   Q => W_reg_24_2
);
W_reg_24_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x108_out_30,
   R => '0',
   Q => W_reg_24_30
);
W_reg_24_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x108_out_31,
   R => '0',
   Q => W_reg_24_31
);
W_reg_24_31_i_1 : CARRY4
 port map (
   CI => W_reg_24_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_24_31_i_4_n_0,
   DI(1) => W_24_31_i_3_n_0,
   DI(2) => W_24_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_24_31_i_8_n_0,
   S(1) => W_24_31_i_7_n_0,
   S(2) => W_24_31_i_6_n_0,
   S(3) => W_24_31_i_5_n_0,
   CO(0) => W_reg_24_31_i_1_n_3,
   CO(1) => W_reg_24_31_i_1_n_2,
   CO(2) => W_reg_24_31_i_1_n_1,
   CO(3) => NLW_W_reg_24_31_i_1_CO_UNCONNECTED_3,
   O(0) => x108_out_28,
   O(1) => x108_out_29,
   O(2) => x108_out_30,
   O(3) => x108_out_31
);
W_reg_24_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x108_out_3,
   R => '0',
   Q => W_reg_24_3
);
W_reg_24_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_24_3_i_5_n_0,
   DI(1) => W_24_3_i_4_n_0,
   DI(2) => W_24_3_i_3_n_0,
   DI(3) => W_24_3_i_2_n_0,
   S(0) => W_24_3_i_9_n_0,
   S(1) => W_24_3_i_8_n_0,
   S(2) => W_24_3_i_7_n_0,
   S(3) => W_24_3_i_6_n_0,
   CO(0) => W_reg_24_3_i_1_n_3,
   CO(1) => W_reg_24_3_i_1_n_2,
   CO(2) => W_reg_24_3_i_1_n_1,
   CO(3) => W_reg_24_3_i_1_n_0,
   O(0) => x108_out_0,
   O(1) => x108_out_1,
   O(2) => x108_out_2,
   O(3) => x108_out_3
);
W_reg_24_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x108_out_4,
   R => '0',
   Q => W_reg_24_4
);
W_reg_24_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x108_out_5,
   R => '0',
   Q => W_reg_24_5
);
W_reg_24_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x108_out_6,
   R => '0',
   Q => W_reg_24_6
);
W_reg_24_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x108_out_7,
   R => '0',
   Q => W_reg_24_7
);
W_reg_24_7_i_1 : CARRY4
 port map (
   CI => W_reg_24_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_24_7_i_5_n_0,
   DI(1) => W_24_7_i_4_n_0,
   DI(2) => W_24_7_i_3_n_0,
   DI(3) => W_24_7_i_2_n_0,
   S(0) => W_24_7_i_9_n_0,
   S(1) => W_24_7_i_8_n_0,
   S(2) => W_24_7_i_7_n_0,
   S(3) => W_24_7_i_6_n_0,
   CO(0) => W_reg_24_7_i_1_n_3,
   CO(1) => W_reg_24_7_i_1_n_2,
   CO(2) => W_reg_24_7_i_1_n_1,
   CO(3) => W_reg_24_7_i_1_n_0,
   O(0) => x108_out_4,
   O(1) => x108_out_5,
   O(2) => x108_out_6,
   O(3) => x108_out_7
);
W_reg_24_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x108_out_8,
   R => '0',
   Q => W_reg_24_8
);
W_reg_24_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x108_out_9,
   R => '0',
   Q => W_reg_24_9
);
W_reg_25_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x106_out_0,
   R => '0',
   Q => W_reg_25_0
);
W_reg_25_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x106_out_10,
   R => '0',
   Q => W_reg_25_10
);
W_reg_25_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x106_out_11,
   R => '0',
   Q => W_reg_25_11
);
W_reg_25_11_i_1 : CARRY4
 port map (
   CI => W_reg_25_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_25_11_i_5_n_0,
   DI(1) => W_25_11_i_4_n_0,
   DI(2) => W_25_11_i_3_n_0,
   DI(3) => W_25_11_i_2_n_0,
   S(0) => W_25_11_i_9_n_0,
   S(1) => W_25_11_i_8_n_0,
   S(2) => W_25_11_i_7_n_0,
   S(3) => W_25_11_i_6_n_0,
   CO(0) => W_reg_25_11_i_1_n_3,
   CO(1) => W_reg_25_11_i_1_n_2,
   CO(2) => W_reg_25_11_i_1_n_1,
   CO(3) => W_reg_25_11_i_1_n_0,
   O(0) => x106_out_8,
   O(1) => x106_out_9,
   O(2) => x106_out_10,
   O(3) => x106_out_11
);
W_reg_25_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x106_out_12,
   R => '0',
   Q => W_reg_25_12
);
W_reg_25_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x106_out_13,
   R => '0',
   Q => W_reg_25_13
);
W_reg_25_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x106_out_14,
   R => '0',
   Q => W_reg_25_14
);
W_reg_25_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x106_out_15,
   R => '0',
   Q => W_reg_25_15
);
W_reg_25_15_i_1 : CARRY4
 port map (
   CI => W_reg_25_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_25_15_i_5_n_0,
   DI(1) => W_25_15_i_4_n_0,
   DI(2) => W_25_15_i_3_n_0,
   DI(3) => W_25_15_i_2_n_0,
   S(0) => W_25_15_i_9_n_0,
   S(1) => W_25_15_i_8_n_0,
   S(2) => W_25_15_i_7_n_0,
   S(3) => W_25_15_i_6_n_0,
   CO(0) => W_reg_25_15_i_1_n_3,
   CO(1) => W_reg_25_15_i_1_n_2,
   CO(2) => W_reg_25_15_i_1_n_1,
   CO(3) => W_reg_25_15_i_1_n_0,
   O(0) => x106_out_12,
   O(1) => x106_out_13,
   O(2) => x106_out_14,
   O(3) => x106_out_15
);
W_reg_25_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x106_out_16,
   R => '0',
   Q => W_reg_25_16
);
W_reg_25_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x106_out_17,
   R => '0',
   Q => W_reg_25_17
);
W_reg_25_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x106_out_18,
   R => '0',
   Q => W_reg_25_18
);
W_reg_25_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x106_out_19,
   R => '0',
   Q => W_reg_25_19
);
W_reg_25_19_i_1 : CARRY4
 port map (
   CI => W_reg_25_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_25_19_i_5_n_0,
   DI(1) => W_25_19_i_4_n_0,
   DI(2) => W_25_19_i_3_n_0,
   DI(3) => W_25_19_i_2_n_0,
   S(0) => W_25_19_i_9_n_0,
   S(1) => W_25_19_i_8_n_0,
   S(2) => W_25_19_i_7_n_0,
   S(3) => W_25_19_i_6_n_0,
   CO(0) => W_reg_25_19_i_1_n_3,
   CO(1) => W_reg_25_19_i_1_n_2,
   CO(2) => W_reg_25_19_i_1_n_1,
   CO(3) => W_reg_25_19_i_1_n_0,
   O(0) => x106_out_16,
   O(1) => x106_out_17,
   O(2) => x106_out_18,
   O(3) => x106_out_19
);
W_reg_25_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x106_out_1,
   R => '0',
   Q => W_reg_25_1
);
W_reg_25_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x106_out_20,
   R => '0',
   Q => W_reg_25_20
);
W_reg_25_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x106_out_21,
   R => '0',
   Q => W_reg_25_21
);
W_reg_25_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x106_out_22,
   R => '0',
   Q => W_reg_25_22
);
W_reg_25_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x106_out_23,
   R => '0',
   Q => W_reg_25_23
);
W_reg_25_23_i_1 : CARRY4
 port map (
   CI => W_reg_25_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_25_23_i_5_n_0,
   DI(1) => W_25_23_i_4_n_0,
   DI(2) => W_25_23_i_3_n_0,
   DI(3) => W_25_23_i_2_n_0,
   S(0) => W_25_23_i_9_n_0,
   S(1) => W_25_23_i_8_n_0,
   S(2) => W_25_23_i_7_n_0,
   S(3) => W_25_23_i_6_n_0,
   CO(0) => W_reg_25_23_i_1_n_3,
   CO(1) => W_reg_25_23_i_1_n_2,
   CO(2) => W_reg_25_23_i_1_n_1,
   CO(3) => W_reg_25_23_i_1_n_0,
   O(0) => x106_out_20,
   O(1) => x106_out_21,
   O(2) => x106_out_22,
   O(3) => x106_out_23
);
W_reg_25_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x106_out_24,
   R => '0',
   Q => W_reg_25_24
);
W_reg_25_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x106_out_25,
   R => '0',
   Q => W_reg_25_25
);
W_reg_25_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x106_out_26,
   R => '0',
   Q => W_reg_25_26
);
W_reg_25_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x106_out_27,
   R => '0',
   Q => W_reg_25_27
);
W_reg_25_27_i_1 : CARRY4
 port map (
   CI => W_reg_25_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_25_27_i_5_n_0,
   DI(1) => W_25_27_i_4_n_0,
   DI(2) => W_25_27_i_3_n_0,
   DI(3) => W_25_27_i_2_n_0,
   S(0) => W_25_27_i_9_n_0,
   S(1) => W_25_27_i_8_n_0,
   S(2) => W_25_27_i_7_n_0,
   S(3) => W_25_27_i_6_n_0,
   CO(0) => W_reg_25_27_i_1_n_3,
   CO(1) => W_reg_25_27_i_1_n_2,
   CO(2) => W_reg_25_27_i_1_n_1,
   CO(3) => W_reg_25_27_i_1_n_0,
   O(0) => x106_out_24,
   O(1) => x106_out_25,
   O(2) => x106_out_26,
   O(3) => x106_out_27
);
W_reg_25_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x106_out_28,
   R => '0',
   Q => W_reg_25_28
);
W_reg_25_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x106_out_29,
   R => '0',
   Q => W_reg_25_29
);
W_reg_25_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x106_out_2,
   R => '0',
   Q => W_reg_25_2
);
W_reg_25_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x106_out_30,
   R => '0',
   Q => W_reg_25_30
);
W_reg_25_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x106_out_31,
   R => '0',
   Q => W_reg_25_31
);
W_reg_25_31_i_1 : CARRY4
 port map (
   CI => W_reg_25_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_25_31_i_4_n_0,
   DI(1) => W_25_31_i_3_n_0,
   DI(2) => W_25_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_25_31_i_8_n_0,
   S(1) => W_25_31_i_7_n_0,
   S(2) => W_25_31_i_6_n_0,
   S(3) => W_25_31_i_5_n_0,
   CO(0) => W_reg_25_31_i_1_n_3,
   CO(1) => W_reg_25_31_i_1_n_2,
   CO(2) => W_reg_25_31_i_1_n_1,
   CO(3) => NLW_W_reg_25_31_i_1_CO_UNCONNECTED_3,
   O(0) => x106_out_28,
   O(1) => x106_out_29,
   O(2) => x106_out_30,
   O(3) => x106_out_31
);
W_reg_25_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x106_out_3,
   R => '0',
   Q => W_reg_25_3
);
W_reg_25_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_25_3_i_5_n_0,
   DI(1) => W_25_3_i_4_n_0,
   DI(2) => W_25_3_i_3_n_0,
   DI(3) => W_25_3_i_2_n_0,
   S(0) => W_25_3_i_9_n_0,
   S(1) => W_25_3_i_8_n_0,
   S(2) => W_25_3_i_7_n_0,
   S(3) => W_25_3_i_6_n_0,
   CO(0) => W_reg_25_3_i_1_n_3,
   CO(1) => W_reg_25_3_i_1_n_2,
   CO(2) => W_reg_25_3_i_1_n_1,
   CO(3) => W_reg_25_3_i_1_n_0,
   O(0) => x106_out_0,
   O(1) => x106_out_1,
   O(2) => x106_out_2,
   O(3) => x106_out_3
);
W_reg_25_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x106_out_4,
   R => '0',
   Q => W_reg_25_4
);
W_reg_25_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x106_out_5,
   R => '0',
   Q => W_reg_25_5
);
W_reg_25_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x106_out_6,
   R => '0',
   Q => W_reg_25_6
);
W_reg_25_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x106_out_7,
   R => '0',
   Q => W_reg_25_7
);
W_reg_25_7_i_1 : CARRY4
 port map (
   CI => W_reg_25_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_25_7_i_5_n_0,
   DI(1) => W_25_7_i_4_n_0,
   DI(2) => W_25_7_i_3_n_0,
   DI(3) => W_25_7_i_2_n_0,
   S(0) => W_25_7_i_9_n_0,
   S(1) => W_25_7_i_8_n_0,
   S(2) => W_25_7_i_7_n_0,
   S(3) => W_25_7_i_6_n_0,
   CO(0) => W_reg_25_7_i_1_n_3,
   CO(1) => W_reg_25_7_i_1_n_2,
   CO(2) => W_reg_25_7_i_1_n_1,
   CO(3) => W_reg_25_7_i_1_n_0,
   O(0) => x106_out_4,
   O(1) => x106_out_5,
   O(2) => x106_out_6,
   O(3) => x106_out_7
);
W_reg_25_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x106_out_8,
   R => '0',
   Q => W_reg_25_8
);
W_reg_25_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x106_out_9,
   R => '0',
   Q => W_reg_25_9
);
W_reg_26_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x104_out_0,
   R => '0',
   Q => W_reg_26_0
);
W_reg_26_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x104_out_10,
   R => '0',
   Q => W_reg_26_10
);
W_reg_26_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x104_out_11,
   R => '0',
   Q => W_reg_26_11
);
W_reg_26_11_i_1 : CARRY4
 port map (
   CI => W_reg_26_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_26_11_i_5_n_0,
   DI(1) => W_26_11_i_4_n_0,
   DI(2) => W_26_11_i_3_n_0,
   DI(3) => W_26_11_i_2_n_0,
   S(0) => W_26_11_i_9_n_0,
   S(1) => W_26_11_i_8_n_0,
   S(2) => W_26_11_i_7_n_0,
   S(3) => W_26_11_i_6_n_0,
   CO(0) => W_reg_26_11_i_1_n_3,
   CO(1) => W_reg_26_11_i_1_n_2,
   CO(2) => W_reg_26_11_i_1_n_1,
   CO(3) => W_reg_26_11_i_1_n_0,
   O(0) => x104_out_8,
   O(1) => x104_out_9,
   O(2) => x104_out_10,
   O(3) => x104_out_11
);
W_reg_26_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x104_out_12,
   R => '0',
   Q => W_reg_26_12
);
W_reg_26_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x104_out_13,
   R => '0',
   Q => W_reg_26_13
);
W_reg_26_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x104_out_14,
   R => '0',
   Q => W_reg_26_14
);
W_reg_26_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x104_out_15,
   R => '0',
   Q => W_reg_26_15
);
W_reg_26_15_i_1 : CARRY4
 port map (
   CI => W_reg_26_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_26_15_i_5_n_0,
   DI(1) => W_26_15_i_4_n_0,
   DI(2) => W_26_15_i_3_n_0,
   DI(3) => W_26_15_i_2_n_0,
   S(0) => W_26_15_i_9_n_0,
   S(1) => W_26_15_i_8_n_0,
   S(2) => W_26_15_i_7_n_0,
   S(3) => W_26_15_i_6_n_0,
   CO(0) => W_reg_26_15_i_1_n_3,
   CO(1) => W_reg_26_15_i_1_n_2,
   CO(2) => W_reg_26_15_i_1_n_1,
   CO(3) => W_reg_26_15_i_1_n_0,
   O(0) => x104_out_12,
   O(1) => x104_out_13,
   O(2) => x104_out_14,
   O(3) => x104_out_15
);
W_reg_26_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x104_out_16,
   R => '0',
   Q => W_reg_26_16
);
W_reg_26_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x104_out_17,
   R => '0',
   Q => W_reg_26_17
);
W_reg_26_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x104_out_18,
   R => '0',
   Q => W_reg_26_18
);
W_reg_26_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x104_out_19,
   R => '0',
   Q => W_reg_26_19
);
W_reg_26_19_i_1 : CARRY4
 port map (
   CI => W_reg_26_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_26_19_i_5_n_0,
   DI(1) => W_26_19_i_4_n_0,
   DI(2) => W_26_19_i_3_n_0,
   DI(3) => W_26_19_i_2_n_0,
   S(0) => W_26_19_i_9_n_0,
   S(1) => W_26_19_i_8_n_0,
   S(2) => W_26_19_i_7_n_0,
   S(3) => W_26_19_i_6_n_0,
   CO(0) => W_reg_26_19_i_1_n_3,
   CO(1) => W_reg_26_19_i_1_n_2,
   CO(2) => W_reg_26_19_i_1_n_1,
   CO(3) => W_reg_26_19_i_1_n_0,
   O(0) => x104_out_16,
   O(1) => x104_out_17,
   O(2) => x104_out_18,
   O(3) => x104_out_19
);
W_reg_26_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x104_out_1,
   R => '0',
   Q => W_reg_26_1
);
W_reg_26_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x104_out_20,
   R => '0',
   Q => W_reg_26_20
);
W_reg_26_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x104_out_21,
   R => '0',
   Q => W_reg_26_21
);
W_reg_26_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x104_out_22,
   R => '0',
   Q => W_reg_26_22
);
W_reg_26_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x104_out_23,
   R => '0',
   Q => W_reg_26_23
);
W_reg_26_23_i_1 : CARRY4
 port map (
   CI => W_reg_26_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_26_23_i_5_n_0,
   DI(1) => W_26_23_i_4_n_0,
   DI(2) => W_26_23_i_3_n_0,
   DI(3) => W_26_23_i_2_n_0,
   S(0) => W_26_23_i_9_n_0,
   S(1) => W_26_23_i_8_n_0,
   S(2) => W_26_23_i_7_n_0,
   S(3) => W_26_23_i_6_n_0,
   CO(0) => W_reg_26_23_i_1_n_3,
   CO(1) => W_reg_26_23_i_1_n_2,
   CO(2) => W_reg_26_23_i_1_n_1,
   CO(3) => W_reg_26_23_i_1_n_0,
   O(0) => x104_out_20,
   O(1) => x104_out_21,
   O(2) => x104_out_22,
   O(3) => x104_out_23
);
W_reg_26_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x104_out_24,
   R => '0',
   Q => W_reg_26_24
);
W_reg_26_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x104_out_25,
   R => '0',
   Q => W_reg_26_25
);
W_reg_26_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x104_out_26,
   R => '0',
   Q => W_reg_26_26
);
W_reg_26_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x104_out_27,
   R => '0',
   Q => W_reg_26_27
);
W_reg_26_27_i_1 : CARRY4
 port map (
   CI => W_reg_26_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_26_27_i_5_n_0,
   DI(1) => W_26_27_i_4_n_0,
   DI(2) => W_26_27_i_3_n_0,
   DI(3) => W_26_27_i_2_n_0,
   S(0) => W_26_27_i_9_n_0,
   S(1) => W_26_27_i_8_n_0,
   S(2) => W_26_27_i_7_n_0,
   S(3) => W_26_27_i_6_n_0,
   CO(0) => W_reg_26_27_i_1_n_3,
   CO(1) => W_reg_26_27_i_1_n_2,
   CO(2) => W_reg_26_27_i_1_n_1,
   CO(3) => W_reg_26_27_i_1_n_0,
   O(0) => x104_out_24,
   O(1) => x104_out_25,
   O(2) => x104_out_26,
   O(3) => x104_out_27
);
W_reg_26_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x104_out_28,
   R => '0',
   Q => W_reg_26_28
);
W_reg_26_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x104_out_29,
   R => '0',
   Q => W_reg_26_29
);
W_reg_26_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x104_out_2,
   R => '0',
   Q => W_reg_26_2
);
W_reg_26_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x104_out_30,
   R => '0',
   Q => W_reg_26_30
);
W_reg_26_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x104_out_31,
   R => '0',
   Q => W_reg_26_31
);
W_reg_26_31_i_1 : CARRY4
 port map (
   CI => W_reg_26_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_26_31_i_4_n_0,
   DI(1) => W_26_31_i_3_n_0,
   DI(2) => W_26_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_26_31_i_8_n_0,
   S(1) => W_26_31_i_7_n_0,
   S(2) => W_26_31_i_6_n_0,
   S(3) => W_26_31_i_5_n_0,
   CO(0) => W_reg_26_31_i_1_n_3,
   CO(1) => W_reg_26_31_i_1_n_2,
   CO(2) => W_reg_26_31_i_1_n_1,
   CO(3) => NLW_W_reg_26_31_i_1_CO_UNCONNECTED_3,
   O(0) => x104_out_28,
   O(1) => x104_out_29,
   O(2) => x104_out_30,
   O(3) => x104_out_31
);
W_reg_26_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x104_out_3,
   R => '0',
   Q => W_reg_26_3
);
W_reg_26_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_26_3_i_5_n_0,
   DI(1) => W_26_3_i_4_n_0,
   DI(2) => W_26_3_i_3_n_0,
   DI(3) => W_26_3_i_2_n_0,
   S(0) => W_26_3_i_9_n_0,
   S(1) => W_26_3_i_8_n_0,
   S(2) => W_26_3_i_7_n_0,
   S(3) => W_26_3_i_6_n_0,
   CO(0) => W_reg_26_3_i_1_n_3,
   CO(1) => W_reg_26_3_i_1_n_2,
   CO(2) => W_reg_26_3_i_1_n_1,
   CO(3) => W_reg_26_3_i_1_n_0,
   O(0) => x104_out_0,
   O(1) => x104_out_1,
   O(2) => x104_out_2,
   O(3) => x104_out_3
);
W_reg_26_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x104_out_4,
   R => '0',
   Q => W_reg_26_4
);
W_reg_26_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x104_out_5,
   R => '0',
   Q => W_reg_26_5
);
W_reg_26_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x104_out_6,
   R => '0',
   Q => W_reg_26_6
);
W_reg_26_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x104_out_7,
   R => '0',
   Q => W_reg_26_7
);
W_reg_26_7_i_1 : CARRY4
 port map (
   CI => W_reg_26_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_26_7_i_5_n_0,
   DI(1) => W_26_7_i_4_n_0,
   DI(2) => W_26_7_i_3_n_0,
   DI(3) => W_26_7_i_2_n_0,
   S(0) => W_26_7_i_9_n_0,
   S(1) => W_26_7_i_8_n_0,
   S(2) => W_26_7_i_7_n_0,
   S(3) => W_26_7_i_6_n_0,
   CO(0) => W_reg_26_7_i_1_n_3,
   CO(1) => W_reg_26_7_i_1_n_2,
   CO(2) => W_reg_26_7_i_1_n_1,
   CO(3) => W_reg_26_7_i_1_n_0,
   O(0) => x104_out_4,
   O(1) => x104_out_5,
   O(2) => x104_out_6,
   O(3) => x104_out_7
);
W_reg_26_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x104_out_8,
   R => '0',
   Q => W_reg_26_8
);
W_reg_26_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x104_out_9,
   R => '0',
   Q => W_reg_26_9
);
W_reg_27_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x102_out_0,
   R => '0',
   Q => W_reg_27_0
);
W_reg_27_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x102_out_10,
   R => '0',
   Q => W_reg_27_10
);
W_reg_27_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x102_out_11,
   R => '0',
   Q => W_reg_27_11
);
W_reg_27_11_i_1 : CARRY4
 port map (
   CI => W_reg_27_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_27_11_i_5_n_0,
   DI(1) => W_27_11_i_4_n_0,
   DI(2) => W_27_11_i_3_n_0,
   DI(3) => W_27_11_i_2_n_0,
   S(0) => W_27_11_i_9_n_0,
   S(1) => W_27_11_i_8_n_0,
   S(2) => W_27_11_i_7_n_0,
   S(3) => W_27_11_i_6_n_0,
   CO(0) => W_reg_27_11_i_1_n_3,
   CO(1) => W_reg_27_11_i_1_n_2,
   CO(2) => W_reg_27_11_i_1_n_1,
   CO(3) => W_reg_27_11_i_1_n_0,
   O(0) => x102_out_8,
   O(1) => x102_out_9,
   O(2) => x102_out_10,
   O(3) => x102_out_11
);
W_reg_27_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x102_out_12,
   R => '0',
   Q => W_reg_27_12
);
W_reg_27_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x102_out_13,
   R => '0',
   Q => W_reg_27_13
);
W_reg_27_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x102_out_14,
   R => '0',
   Q => W_reg_27_14
);
W_reg_27_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x102_out_15,
   R => '0',
   Q => W_reg_27_15
);
W_reg_27_15_i_1 : CARRY4
 port map (
   CI => W_reg_27_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_27_15_i_5_n_0,
   DI(1) => W_27_15_i_4_n_0,
   DI(2) => W_27_15_i_3_n_0,
   DI(3) => W_27_15_i_2_n_0,
   S(0) => W_27_15_i_9_n_0,
   S(1) => W_27_15_i_8_n_0,
   S(2) => W_27_15_i_7_n_0,
   S(3) => W_27_15_i_6_n_0,
   CO(0) => W_reg_27_15_i_1_n_3,
   CO(1) => W_reg_27_15_i_1_n_2,
   CO(2) => W_reg_27_15_i_1_n_1,
   CO(3) => W_reg_27_15_i_1_n_0,
   O(0) => x102_out_12,
   O(1) => x102_out_13,
   O(2) => x102_out_14,
   O(3) => x102_out_15
);
W_reg_27_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x102_out_16,
   R => '0',
   Q => W_reg_27_16
);
W_reg_27_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x102_out_17,
   R => '0',
   Q => W_reg_27_17
);
W_reg_27_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x102_out_18,
   R => '0',
   Q => W_reg_27_18
);
W_reg_27_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x102_out_19,
   R => '0',
   Q => W_reg_27_19
);
W_reg_27_19_i_1 : CARRY4
 port map (
   CI => W_reg_27_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_27_19_i_5_n_0,
   DI(1) => W_27_19_i_4_n_0,
   DI(2) => W_27_19_i_3_n_0,
   DI(3) => W_27_19_i_2_n_0,
   S(0) => W_27_19_i_9_n_0,
   S(1) => W_27_19_i_8_n_0,
   S(2) => W_27_19_i_7_n_0,
   S(3) => W_27_19_i_6_n_0,
   CO(0) => W_reg_27_19_i_1_n_3,
   CO(1) => W_reg_27_19_i_1_n_2,
   CO(2) => W_reg_27_19_i_1_n_1,
   CO(3) => W_reg_27_19_i_1_n_0,
   O(0) => x102_out_16,
   O(1) => x102_out_17,
   O(2) => x102_out_18,
   O(3) => x102_out_19
);
W_reg_27_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x102_out_1,
   R => '0',
   Q => W_reg_27_1
);
W_reg_27_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x102_out_20,
   R => '0',
   Q => W_reg_27_20
);
W_reg_27_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x102_out_21,
   R => '0',
   Q => W_reg_27_21
);
W_reg_27_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x102_out_22,
   R => '0',
   Q => W_reg_27_22
);
W_reg_27_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x102_out_23,
   R => '0',
   Q => W_reg_27_23
);
W_reg_27_23_i_1 : CARRY4
 port map (
   CI => W_reg_27_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_27_23_i_5_n_0,
   DI(1) => W_27_23_i_4_n_0,
   DI(2) => W_27_23_i_3_n_0,
   DI(3) => W_27_23_i_2_n_0,
   S(0) => W_27_23_i_9_n_0,
   S(1) => W_27_23_i_8_n_0,
   S(2) => W_27_23_i_7_n_0,
   S(3) => W_27_23_i_6_n_0,
   CO(0) => W_reg_27_23_i_1_n_3,
   CO(1) => W_reg_27_23_i_1_n_2,
   CO(2) => W_reg_27_23_i_1_n_1,
   CO(3) => W_reg_27_23_i_1_n_0,
   O(0) => x102_out_20,
   O(1) => x102_out_21,
   O(2) => x102_out_22,
   O(3) => x102_out_23
);
W_reg_27_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x102_out_24,
   R => '0',
   Q => W_reg_27_24
);
W_reg_27_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x102_out_25,
   R => '0',
   Q => W_reg_27_25
);
W_reg_27_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x102_out_26,
   R => '0',
   Q => W_reg_27_26
);
W_reg_27_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x102_out_27,
   R => '0',
   Q => W_reg_27_27
);
W_reg_27_27_i_1 : CARRY4
 port map (
   CI => W_reg_27_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_27_27_i_5_n_0,
   DI(1) => W_27_27_i_4_n_0,
   DI(2) => W_27_27_i_3_n_0,
   DI(3) => W_27_27_i_2_n_0,
   S(0) => W_27_27_i_9_n_0,
   S(1) => W_27_27_i_8_n_0,
   S(2) => W_27_27_i_7_n_0,
   S(3) => W_27_27_i_6_n_0,
   CO(0) => W_reg_27_27_i_1_n_3,
   CO(1) => W_reg_27_27_i_1_n_2,
   CO(2) => W_reg_27_27_i_1_n_1,
   CO(3) => W_reg_27_27_i_1_n_0,
   O(0) => x102_out_24,
   O(1) => x102_out_25,
   O(2) => x102_out_26,
   O(3) => x102_out_27
);
W_reg_27_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x102_out_28,
   R => '0',
   Q => W_reg_27_28
);
W_reg_27_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x102_out_29,
   R => '0',
   Q => W_reg_27_29
);
W_reg_27_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x102_out_2,
   R => '0',
   Q => W_reg_27_2
);
W_reg_27_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x102_out_30,
   R => '0',
   Q => W_reg_27_30
);
W_reg_27_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x102_out_31,
   R => '0',
   Q => W_reg_27_31
);
W_reg_27_31_i_1 : CARRY4
 port map (
   CI => W_reg_27_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_27_31_i_4_n_0,
   DI(1) => W_27_31_i_3_n_0,
   DI(2) => W_27_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_27_31_i_8_n_0,
   S(1) => W_27_31_i_7_n_0,
   S(2) => W_27_31_i_6_n_0,
   S(3) => W_27_31_i_5_n_0,
   CO(0) => W_reg_27_31_i_1_n_3,
   CO(1) => W_reg_27_31_i_1_n_2,
   CO(2) => W_reg_27_31_i_1_n_1,
   CO(3) => NLW_W_reg_27_31_i_1_CO_UNCONNECTED_3,
   O(0) => x102_out_28,
   O(1) => x102_out_29,
   O(2) => x102_out_30,
   O(3) => x102_out_31
);
W_reg_27_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x102_out_3,
   R => '0',
   Q => W_reg_27_3
);
W_reg_27_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_27_3_i_5_n_0,
   DI(1) => W_27_3_i_4_n_0,
   DI(2) => W_27_3_i_3_n_0,
   DI(3) => W_27_3_i_2_n_0,
   S(0) => W_27_3_i_9_n_0,
   S(1) => W_27_3_i_8_n_0,
   S(2) => W_27_3_i_7_n_0,
   S(3) => W_27_3_i_6_n_0,
   CO(0) => W_reg_27_3_i_1_n_3,
   CO(1) => W_reg_27_3_i_1_n_2,
   CO(2) => W_reg_27_3_i_1_n_1,
   CO(3) => W_reg_27_3_i_1_n_0,
   O(0) => x102_out_0,
   O(1) => x102_out_1,
   O(2) => x102_out_2,
   O(3) => x102_out_3
);
W_reg_27_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x102_out_4,
   R => '0',
   Q => W_reg_27_4
);
W_reg_27_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x102_out_5,
   R => '0',
   Q => W_reg_27_5
);
W_reg_27_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x102_out_6,
   R => '0',
   Q => W_reg_27_6
);
W_reg_27_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x102_out_7,
   R => '0',
   Q => W_reg_27_7
);
W_reg_27_7_i_1 : CARRY4
 port map (
   CI => W_reg_27_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_27_7_i_5_n_0,
   DI(1) => W_27_7_i_4_n_0,
   DI(2) => W_27_7_i_3_n_0,
   DI(3) => W_27_7_i_2_n_0,
   S(0) => W_27_7_i_9_n_0,
   S(1) => W_27_7_i_8_n_0,
   S(2) => W_27_7_i_7_n_0,
   S(3) => W_27_7_i_6_n_0,
   CO(0) => W_reg_27_7_i_1_n_3,
   CO(1) => W_reg_27_7_i_1_n_2,
   CO(2) => W_reg_27_7_i_1_n_1,
   CO(3) => W_reg_27_7_i_1_n_0,
   O(0) => x102_out_4,
   O(1) => x102_out_5,
   O(2) => x102_out_6,
   O(3) => x102_out_7
);
W_reg_27_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x102_out_8,
   R => '0',
   Q => W_reg_27_8
);
W_reg_27_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x102_out_9,
   R => '0',
   Q => W_reg_27_9
);
W_reg_28_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x100_out_0,
   R => '0',
   Q => W_reg_28_0
);
W_reg_28_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x100_out_10,
   R => '0',
   Q => W_reg_28_10
);
W_reg_28_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x100_out_11,
   R => '0',
   Q => W_reg_28_11
);
W_reg_28_11_i_1 : CARRY4
 port map (
   CI => W_reg_28_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_28_11_i_5_n_0,
   DI(1) => W_28_11_i_4_n_0,
   DI(2) => W_28_11_i_3_n_0,
   DI(3) => W_28_11_i_2_n_0,
   S(0) => W_28_11_i_9_n_0,
   S(1) => W_28_11_i_8_n_0,
   S(2) => W_28_11_i_7_n_0,
   S(3) => W_28_11_i_6_n_0,
   CO(0) => W_reg_28_11_i_1_n_3,
   CO(1) => W_reg_28_11_i_1_n_2,
   CO(2) => W_reg_28_11_i_1_n_1,
   CO(3) => W_reg_28_11_i_1_n_0,
   O(0) => x100_out_8,
   O(1) => x100_out_9,
   O(2) => x100_out_10,
   O(3) => x100_out_11
);
W_reg_28_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x100_out_12,
   R => '0',
   Q => W_reg_28_12
);
W_reg_28_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x100_out_13,
   R => '0',
   Q => W_reg_28_13
);
W_reg_28_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x100_out_14,
   R => '0',
   Q => W_reg_28_14
);
W_reg_28_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x100_out_15,
   R => '0',
   Q => W_reg_28_15
);
W_reg_28_15_i_1 : CARRY4
 port map (
   CI => W_reg_28_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_28_15_i_5_n_0,
   DI(1) => W_28_15_i_4_n_0,
   DI(2) => W_28_15_i_3_n_0,
   DI(3) => W_28_15_i_2_n_0,
   S(0) => W_28_15_i_9_n_0,
   S(1) => W_28_15_i_8_n_0,
   S(2) => W_28_15_i_7_n_0,
   S(3) => W_28_15_i_6_n_0,
   CO(0) => W_reg_28_15_i_1_n_3,
   CO(1) => W_reg_28_15_i_1_n_2,
   CO(2) => W_reg_28_15_i_1_n_1,
   CO(3) => W_reg_28_15_i_1_n_0,
   O(0) => x100_out_12,
   O(1) => x100_out_13,
   O(2) => x100_out_14,
   O(3) => x100_out_15
);
W_reg_28_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x100_out_16,
   R => '0',
   Q => W_reg_28_16
);
W_reg_28_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x100_out_17,
   R => '0',
   Q => W_reg_28_17
);
W_reg_28_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x100_out_18,
   R => '0',
   Q => W_reg_28_18
);
W_reg_28_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x100_out_19,
   R => '0',
   Q => W_reg_28_19
);
W_reg_28_19_i_1 : CARRY4
 port map (
   CI => W_reg_28_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_28_19_i_5_n_0,
   DI(1) => W_28_19_i_4_n_0,
   DI(2) => W_28_19_i_3_n_0,
   DI(3) => W_28_19_i_2_n_0,
   S(0) => W_28_19_i_9_n_0,
   S(1) => W_28_19_i_8_n_0,
   S(2) => W_28_19_i_7_n_0,
   S(3) => W_28_19_i_6_n_0,
   CO(0) => W_reg_28_19_i_1_n_3,
   CO(1) => W_reg_28_19_i_1_n_2,
   CO(2) => W_reg_28_19_i_1_n_1,
   CO(3) => W_reg_28_19_i_1_n_0,
   O(0) => x100_out_16,
   O(1) => x100_out_17,
   O(2) => x100_out_18,
   O(3) => x100_out_19
);
W_reg_28_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x100_out_1,
   R => '0',
   Q => W_reg_28_1
);
W_reg_28_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x100_out_20,
   R => '0',
   Q => W_reg_28_20
);
W_reg_28_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x100_out_21,
   R => '0',
   Q => W_reg_28_21
);
W_reg_28_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x100_out_22,
   R => '0',
   Q => W_reg_28_22
);
W_reg_28_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x100_out_23,
   R => '0',
   Q => W_reg_28_23
);
W_reg_28_23_i_1 : CARRY4
 port map (
   CI => W_reg_28_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_28_23_i_5_n_0,
   DI(1) => W_28_23_i_4_n_0,
   DI(2) => W_28_23_i_3_n_0,
   DI(3) => W_28_23_i_2_n_0,
   S(0) => W_28_23_i_9_n_0,
   S(1) => W_28_23_i_8_n_0,
   S(2) => W_28_23_i_7_n_0,
   S(3) => W_28_23_i_6_n_0,
   CO(0) => W_reg_28_23_i_1_n_3,
   CO(1) => W_reg_28_23_i_1_n_2,
   CO(2) => W_reg_28_23_i_1_n_1,
   CO(3) => W_reg_28_23_i_1_n_0,
   O(0) => x100_out_20,
   O(1) => x100_out_21,
   O(2) => x100_out_22,
   O(3) => x100_out_23
);
W_reg_28_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x100_out_24,
   R => '0',
   Q => W_reg_28_24
);
W_reg_28_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x100_out_25,
   R => '0',
   Q => W_reg_28_25
);
W_reg_28_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x100_out_26,
   R => '0',
   Q => W_reg_28_26
);
W_reg_28_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x100_out_27,
   R => '0',
   Q => W_reg_28_27
);
W_reg_28_27_i_1 : CARRY4
 port map (
   CI => W_reg_28_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_28_27_i_5_n_0,
   DI(1) => W_28_27_i_4_n_0,
   DI(2) => W_28_27_i_3_n_0,
   DI(3) => W_28_27_i_2_n_0,
   S(0) => W_28_27_i_9_n_0,
   S(1) => W_28_27_i_8_n_0,
   S(2) => W_28_27_i_7_n_0,
   S(3) => W_28_27_i_6_n_0,
   CO(0) => W_reg_28_27_i_1_n_3,
   CO(1) => W_reg_28_27_i_1_n_2,
   CO(2) => W_reg_28_27_i_1_n_1,
   CO(3) => W_reg_28_27_i_1_n_0,
   O(0) => x100_out_24,
   O(1) => x100_out_25,
   O(2) => x100_out_26,
   O(3) => x100_out_27
);
W_reg_28_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x100_out_28,
   R => '0',
   Q => W_reg_28_28
);
W_reg_28_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x100_out_29,
   R => '0',
   Q => W_reg_28_29
);
W_reg_28_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x100_out_2,
   R => '0',
   Q => W_reg_28_2
);
W_reg_28_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x100_out_30,
   R => '0',
   Q => W_reg_28_30
);
W_reg_28_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x100_out_31,
   R => '0',
   Q => W_reg_28_31
);
W_reg_28_31_i_1 : CARRY4
 port map (
   CI => W_reg_28_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_28_31_i_4_n_0,
   DI(1) => W_28_31_i_3_n_0,
   DI(2) => W_28_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_28_31_i_8_n_0,
   S(1) => W_28_31_i_7_n_0,
   S(2) => W_28_31_i_6_n_0,
   S(3) => W_28_31_i_5_n_0,
   CO(0) => W_reg_28_31_i_1_n_3,
   CO(1) => W_reg_28_31_i_1_n_2,
   CO(2) => W_reg_28_31_i_1_n_1,
   CO(3) => NLW_W_reg_28_31_i_1_CO_UNCONNECTED_3,
   O(0) => x100_out_28,
   O(1) => x100_out_29,
   O(2) => x100_out_30,
   O(3) => x100_out_31
);
W_reg_28_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x100_out_3,
   R => '0',
   Q => W_reg_28_3
);
W_reg_28_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_28_3_i_5_n_0,
   DI(1) => W_28_3_i_4_n_0,
   DI(2) => W_28_3_i_3_n_0,
   DI(3) => W_28_3_i_2_n_0,
   S(0) => W_28_3_i_9_n_0,
   S(1) => W_28_3_i_8_n_0,
   S(2) => W_28_3_i_7_n_0,
   S(3) => W_28_3_i_6_n_0,
   CO(0) => W_reg_28_3_i_1_n_3,
   CO(1) => W_reg_28_3_i_1_n_2,
   CO(2) => W_reg_28_3_i_1_n_1,
   CO(3) => W_reg_28_3_i_1_n_0,
   O(0) => x100_out_0,
   O(1) => x100_out_1,
   O(2) => x100_out_2,
   O(3) => x100_out_3
);
W_reg_28_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x100_out_4,
   R => '0',
   Q => W_reg_28_4
);
W_reg_28_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x100_out_5,
   R => '0',
   Q => W_reg_28_5
);
W_reg_28_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x100_out_6,
   R => '0',
   Q => W_reg_28_6
);
W_reg_28_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x100_out_7,
   R => '0',
   Q => W_reg_28_7
);
W_reg_28_7_i_1 : CARRY4
 port map (
   CI => W_reg_28_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_28_7_i_5_n_0,
   DI(1) => W_28_7_i_4_n_0,
   DI(2) => W_28_7_i_3_n_0,
   DI(3) => W_28_7_i_2_n_0,
   S(0) => W_28_7_i_9_n_0,
   S(1) => W_28_7_i_8_n_0,
   S(2) => W_28_7_i_7_n_0,
   S(3) => W_28_7_i_6_n_0,
   CO(0) => W_reg_28_7_i_1_n_3,
   CO(1) => W_reg_28_7_i_1_n_2,
   CO(2) => W_reg_28_7_i_1_n_1,
   CO(3) => W_reg_28_7_i_1_n_0,
   O(0) => x100_out_4,
   O(1) => x100_out_5,
   O(2) => x100_out_6,
   O(3) => x100_out_7
);
W_reg_28_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x100_out_8,
   R => '0',
   Q => W_reg_28_8
);
W_reg_28_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x100_out_9,
   R => '0',
   Q => W_reg_28_9
);
W_reg_29_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x98_out_0,
   R => '0',
   Q => W_reg_29_0
);
W_reg_29_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x98_out_10,
   R => '0',
   Q => W_reg_29_10
);
W_reg_29_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x98_out_11,
   R => '0',
   Q => W_reg_29_11
);
W_reg_29_11_i_1 : CARRY4
 port map (
   CI => W_reg_29_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_29_11_i_5_n_0,
   DI(1) => W_29_11_i_4_n_0,
   DI(2) => W_29_11_i_3_n_0,
   DI(3) => W_29_11_i_2_n_0,
   S(0) => W_29_11_i_9_n_0,
   S(1) => W_29_11_i_8_n_0,
   S(2) => W_29_11_i_7_n_0,
   S(3) => W_29_11_i_6_n_0,
   CO(0) => W_reg_29_11_i_1_n_3,
   CO(1) => W_reg_29_11_i_1_n_2,
   CO(2) => W_reg_29_11_i_1_n_1,
   CO(3) => W_reg_29_11_i_1_n_0,
   O(0) => x98_out_8,
   O(1) => x98_out_9,
   O(2) => x98_out_10,
   O(3) => x98_out_11
);
W_reg_29_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x98_out_12,
   R => '0',
   Q => W_reg_29_12
);
W_reg_29_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x98_out_13,
   R => '0',
   Q => W_reg_29_13
);
W_reg_29_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x98_out_14,
   R => '0',
   Q => W_reg_29_14
);
W_reg_29_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x98_out_15,
   R => '0',
   Q => W_reg_29_15
);
W_reg_29_15_i_1 : CARRY4
 port map (
   CI => W_reg_29_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_29_15_i_5_n_0,
   DI(1) => W_29_15_i_4_n_0,
   DI(2) => W_29_15_i_3_n_0,
   DI(3) => W_29_15_i_2_n_0,
   S(0) => W_29_15_i_9_n_0,
   S(1) => W_29_15_i_8_n_0,
   S(2) => W_29_15_i_7_n_0,
   S(3) => W_29_15_i_6_n_0,
   CO(0) => W_reg_29_15_i_1_n_3,
   CO(1) => W_reg_29_15_i_1_n_2,
   CO(2) => W_reg_29_15_i_1_n_1,
   CO(3) => W_reg_29_15_i_1_n_0,
   O(0) => x98_out_12,
   O(1) => x98_out_13,
   O(2) => x98_out_14,
   O(3) => x98_out_15
);
W_reg_29_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x98_out_16,
   R => '0',
   Q => W_reg_29_16
);
W_reg_29_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x98_out_17,
   R => '0',
   Q => W_reg_29_17
);
W_reg_29_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x98_out_18,
   R => '0',
   Q => W_reg_29_18
);
W_reg_29_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x98_out_19,
   R => '0',
   Q => W_reg_29_19
);
W_reg_29_19_i_1 : CARRY4
 port map (
   CI => W_reg_29_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_29_19_i_5_n_0,
   DI(1) => W_29_19_i_4_n_0,
   DI(2) => W_29_19_i_3_n_0,
   DI(3) => W_29_19_i_2_n_0,
   S(0) => W_29_19_i_9_n_0,
   S(1) => W_29_19_i_8_n_0,
   S(2) => W_29_19_i_7_n_0,
   S(3) => W_29_19_i_6_n_0,
   CO(0) => W_reg_29_19_i_1_n_3,
   CO(1) => W_reg_29_19_i_1_n_2,
   CO(2) => W_reg_29_19_i_1_n_1,
   CO(3) => W_reg_29_19_i_1_n_0,
   O(0) => x98_out_16,
   O(1) => x98_out_17,
   O(2) => x98_out_18,
   O(3) => x98_out_19
);
W_reg_29_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x98_out_1,
   R => '0',
   Q => W_reg_29_1
);
W_reg_29_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x98_out_20,
   R => '0',
   Q => W_reg_29_20
);
W_reg_29_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x98_out_21,
   R => '0',
   Q => W_reg_29_21
);
W_reg_29_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x98_out_22,
   R => '0',
   Q => W_reg_29_22
);
W_reg_29_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x98_out_23,
   R => '0',
   Q => W_reg_29_23
);
W_reg_29_23_i_1 : CARRY4
 port map (
   CI => W_reg_29_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_29_23_i_5_n_0,
   DI(1) => W_29_23_i_4_n_0,
   DI(2) => W_29_23_i_3_n_0,
   DI(3) => W_29_23_i_2_n_0,
   S(0) => W_29_23_i_9_n_0,
   S(1) => W_29_23_i_8_n_0,
   S(2) => W_29_23_i_7_n_0,
   S(3) => W_29_23_i_6_n_0,
   CO(0) => W_reg_29_23_i_1_n_3,
   CO(1) => W_reg_29_23_i_1_n_2,
   CO(2) => W_reg_29_23_i_1_n_1,
   CO(3) => W_reg_29_23_i_1_n_0,
   O(0) => x98_out_20,
   O(1) => x98_out_21,
   O(2) => x98_out_22,
   O(3) => x98_out_23
);
W_reg_29_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x98_out_24,
   R => '0',
   Q => W_reg_29_24
);
W_reg_29_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x98_out_25,
   R => '0',
   Q => W_reg_29_25
);
W_reg_29_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x98_out_26,
   R => '0',
   Q => W_reg_29_26
);
W_reg_29_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x98_out_27,
   R => '0',
   Q => W_reg_29_27
);
W_reg_29_27_i_1 : CARRY4
 port map (
   CI => W_reg_29_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_29_27_i_5_n_0,
   DI(1) => W_29_27_i_4_n_0,
   DI(2) => W_29_27_i_3_n_0,
   DI(3) => W_29_27_i_2_n_0,
   S(0) => W_29_27_i_9_n_0,
   S(1) => W_29_27_i_8_n_0,
   S(2) => W_29_27_i_7_n_0,
   S(3) => W_29_27_i_6_n_0,
   CO(0) => W_reg_29_27_i_1_n_3,
   CO(1) => W_reg_29_27_i_1_n_2,
   CO(2) => W_reg_29_27_i_1_n_1,
   CO(3) => W_reg_29_27_i_1_n_0,
   O(0) => x98_out_24,
   O(1) => x98_out_25,
   O(2) => x98_out_26,
   O(3) => x98_out_27
);
W_reg_29_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x98_out_28,
   R => '0',
   Q => W_reg_29_28
);
W_reg_29_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x98_out_29,
   R => '0',
   Q => W_reg_29_29
);
W_reg_29_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x98_out_2,
   R => '0',
   Q => W_reg_29_2
);
W_reg_29_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x98_out_30,
   R => '0',
   Q => W_reg_29_30
);
W_reg_29_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x98_out_31,
   R => '0',
   Q => W_reg_29_31
);
W_reg_29_31_i_1 : CARRY4
 port map (
   CI => W_reg_29_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_29_31_i_4_n_0,
   DI(1) => W_29_31_i_3_n_0,
   DI(2) => W_29_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_29_31_i_8_n_0,
   S(1) => W_29_31_i_7_n_0,
   S(2) => W_29_31_i_6_n_0,
   S(3) => W_29_31_i_5_n_0,
   CO(0) => W_reg_29_31_i_1_n_3,
   CO(1) => W_reg_29_31_i_1_n_2,
   CO(2) => W_reg_29_31_i_1_n_1,
   CO(3) => NLW_W_reg_29_31_i_1_CO_UNCONNECTED_3,
   O(0) => x98_out_28,
   O(1) => x98_out_29,
   O(2) => x98_out_30,
   O(3) => x98_out_31
);
W_reg_29_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x98_out_3,
   R => '0',
   Q => W_reg_29_3
);
W_reg_29_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_29_3_i_5_n_0,
   DI(1) => W_29_3_i_4_n_0,
   DI(2) => W_29_3_i_3_n_0,
   DI(3) => W_29_3_i_2_n_0,
   S(0) => W_29_3_i_9_n_0,
   S(1) => W_29_3_i_8_n_0,
   S(2) => W_29_3_i_7_n_0,
   S(3) => W_29_3_i_6_n_0,
   CO(0) => W_reg_29_3_i_1_n_3,
   CO(1) => W_reg_29_3_i_1_n_2,
   CO(2) => W_reg_29_3_i_1_n_1,
   CO(3) => W_reg_29_3_i_1_n_0,
   O(0) => x98_out_0,
   O(1) => x98_out_1,
   O(2) => x98_out_2,
   O(3) => x98_out_3
);
W_reg_29_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x98_out_4,
   R => '0',
   Q => W_reg_29_4
);
W_reg_29_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x98_out_5,
   R => '0',
   Q => W_reg_29_5
);
W_reg_29_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x98_out_6,
   R => '0',
   Q => W_reg_29_6
);
W_reg_29_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x98_out_7,
   R => '0',
   Q => W_reg_29_7
);
W_reg_29_7_i_1 : CARRY4
 port map (
   CI => W_reg_29_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_29_7_i_5_n_0,
   DI(1) => W_29_7_i_4_n_0,
   DI(2) => W_29_7_i_3_n_0,
   DI(3) => W_29_7_i_2_n_0,
   S(0) => W_29_7_i_9_n_0,
   S(1) => W_29_7_i_8_n_0,
   S(2) => W_29_7_i_7_n_0,
   S(3) => W_29_7_i_6_n_0,
   CO(0) => W_reg_29_7_i_1_n_3,
   CO(1) => W_reg_29_7_i_1_n_2,
   CO(2) => W_reg_29_7_i_1_n_1,
   CO(3) => W_reg_29_7_i_1_n_0,
   O(0) => x98_out_4,
   O(1) => x98_out_5,
   O(2) => x98_out_6,
   O(3) => x98_out_7
);
W_reg_29_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x98_out_8,
   R => '0',
   Q => W_reg_29_8
);
W_reg_29_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x98_out_9,
   R => '0',
   Q => W_reg_29_9
);
W_reg_2_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_2_0,
   R => '0',
   Q => W_reg_2_0
);
W_reg_2_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_2_10,
   R => '0',
   Q => W_reg_2_10
);
W_reg_2_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_2_11,
   R => '0',
   Q => W_reg_2_11
);
W_reg_2_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_2_12,
   R => '0',
   Q => W_reg_2_12
);
W_reg_2_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_2_13,
   R => '0',
   Q => W_reg_2_13
);
W_reg_2_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_2_14,
   R => '0',
   Q => W_reg_2_14
);
W_reg_2_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_2_15,
   R => '0',
   Q => W_reg_2_15
);
W_reg_2_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_2_16,
   R => '0',
   Q => W_reg_2_16
);
W_reg_2_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_2_17,
   R => '0',
   Q => W_reg_2_17
);
W_reg_2_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_2_18,
   R => '0',
   Q => W_reg_2_18
);
W_reg_2_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_2_19,
   R => '0',
   Q => W_reg_2_19
);
W_reg_2_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_2_1,
   R => '0',
   Q => W_reg_2_1
);
W_reg_2_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_2_20,
   R => '0',
   Q => W_reg_2_20
);
W_reg_2_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_2_21,
   R => '0',
   Q => W_reg_2_21
);
W_reg_2_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_2_22,
   R => '0',
   Q => W_reg_2_22
);
W_reg_2_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_2_23,
   R => '0',
   Q => W_reg_2_23
);
W_reg_2_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_2_24,
   R => '0',
   Q => W_reg_2_24
);
W_reg_2_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_2_25,
   R => '0',
   Q => W_reg_2_25
);
W_reg_2_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_2_26,
   R => '0',
   Q => W_reg_2_26
);
W_reg_2_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_2_27,
   R => '0',
   Q => W_reg_2_27
);
W_reg_2_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_2_28,
   R => '0',
   Q => W_reg_2_28
);
W_reg_2_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_2_29,
   R => '0',
   Q => W_reg_2_29
);
W_reg_2_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_2_2,
   R => '0',
   Q => W_reg_2_2
);
W_reg_2_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_2_30,
   R => '0',
   Q => W_reg_2_30
);
W_reg_2_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_2_31,
   R => '0',
   Q => W_reg_2_31
);
W_reg_2_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_2_3,
   R => '0',
   Q => W_reg_2_3
);
W_reg_2_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_2_4,
   R => '0',
   Q => W_reg_2_4
);
W_reg_2_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_2_5,
   R => '0',
   Q => W_reg_2_5
);
W_reg_2_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_2_6,
   R => '0',
   Q => W_reg_2_6
);
W_reg_2_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_2_7,
   R => '0',
   Q => W_reg_2_7
);
W_reg_2_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_2_8,
   R => '0',
   Q => W_reg_2_8
);
W_reg_2_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_2_9,
   R => '0',
   Q => W_reg_2_9
);
W_reg_30_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x96_out_0,
   R => '0',
   Q => W_reg_30_0
);
W_reg_30_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x96_out_10,
   R => '0',
   Q => W_reg_30_10
);
W_reg_30_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x96_out_11,
   R => '0',
   Q => W_reg_30_11
);
W_reg_30_11_i_1 : CARRY4
 port map (
   CI => W_reg_30_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_30_11_i_5_n_0,
   DI(1) => W_30_11_i_4_n_0,
   DI(2) => W_30_11_i_3_n_0,
   DI(3) => W_30_11_i_2_n_0,
   S(0) => W_30_11_i_9_n_0,
   S(1) => W_30_11_i_8_n_0,
   S(2) => W_30_11_i_7_n_0,
   S(3) => W_30_11_i_6_n_0,
   CO(0) => W_reg_30_11_i_1_n_3,
   CO(1) => W_reg_30_11_i_1_n_2,
   CO(2) => W_reg_30_11_i_1_n_1,
   CO(3) => W_reg_30_11_i_1_n_0,
   O(0) => x96_out_8,
   O(1) => x96_out_9,
   O(2) => x96_out_10,
   O(3) => x96_out_11
);
W_reg_30_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x96_out_12,
   R => '0',
   Q => W_reg_30_12
);
W_reg_30_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x96_out_13,
   R => '0',
   Q => W_reg_30_13
);
W_reg_30_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x96_out_14,
   R => '0',
   Q => W_reg_30_14
);
W_reg_30_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x96_out_15,
   R => '0',
   Q => W_reg_30_15
);
W_reg_30_15_i_1 : CARRY4
 port map (
   CI => W_reg_30_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_30_15_i_5_n_0,
   DI(1) => W_30_15_i_4_n_0,
   DI(2) => W_30_15_i_3_n_0,
   DI(3) => W_30_15_i_2_n_0,
   S(0) => W_30_15_i_9_n_0,
   S(1) => W_30_15_i_8_n_0,
   S(2) => W_30_15_i_7_n_0,
   S(3) => W_30_15_i_6_n_0,
   CO(0) => W_reg_30_15_i_1_n_3,
   CO(1) => W_reg_30_15_i_1_n_2,
   CO(2) => W_reg_30_15_i_1_n_1,
   CO(3) => W_reg_30_15_i_1_n_0,
   O(0) => x96_out_12,
   O(1) => x96_out_13,
   O(2) => x96_out_14,
   O(3) => x96_out_15
);
W_reg_30_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x96_out_16,
   R => '0',
   Q => W_reg_30_16
);
W_reg_30_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x96_out_17,
   R => '0',
   Q => W_reg_30_17
);
W_reg_30_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x96_out_18,
   R => '0',
   Q => W_reg_30_18
);
W_reg_30_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x96_out_19,
   R => '0',
   Q => W_reg_30_19
);
W_reg_30_19_i_1 : CARRY4
 port map (
   CI => W_reg_30_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_30_19_i_5_n_0,
   DI(1) => W_30_19_i_4_n_0,
   DI(2) => W_30_19_i_3_n_0,
   DI(3) => W_30_19_i_2_n_0,
   S(0) => W_30_19_i_9_n_0,
   S(1) => W_30_19_i_8_n_0,
   S(2) => W_30_19_i_7_n_0,
   S(3) => W_30_19_i_6_n_0,
   CO(0) => W_reg_30_19_i_1_n_3,
   CO(1) => W_reg_30_19_i_1_n_2,
   CO(2) => W_reg_30_19_i_1_n_1,
   CO(3) => W_reg_30_19_i_1_n_0,
   O(0) => x96_out_16,
   O(1) => x96_out_17,
   O(2) => x96_out_18,
   O(3) => x96_out_19
);
W_reg_30_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x96_out_1,
   R => '0',
   Q => W_reg_30_1
);
W_reg_30_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x96_out_20,
   R => '0',
   Q => W_reg_30_20
);
W_reg_30_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x96_out_21,
   R => '0',
   Q => W_reg_30_21
);
W_reg_30_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x96_out_22,
   R => '0',
   Q => W_reg_30_22
);
W_reg_30_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x96_out_23,
   R => '0',
   Q => W_reg_30_23
);
W_reg_30_23_i_1 : CARRY4
 port map (
   CI => W_reg_30_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_30_23_i_5_n_0,
   DI(1) => W_30_23_i_4_n_0,
   DI(2) => W_30_23_i_3_n_0,
   DI(3) => W_30_23_i_2_n_0,
   S(0) => W_30_23_i_9_n_0,
   S(1) => W_30_23_i_8_n_0,
   S(2) => W_30_23_i_7_n_0,
   S(3) => W_30_23_i_6_n_0,
   CO(0) => W_reg_30_23_i_1_n_3,
   CO(1) => W_reg_30_23_i_1_n_2,
   CO(2) => W_reg_30_23_i_1_n_1,
   CO(3) => W_reg_30_23_i_1_n_0,
   O(0) => x96_out_20,
   O(1) => x96_out_21,
   O(2) => x96_out_22,
   O(3) => x96_out_23
);
W_reg_30_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x96_out_24,
   R => '0',
   Q => W_reg_30_24
);
W_reg_30_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x96_out_25,
   R => '0',
   Q => W_reg_30_25
);
W_reg_30_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x96_out_26,
   R => '0',
   Q => W_reg_30_26
);
W_reg_30_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x96_out_27,
   R => '0',
   Q => W_reg_30_27
);
W_reg_30_27_i_1 : CARRY4
 port map (
   CI => W_reg_30_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_30_27_i_5_n_0,
   DI(1) => W_30_27_i_4_n_0,
   DI(2) => W_30_27_i_3_n_0,
   DI(3) => W_30_27_i_2_n_0,
   S(0) => W_30_27_i_9_n_0,
   S(1) => W_30_27_i_8_n_0,
   S(2) => W_30_27_i_7_n_0,
   S(3) => W_30_27_i_6_n_0,
   CO(0) => W_reg_30_27_i_1_n_3,
   CO(1) => W_reg_30_27_i_1_n_2,
   CO(2) => W_reg_30_27_i_1_n_1,
   CO(3) => W_reg_30_27_i_1_n_0,
   O(0) => x96_out_24,
   O(1) => x96_out_25,
   O(2) => x96_out_26,
   O(3) => x96_out_27
);
W_reg_30_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x96_out_28,
   R => '0',
   Q => W_reg_30_28
);
W_reg_30_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x96_out_29,
   R => '0',
   Q => W_reg_30_29
);
W_reg_30_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x96_out_2,
   R => '0',
   Q => W_reg_30_2
);
W_reg_30_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x96_out_30,
   R => '0',
   Q => W_reg_30_30
);
W_reg_30_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x96_out_31,
   R => '0',
   Q => W_reg_30_31
);
W_reg_30_31_i_1 : CARRY4
 port map (
   CI => W_reg_30_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_30_31_i_4_n_0,
   DI(1) => W_30_31_i_3_n_0,
   DI(2) => W_30_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_30_31_i_8_n_0,
   S(1) => W_30_31_i_7_n_0,
   S(2) => W_30_31_i_6_n_0,
   S(3) => W_30_31_i_5_n_0,
   CO(0) => W_reg_30_31_i_1_n_3,
   CO(1) => W_reg_30_31_i_1_n_2,
   CO(2) => W_reg_30_31_i_1_n_1,
   CO(3) => NLW_W_reg_30_31_i_1_CO_UNCONNECTED_3,
   O(0) => x96_out_28,
   O(1) => x96_out_29,
   O(2) => x96_out_30,
   O(3) => x96_out_31
);
W_reg_30_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x96_out_3,
   R => '0',
   Q => W_reg_30_3
);
W_reg_30_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_30_3_i_5_n_0,
   DI(1) => W_30_3_i_4_n_0,
   DI(2) => W_30_3_i_3_n_0,
   DI(3) => W_30_3_i_2_n_0,
   S(0) => W_30_3_i_9_n_0,
   S(1) => W_30_3_i_8_n_0,
   S(2) => W_30_3_i_7_n_0,
   S(3) => W_30_3_i_6_n_0,
   CO(0) => W_reg_30_3_i_1_n_3,
   CO(1) => W_reg_30_3_i_1_n_2,
   CO(2) => W_reg_30_3_i_1_n_1,
   CO(3) => W_reg_30_3_i_1_n_0,
   O(0) => x96_out_0,
   O(1) => x96_out_1,
   O(2) => x96_out_2,
   O(3) => x96_out_3
);
W_reg_30_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x96_out_4,
   R => '0',
   Q => W_reg_30_4
);
W_reg_30_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x96_out_5,
   R => '0',
   Q => W_reg_30_5
);
W_reg_30_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x96_out_6,
   R => '0',
   Q => W_reg_30_6
);
W_reg_30_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x96_out_7,
   R => '0',
   Q => W_reg_30_7
);
W_reg_30_7_i_1 : CARRY4
 port map (
   CI => W_reg_30_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_30_7_i_5_n_0,
   DI(1) => W_30_7_i_4_n_0,
   DI(2) => W_30_7_i_3_n_0,
   DI(3) => W_30_7_i_2_n_0,
   S(0) => W_30_7_i_9_n_0,
   S(1) => W_30_7_i_8_n_0,
   S(2) => W_30_7_i_7_n_0,
   S(3) => W_30_7_i_6_n_0,
   CO(0) => W_reg_30_7_i_1_n_3,
   CO(1) => W_reg_30_7_i_1_n_2,
   CO(2) => W_reg_30_7_i_1_n_1,
   CO(3) => W_reg_30_7_i_1_n_0,
   O(0) => x96_out_4,
   O(1) => x96_out_5,
   O(2) => x96_out_6,
   O(3) => x96_out_7
);
W_reg_30_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x96_out_8,
   R => '0',
   Q => W_reg_30_8
);
W_reg_30_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x96_out_9,
   R => '0',
   Q => W_reg_30_9
);
W_reg_31_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x94_out_0,
   R => '0',
   Q => W_reg_31_0
);
W_reg_31_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x94_out_10,
   R => '0',
   Q => W_reg_31_10
);
W_reg_31_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x94_out_11,
   R => '0',
   Q => W_reg_31_11
);
W_reg_31_11_i_1 : CARRY4
 port map (
   CI => W_reg_31_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_31_11_i_5_n_0,
   DI(1) => W_31_11_i_4_n_0,
   DI(2) => W_31_11_i_3_n_0,
   DI(3) => W_31_11_i_2_n_0,
   S(0) => W_31_11_i_9_n_0,
   S(1) => W_31_11_i_8_n_0,
   S(2) => W_31_11_i_7_n_0,
   S(3) => W_31_11_i_6_n_0,
   CO(0) => W_reg_31_11_i_1_n_3,
   CO(1) => W_reg_31_11_i_1_n_2,
   CO(2) => W_reg_31_11_i_1_n_1,
   CO(3) => W_reg_31_11_i_1_n_0,
   O(0) => x94_out_8,
   O(1) => x94_out_9,
   O(2) => x94_out_10,
   O(3) => x94_out_11
);
W_reg_31_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x94_out_12,
   R => '0',
   Q => W_reg_31_12
);
W_reg_31_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x94_out_13,
   R => '0',
   Q => W_reg_31_13
);
W_reg_31_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x94_out_14,
   R => '0',
   Q => W_reg_31_14
);
W_reg_31_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x94_out_15,
   R => '0',
   Q => W_reg_31_15
);
W_reg_31_15_i_1 : CARRY4
 port map (
   CI => W_reg_31_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_31_15_i_5_n_0,
   DI(1) => W_31_15_i_4_n_0,
   DI(2) => W_31_15_i_3_n_0,
   DI(3) => W_31_15_i_2_n_0,
   S(0) => W_31_15_i_9_n_0,
   S(1) => W_31_15_i_8_n_0,
   S(2) => W_31_15_i_7_n_0,
   S(3) => W_31_15_i_6_n_0,
   CO(0) => W_reg_31_15_i_1_n_3,
   CO(1) => W_reg_31_15_i_1_n_2,
   CO(2) => W_reg_31_15_i_1_n_1,
   CO(3) => W_reg_31_15_i_1_n_0,
   O(0) => x94_out_12,
   O(1) => x94_out_13,
   O(2) => x94_out_14,
   O(3) => x94_out_15
);
W_reg_31_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x94_out_16,
   R => '0',
   Q => W_reg_31_16
);
W_reg_31_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x94_out_17,
   R => '0',
   Q => W_reg_31_17
);
W_reg_31_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x94_out_18,
   R => '0',
   Q => W_reg_31_18
);
W_reg_31_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x94_out_19,
   R => '0',
   Q => W_reg_31_19
);
W_reg_31_19_i_1 : CARRY4
 port map (
   CI => W_reg_31_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_31_19_i_5_n_0,
   DI(1) => W_31_19_i_4_n_0,
   DI(2) => W_31_19_i_3_n_0,
   DI(3) => W_31_19_i_2_n_0,
   S(0) => W_31_19_i_9_n_0,
   S(1) => W_31_19_i_8_n_0,
   S(2) => W_31_19_i_7_n_0,
   S(3) => W_31_19_i_6_n_0,
   CO(0) => W_reg_31_19_i_1_n_3,
   CO(1) => W_reg_31_19_i_1_n_2,
   CO(2) => W_reg_31_19_i_1_n_1,
   CO(3) => W_reg_31_19_i_1_n_0,
   O(0) => x94_out_16,
   O(1) => x94_out_17,
   O(2) => x94_out_18,
   O(3) => x94_out_19
);
W_reg_31_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x94_out_1,
   R => '0',
   Q => W_reg_31_1
);
W_reg_31_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x94_out_20,
   R => '0',
   Q => W_reg_31_20
);
W_reg_31_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x94_out_21,
   R => '0',
   Q => W_reg_31_21
);
W_reg_31_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x94_out_22,
   R => '0',
   Q => W_reg_31_22
);
W_reg_31_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x94_out_23,
   R => '0',
   Q => W_reg_31_23
);
W_reg_31_23_i_1 : CARRY4
 port map (
   CI => W_reg_31_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_31_23_i_5_n_0,
   DI(1) => W_31_23_i_4_n_0,
   DI(2) => W_31_23_i_3_n_0,
   DI(3) => W_31_23_i_2_n_0,
   S(0) => W_31_23_i_9_n_0,
   S(1) => W_31_23_i_8_n_0,
   S(2) => W_31_23_i_7_n_0,
   S(3) => W_31_23_i_6_n_0,
   CO(0) => W_reg_31_23_i_1_n_3,
   CO(1) => W_reg_31_23_i_1_n_2,
   CO(2) => W_reg_31_23_i_1_n_1,
   CO(3) => W_reg_31_23_i_1_n_0,
   O(0) => x94_out_20,
   O(1) => x94_out_21,
   O(2) => x94_out_22,
   O(3) => x94_out_23
);
W_reg_31_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x94_out_24,
   R => '0',
   Q => W_reg_31_24
);
W_reg_31_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x94_out_25,
   R => '0',
   Q => W_reg_31_25
);
W_reg_31_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x94_out_26,
   R => '0',
   Q => W_reg_31_26
);
W_reg_31_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x94_out_27,
   R => '0',
   Q => W_reg_31_27
);
W_reg_31_27_i_1 : CARRY4
 port map (
   CI => W_reg_31_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_31_27_i_5_n_0,
   DI(1) => W_31_27_i_4_n_0,
   DI(2) => W_31_27_i_3_n_0,
   DI(3) => W_31_27_i_2_n_0,
   S(0) => W_31_27_i_9_n_0,
   S(1) => W_31_27_i_8_n_0,
   S(2) => W_31_27_i_7_n_0,
   S(3) => W_31_27_i_6_n_0,
   CO(0) => W_reg_31_27_i_1_n_3,
   CO(1) => W_reg_31_27_i_1_n_2,
   CO(2) => W_reg_31_27_i_1_n_1,
   CO(3) => W_reg_31_27_i_1_n_0,
   O(0) => x94_out_24,
   O(1) => x94_out_25,
   O(2) => x94_out_26,
   O(3) => x94_out_27
);
W_reg_31_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x94_out_28,
   R => '0',
   Q => W_reg_31_28
);
W_reg_31_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x94_out_29,
   R => '0',
   Q => W_reg_31_29
);
W_reg_31_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x94_out_2,
   R => '0',
   Q => W_reg_31_2
);
W_reg_31_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x94_out_30,
   R => '0',
   Q => W_reg_31_30
);
W_reg_31_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x94_out_31,
   R => '0',
   Q => W_reg_31_31
);
W_reg_31_31_i_1 : CARRY4
 port map (
   CI => W_reg_31_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_31_31_i_4_n_0,
   DI(1) => W_31_31_i_3_n_0,
   DI(2) => W_31_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_31_31_i_8_n_0,
   S(1) => W_31_31_i_7_n_0,
   S(2) => W_31_31_i_6_n_0,
   S(3) => W_31_31_i_5_n_0,
   CO(0) => W_reg_31_31_i_1_n_3,
   CO(1) => W_reg_31_31_i_1_n_2,
   CO(2) => W_reg_31_31_i_1_n_1,
   CO(3) => NLW_W_reg_31_31_i_1_CO_UNCONNECTED_3,
   O(0) => x94_out_28,
   O(1) => x94_out_29,
   O(2) => x94_out_30,
   O(3) => x94_out_31
);
W_reg_31_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x94_out_3,
   R => '0',
   Q => W_reg_31_3
);
W_reg_31_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_31_3_i_5_n_0,
   DI(1) => W_31_3_i_4_n_0,
   DI(2) => W_31_3_i_3_n_0,
   DI(3) => W_31_3_i_2_n_0,
   S(0) => W_31_3_i_9_n_0,
   S(1) => W_31_3_i_8_n_0,
   S(2) => W_31_3_i_7_n_0,
   S(3) => W_31_3_i_6_n_0,
   CO(0) => W_reg_31_3_i_1_n_3,
   CO(1) => W_reg_31_3_i_1_n_2,
   CO(2) => W_reg_31_3_i_1_n_1,
   CO(3) => W_reg_31_3_i_1_n_0,
   O(0) => x94_out_0,
   O(1) => x94_out_1,
   O(2) => x94_out_2,
   O(3) => x94_out_3
);
W_reg_31_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x94_out_4,
   R => '0',
   Q => W_reg_31_4
);
W_reg_31_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x94_out_5,
   R => '0',
   Q => W_reg_31_5
);
W_reg_31_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x94_out_6,
   R => '0',
   Q => W_reg_31_6
);
W_reg_31_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x94_out_7,
   R => '0',
   Q => W_reg_31_7
);
W_reg_31_7_i_1 : CARRY4
 port map (
   CI => W_reg_31_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_31_7_i_5_n_0,
   DI(1) => W_31_7_i_4_n_0,
   DI(2) => W_31_7_i_3_n_0,
   DI(3) => W_31_7_i_2_n_0,
   S(0) => W_31_7_i_9_n_0,
   S(1) => W_31_7_i_8_n_0,
   S(2) => W_31_7_i_7_n_0,
   S(3) => W_31_7_i_6_n_0,
   CO(0) => W_reg_31_7_i_1_n_3,
   CO(1) => W_reg_31_7_i_1_n_2,
   CO(2) => W_reg_31_7_i_1_n_1,
   CO(3) => W_reg_31_7_i_1_n_0,
   O(0) => x94_out_4,
   O(1) => x94_out_5,
   O(2) => x94_out_6,
   O(3) => x94_out_7
);
W_reg_31_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x94_out_8,
   R => '0',
   Q => W_reg_31_8
);
W_reg_31_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_16_0,
   D => x94_out_9,
   R => '0',
   Q => W_reg_31_9
);
W_reg_32_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x92_out_0,
   R => '0',
   Q => W_reg_32_0
);
W_reg_32_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x92_out_10,
   R => '0',
   Q => W_reg_32_10
);
W_reg_32_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x92_out_11,
   R => '0',
   Q => W_reg_32_11
);
W_reg_32_11_i_1 : CARRY4
 port map (
   CI => W_reg_32_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_32_11_i_5_n_0,
   DI(1) => W_32_11_i_4_n_0,
   DI(2) => W_32_11_i_3_n_0,
   DI(3) => W_32_11_i_2_n_0,
   S(0) => W_32_11_i_9_n_0,
   S(1) => W_32_11_i_8_n_0,
   S(2) => W_32_11_i_7_n_0,
   S(3) => W_32_11_i_6_n_0,
   CO(0) => W_reg_32_11_i_1_n_3,
   CO(1) => W_reg_32_11_i_1_n_2,
   CO(2) => W_reg_32_11_i_1_n_1,
   CO(3) => W_reg_32_11_i_1_n_0,
   O(0) => x92_out_8,
   O(1) => x92_out_9,
   O(2) => x92_out_10,
   O(3) => x92_out_11
);
W_reg_32_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x92_out_12,
   R => '0',
   Q => W_reg_32_12
);
W_reg_32_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x92_out_13,
   R => '0',
   Q => W_reg_32_13
);
W_reg_32_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x92_out_14,
   R => '0',
   Q => W_reg_32_14
);
W_reg_32_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x92_out_15,
   R => '0',
   Q => W_reg_32_15
);
W_reg_32_15_i_1 : CARRY4
 port map (
   CI => W_reg_32_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_32_15_i_5_n_0,
   DI(1) => W_32_15_i_4_n_0,
   DI(2) => W_32_15_i_3_n_0,
   DI(3) => W_32_15_i_2_n_0,
   S(0) => W_32_15_i_9_n_0,
   S(1) => W_32_15_i_8_n_0,
   S(2) => W_32_15_i_7_n_0,
   S(3) => W_32_15_i_6_n_0,
   CO(0) => W_reg_32_15_i_1_n_3,
   CO(1) => W_reg_32_15_i_1_n_2,
   CO(2) => W_reg_32_15_i_1_n_1,
   CO(3) => W_reg_32_15_i_1_n_0,
   O(0) => x92_out_12,
   O(1) => x92_out_13,
   O(2) => x92_out_14,
   O(3) => x92_out_15
);
W_reg_32_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x92_out_16,
   R => '0',
   Q => W_reg_32_16
);
W_reg_32_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x92_out_17,
   R => '0',
   Q => W_reg_32_17
);
W_reg_32_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x92_out_18,
   R => '0',
   Q => W_reg_32_18
);
W_reg_32_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x92_out_19,
   R => '0',
   Q => W_reg_32_19
);
W_reg_32_19_i_1 : CARRY4
 port map (
   CI => W_reg_32_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_32_19_i_5_n_0,
   DI(1) => W_32_19_i_4_n_0,
   DI(2) => W_32_19_i_3_n_0,
   DI(3) => W_32_19_i_2_n_0,
   S(0) => W_32_19_i_9_n_0,
   S(1) => W_32_19_i_8_n_0,
   S(2) => W_32_19_i_7_n_0,
   S(3) => W_32_19_i_6_n_0,
   CO(0) => W_reg_32_19_i_1_n_3,
   CO(1) => W_reg_32_19_i_1_n_2,
   CO(2) => W_reg_32_19_i_1_n_1,
   CO(3) => W_reg_32_19_i_1_n_0,
   O(0) => x92_out_16,
   O(1) => x92_out_17,
   O(2) => x92_out_18,
   O(3) => x92_out_19
);
W_reg_32_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x92_out_1,
   R => '0',
   Q => W_reg_32_1
);
W_reg_32_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x92_out_20,
   R => '0',
   Q => W_reg_32_20
);
W_reg_32_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x92_out_21,
   R => '0',
   Q => W_reg_32_21
);
W_reg_32_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x92_out_22,
   R => '0',
   Q => W_reg_32_22
);
W_reg_32_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x92_out_23,
   R => '0',
   Q => W_reg_32_23
);
W_reg_32_23_i_1 : CARRY4
 port map (
   CI => W_reg_32_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_32_23_i_5_n_0,
   DI(1) => W_32_23_i_4_n_0,
   DI(2) => W_32_23_i_3_n_0,
   DI(3) => W_32_23_i_2_n_0,
   S(0) => W_32_23_i_9_n_0,
   S(1) => W_32_23_i_8_n_0,
   S(2) => W_32_23_i_7_n_0,
   S(3) => W_32_23_i_6_n_0,
   CO(0) => W_reg_32_23_i_1_n_3,
   CO(1) => W_reg_32_23_i_1_n_2,
   CO(2) => W_reg_32_23_i_1_n_1,
   CO(3) => W_reg_32_23_i_1_n_0,
   O(0) => x92_out_20,
   O(1) => x92_out_21,
   O(2) => x92_out_22,
   O(3) => x92_out_23
);
W_reg_32_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x92_out_24,
   R => '0',
   Q => W_reg_32_24
);
W_reg_32_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x92_out_25,
   R => '0',
   Q => W_reg_32_25
);
W_reg_32_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x92_out_26,
   R => '0',
   Q => W_reg_32_26
);
W_reg_32_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x92_out_27,
   R => '0',
   Q => W_reg_32_27
);
W_reg_32_27_i_1 : CARRY4
 port map (
   CI => W_reg_32_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_32_27_i_5_n_0,
   DI(1) => W_32_27_i_4_n_0,
   DI(2) => W_32_27_i_3_n_0,
   DI(3) => W_32_27_i_2_n_0,
   S(0) => W_32_27_i_9_n_0,
   S(1) => W_32_27_i_8_n_0,
   S(2) => W_32_27_i_7_n_0,
   S(3) => W_32_27_i_6_n_0,
   CO(0) => W_reg_32_27_i_1_n_3,
   CO(1) => W_reg_32_27_i_1_n_2,
   CO(2) => W_reg_32_27_i_1_n_1,
   CO(3) => W_reg_32_27_i_1_n_0,
   O(0) => x92_out_24,
   O(1) => x92_out_25,
   O(2) => x92_out_26,
   O(3) => x92_out_27
);
W_reg_32_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x92_out_28,
   R => '0',
   Q => W_reg_32_28
);
W_reg_32_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x92_out_29,
   R => '0',
   Q => W_reg_32_29
);
W_reg_32_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x92_out_2,
   R => '0',
   Q => W_reg_32_2
);
W_reg_32_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x92_out_30,
   R => '0',
   Q => W_reg_32_30
);
W_reg_32_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x92_out_31,
   R => '0',
   Q => W_reg_32_31
);
W_reg_32_31_i_2 : CARRY4
 port map (
   CI => W_reg_32_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_32_31_i_5_n_0,
   DI(1) => W_32_31_i_4_n_0,
   DI(2) => W_32_31_i_3_n_0,
   DI(3) => '0',
   S(0) => W_32_31_i_9_n_0,
   S(1) => W_32_31_i_8_n_0,
   S(2) => W_32_31_i_7_n_0,
   S(3) => W_32_31_i_6_n_0,
   CO(0) => W_reg_32_31_i_2_n_3,
   CO(1) => W_reg_32_31_i_2_n_2,
   CO(2) => W_reg_32_31_i_2_n_1,
   CO(3) => NLW_W_reg_32_31_i_2_CO_UNCONNECTED_3,
   O(0) => x92_out_28,
   O(1) => x92_out_29,
   O(2) => x92_out_30,
   O(3) => x92_out_31
);
W_reg_32_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x92_out_3,
   R => '0',
   Q => W_reg_32_3
);
W_reg_32_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_32_3_i_5_n_0,
   DI(1) => W_32_3_i_4_n_0,
   DI(2) => W_32_3_i_3_n_0,
   DI(3) => W_32_3_i_2_n_0,
   S(0) => W_32_3_i_9_n_0,
   S(1) => W_32_3_i_8_n_0,
   S(2) => W_32_3_i_7_n_0,
   S(3) => W_32_3_i_6_n_0,
   CO(0) => W_reg_32_3_i_1_n_3,
   CO(1) => W_reg_32_3_i_1_n_2,
   CO(2) => W_reg_32_3_i_1_n_1,
   CO(3) => W_reg_32_3_i_1_n_0,
   O(0) => x92_out_0,
   O(1) => x92_out_1,
   O(2) => x92_out_2,
   O(3) => x92_out_3
);
W_reg_32_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x92_out_4,
   R => '0',
   Q => W_reg_32_4
);
W_reg_32_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x92_out_5,
   R => '0',
   Q => W_reg_32_5
);
W_reg_32_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x92_out_6,
   R => '0',
   Q => W_reg_32_6
);
W_reg_32_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x92_out_7,
   R => '0',
   Q => W_reg_32_7
);
W_reg_32_7_i_1 : CARRY4
 port map (
   CI => W_reg_32_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_32_7_i_5_n_0,
   DI(1) => W_32_7_i_4_n_0,
   DI(2) => W_32_7_i_3_n_0,
   DI(3) => W_32_7_i_2_n_0,
   S(0) => W_32_7_i_9_n_0,
   S(1) => W_32_7_i_8_n_0,
   S(2) => W_32_7_i_7_n_0,
   S(3) => W_32_7_i_6_n_0,
   CO(0) => W_reg_32_7_i_1_n_3,
   CO(1) => W_reg_32_7_i_1_n_2,
   CO(2) => W_reg_32_7_i_1_n_1,
   CO(3) => W_reg_32_7_i_1_n_0,
   O(0) => x92_out_4,
   O(1) => x92_out_5,
   O(2) => x92_out_6,
   O(3) => x92_out_7
);
W_reg_32_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x92_out_8,
   R => '0',
   Q => W_reg_32_8
);
W_reg_32_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x92_out_9,
   R => '0',
   Q => W_reg_32_9
);
W_reg_33_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x89_out_0,
   R => '0',
   Q => W_reg_33_0
);
W_reg_33_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x89_out_10,
   R => '0',
   Q => W_reg_33_10
);
W_reg_33_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x89_out_11,
   R => '0',
   Q => W_reg_33_11
);
W_reg_33_11_i_1 : CARRY4
 port map (
   CI => W_reg_33_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_33_11_i_5_n_0,
   DI(1) => W_33_11_i_4_n_0,
   DI(2) => W_33_11_i_3_n_0,
   DI(3) => W_33_11_i_2_n_0,
   S(0) => W_33_11_i_9_n_0,
   S(1) => W_33_11_i_8_n_0,
   S(2) => W_33_11_i_7_n_0,
   S(3) => W_33_11_i_6_n_0,
   CO(0) => W_reg_33_11_i_1_n_3,
   CO(1) => W_reg_33_11_i_1_n_2,
   CO(2) => W_reg_33_11_i_1_n_1,
   CO(3) => W_reg_33_11_i_1_n_0,
   O(0) => x89_out_8,
   O(1) => x89_out_9,
   O(2) => x89_out_10,
   O(3) => x89_out_11
);
W_reg_33_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x89_out_12,
   R => '0',
   Q => W_reg_33_12
);
W_reg_33_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x89_out_13,
   R => '0',
   Q => W_reg_33_13
);
W_reg_33_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x89_out_14,
   R => '0',
   Q => W_reg_33_14
);
W_reg_33_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x89_out_15,
   R => '0',
   Q => W_reg_33_15
);
W_reg_33_15_i_1 : CARRY4
 port map (
   CI => W_reg_33_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_33_15_i_5_n_0,
   DI(1) => W_33_15_i_4_n_0,
   DI(2) => W_33_15_i_3_n_0,
   DI(3) => W_33_15_i_2_n_0,
   S(0) => W_33_15_i_9_n_0,
   S(1) => W_33_15_i_8_n_0,
   S(2) => W_33_15_i_7_n_0,
   S(3) => W_33_15_i_6_n_0,
   CO(0) => W_reg_33_15_i_1_n_3,
   CO(1) => W_reg_33_15_i_1_n_2,
   CO(2) => W_reg_33_15_i_1_n_1,
   CO(3) => W_reg_33_15_i_1_n_0,
   O(0) => x89_out_12,
   O(1) => x89_out_13,
   O(2) => x89_out_14,
   O(3) => x89_out_15
);
W_reg_33_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x89_out_16,
   R => '0',
   Q => W_reg_33_16
);
W_reg_33_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x89_out_17,
   R => '0',
   Q => W_reg_33_17
);
W_reg_33_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x89_out_18,
   R => '0',
   Q => W_reg_33_18
);
W_reg_33_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x89_out_19,
   R => '0',
   Q => W_reg_33_19
);
W_reg_33_19_i_1 : CARRY4
 port map (
   CI => W_reg_33_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_33_19_i_5_n_0,
   DI(1) => W_33_19_i_4_n_0,
   DI(2) => W_33_19_i_3_n_0,
   DI(3) => W_33_19_i_2_n_0,
   S(0) => W_33_19_i_9_n_0,
   S(1) => W_33_19_i_8_n_0,
   S(2) => W_33_19_i_7_n_0,
   S(3) => W_33_19_i_6_n_0,
   CO(0) => W_reg_33_19_i_1_n_3,
   CO(1) => W_reg_33_19_i_1_n_2,
   CO(2) => W_reg_33_19_i_1_n_1,
   CO(3) => W_reg_33_19_i_1_n_0,
   O(0) => x89_out_16,
   O(1) => x89_out_17,
   O(2) => x89_out_18,
   O(3) => x89_out_19
);
W_reg_33_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x89_out_1,
   R => '0',
   Q => W_reg_33_1
);
W_reg_33_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x89_out_20,
   R => '0',
   Q => W_reg_33_20
);
W_reg_33_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x89_out_21,
   R => '0',
   Q => W_reg_33_21
);
W_reg_33_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x89_out_22,
   R => '0',
   Q => W_reg_33_22
);
W_reg_33_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x89_out_23,
   R => '0',
   Q => W_reg_33_23
);
W_reg_33_23_i_1 : CARRY4
 port map (
   CI => W_reg_33_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_33_23_i_5_n_0,
   DI(1) => W_33_23_i_4_n_0,
   DI(2) => W_33_23_i_3_n_0,
   DI(3) => W_33_23_i_2_n_0,
   S(0) => W_33_23_i_9_n_0,
   S(1) => W_33_23_i_8_n_0,
   S(2) => W_33_23_i_7_n_0,
   S(3) => W_33_23_i_6_n_0,
   CO(0) => W_reg_33_23_i_1_n_3,
   CO(1) => W_reg_33_23_i_1_n_2,
   CO(2) => W_reg_33_23_i_1_n_1,
   CO(3) => W_reg_33_23_i_1_n_0,
   O(0) => x89_out_20,
   O(1) => x89_out_21,
   O(2) => x89_out_22,
   O(3) => x89_out_23
);
W_reg_33_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x89_out_24,
   R => '0',
   Q => W_reg_33_24
);
W_reg_33_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x89_out_25,
   R => '0',
   Q => W_reg_33_25
);
W_reg_33_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x89_out_26,
   R => '0',
   Q => W_reg_33_26
);
W_reg_33_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x89_out_27,
   R => '0',
   Q => W_reg_33_27
);
W_reg_33_27_i_1 : CARRY4
 port map (
   CI => W_reg_33_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_33_27_i_5_n_0,
   DI(1) => W_33_27_i_4_n_0,
   DI(2) => W_33_27_i_3_n_0,
   DI(3) => W_33_27_i_2_n_0,
   S(0) => W_33_27_i_9_n_0,
   S(1) => W_33_27_i_8_n_0,
   S(2) => W_33_27_i_7_n_0,
   S(3) => W_33_27_i_6_n_0,
   CO(0) => W_reg_33_27_i_1_n_3,
   CO(1) => W_reg_33_27_i_1_n_2,
   CO(2) => W_reg_33_27_i_1_n_1,
   CO(3) => W_reg_33_27_i_1_n_0,
   O(0) => x89_out_24,
   O(1) => x89_out_25,
   O(2) => x89_out_26,
   O(3) => x89_out_27
);
W_reg_33_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x89_out_28,
   R => '0',
   Q => W_reg_33_28
);
W_reg_33_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x89_out_29,
   R => '0',
   Q => W_reg_33_29
);
W_reg_33_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x89_out_2,
   R => '0',
   Q => W_reg_33_2
);
W_reg_33_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x89_out_30,
   R => '0',
   Q => W_reg_33_30
);
W_reg_33_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x89_out_31,
   R => '0',
   Q => W_reg_33_31
);
W_reg_33_31_i_1 : CARRY4
 port map (
   CI => W_reg_33_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_33_31_i_4_n_0,
   DI(1) => W_33_31_i_3_n_0,
   DI(2) => W_33_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_33_31_i_8_n_0,
   S(1) => W_33_31_i_7_n_0,
   S(2) => W_33_31_i_6_n_0,
   S(3) => W_33_31_i_5_n_0,
   CO(0) => W_reg_33_31_i_1_n_3,
   CO(1) => W_reg_33_31_i_1_n_2,
   CO(2) => W_reg_33_31_i_1_n_1,
   CO(3) => NLW_W_reg_33_31_i_1_CO_UNCONNECTED_3,
   O(0) => x89_out_28,
   O(1) => x89_out_29,
   O(2) => x89_out_30,
   O(3) => x89_out_31
);
W_reg_33_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x89_out_3,
   R => '0',
   Q => W_reg_33_3
);
W_reg_33_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_33_3_i_5_n_0,
   DI(1) => W_33_3_i_4_n_0,
   DI(2) => W_33_3_i_3_n_0,
   DI(3) => W_33_3_i_2_n_0,
   S(0) => W_33_3_i_9_n_0,
   S(1) => W_33_3_i_8_n_0,
   S(2) => W_33_3_i_7_n_0,
   S(3) => W_33_3_i_6_n_0,
   CO(0) => W_reg_33_3_i_1_n_3,
   CO(1) => W_reg_33_3_i_1_n_2,
   CO(2) => W_reg_33_3_i_1_n_1,
   CO(3) => W_reg_33_3_i_1_n_0,
   O(0) => x89_out_0,
   O(1) => x89_out_1,
   O(2) => x89_out_2,
   O(3) => x89_out_3
);
W_reg_33_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x89_out_4,
   R => '0',
   Q => W_reg_33_4
);
W_reg_33_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x89_out_5,
   R => '0',
   Q => W_reg_33_5
);
W_reg_33_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x89_out_6,
   R => '0',
   Q => W_reg_33_6
);
W_reg_33_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x89_out_7,
   R => '0',
   Q => W_reg_33_7
);
W_reg_33_7_i_1 : CARRY4
 port map (
   CI => W_reg_33_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_33_7_i_5_n_0,
   DI(1) => W_33_7_i_4_n_0,
   DI(2) => W_33_7_i_3_n_0,
   DI(3) => W_33_7_i_2_n_0,
   S(0) => W_33_7_i_9_n_0,
   S(1) => W_33_7_i_8_n_0,
   S(2) => W_33_7_i_7_n_0,
   S(3) => W_33_7_i_6_n_0,
   CO(0) => W_reg_33_7_i_1_n_3,
   CO(1) => W_reg_33_7_i_1_n_2,
   CO(2) => W_reg_33_7_i_1_n_1,
   CO(3) => W_reg_33_7_i_1_n_0,
   O(0) => x89_out_4,
   O(1) => x89_out_5,
   O(2) => x89_out_6,
   O(3) => x89_out_7
);
W_reg_33_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x89_out_8,
   R => '0',
   Q => W_reg_33_8
);
W_reg_33_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x89_out_9,
   R => '0',
   Q => W_reg_33_9
);
W_reg_34_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x86_out_0,
   R => '0',
   Q => W_reg_34_0
);
W_reg_34_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x86_out_10,
   R => '0',
   Q => W_reg_34_10
);
W_reg_34_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x86_out_11,
   R => '0',
   Q => W_reg_34_11
);
W_reg_34_11_i_1 : CARRY4
 port map (
   CI => W_reg_34_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_34_11_i_5_n_0,
   DI(1) => W_34_11_i_4_n_0,
   DI(2) => W_34_11_i_3_n_0,
   DI(3) => W_34_11_i_2_n_0,
   S(0) => W_34_11_i_9_n_0,
   S(1) => W_34_11_i_8_n_0,
   S(2) => W_34_11_i_7_n_0,
   S(3) => W_34_11_i_6_n_0,
   CO(0) => W_reg_34_11_i_1_n_3,
   CO(1) => W_reg_34_11_i_1_n_2,
   CO(2) => W_reg_34_11_i_1_n_1,
   CO(3) => W_reg_34_11_i_1_n_0,
   O(0) => x86_out_8,
   O(1) => x86_out_9,
   O(2) => x86_out_10,
   O(3) => x86_out_11
);
W_reg_34_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x86_out_12,
   R => '0',
   Q => W_reg_34_12
);
W_reg_34_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x86_out_13,
   R => '0',
   Q => W_reg_34_13
);
W_reg_34_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x86_out_14,
   R => '0',
   Q => W_reg_34_14
);
W_reg_34_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x86_out_15,
   R => '0',
   Q => W_reg_34_15
);
W_reg_34_15_i_1 : CARRY4
 port map (
   CI => W_reg_34_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_34_15_i_5_n_0,
   DI(1) => W_34_15_i_4_n_0,
   DI(2) => W_34_15_i_3_n_0,
   DI(3) => W_34_15_i_2_n_0,
   S(0) => W_34_15_i_9_n_0,
   S(1) => W_34_15_i_8_n_0,
   S(2) => W_34_15_i_7_n_0,
   S(3) => W_34_15_i_6_n_0,
   CO(0) => W_reg_34_15_i_1_n_3,
   CO(1) => W_reg_34_15_i_1_n_2,
   CO(2) => W_reg_34_15_i_1_n_1,
   CO(3) => W_reg_34_15_i_1_n_0,
   O(0) => x86_out_12,
   O(1) => x86_out_13,
   O(2) => x86_out_14,
   O(3) => x86_out_15
);
W_reg_34_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x86_out_16,
   R => '0',
   Q => W_reg_34_16
);
W_reg_34_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x86_out_17,
   R => '0',
   Q => W_reg_34_17
);
W_reg_34_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x86_out_18,
   R => '0',
   Q => W_reg_34_18
);
W_reg_34_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x86_out_19,
   R => '0',
   Q => W_reg_34_19
);
W_reg_34_19_i_1 : CARRY4
 port map (
   CI => W_reg_34_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_34_19_i_5_n_0,
   DI(1) => W_34_19_i_4_n_0,
   DI(2) => W_34_19_i_3_n_0,
   DI(3) => W_34_19_i_2_n_0,
   S(0) => W_34_19_i_9_n_0,
   S(1) => W_34_19_i_8_n_0,
   S(2) => W_34_19_i_7_n_0,
   S(3) => W_34_19_i_6_n_0,
   CO(0) => W_reg_34_19_i_1_n_3,
   CO(1) => W_reg_34_19_i_1_n_2,
   CO(2) => W_reg_34_19_i_1_n_1,
   CO(3) => W_reg_34_19_i_1_n_0,
   O(0) => x86_out_16,
   O(1) => x86_out_17,
   O(2) => x86_out_18,
   O(3) => x86_out_19
);
W_reg_34_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x86_out_1,
   R => '0',
   Q => W_reg_34_1
);
W_reg_34_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x86_out_20,
   R => '0',
   Q => W_reg_34_20
);
W_reg_34_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x86_out_21,
   R => '0',
   Q => W_reg_34_21
);
W_reg_34_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x86_out_22,
   R => '0',
   Q => W_reg_34_22
);
W_reg_34_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x86_out_23,
   R => '0',
   Q => W_reg_34_23
);
W_reg_34_23_i_1 : CARRY4
 port map (
   CI => W_reg_34_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_34_23_i_5_n_0,
   DI(1) => W_34_23_i_4_n_0,
   DI(2) => W_34_23_i_3_n_0,
   DI(3) => W_34_23_i_2_n_0,
   S(0) => W_34_23_i_9_n_0,
   S(1) => W_34_23_i_8_n_0,
   S(2) => W_34_23_i_7_n_0,
   S(3) => W_34_23_i_6_n_0,
   CO(0) => W_reg_34_23_i_1_n_3,
   CO(1) => W_reg_34_23_i_1_n_2,
   CO(2) => W_reg_34_23_i_1_n_1,
   CO(3) => W_reg_34_23_i_1_n_0,
   O(0) => x86_out_20,
   O(1) => x86_out_21,
   O(2) => x86_out_22,
   O(3) => x86_out_23
);
W_reg_34_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x86_out_24,
   R => '0',
   Q => W_reg_34_24
);
W_reg_34_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x86_out_25,
   R => '0',
   Q => W_reg_34_25
);
W_reg_34_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x86_out_26,
   R => '0',
   Q => W_reg_34_26
);
W_reg_34_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x86_out_27,
   R => '0',
   Q => W_reg_34_27
);
W_reg_34_27_i_1 : CARRY4
 port map (
   CI => W_reg_34_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_34_27_i_5_n_0,
   DI(1) => W_34_27_i_4_n_0,
   DI(2) => W_34_27_i_3_n_0,
   DI(3) => W_34_27_i_2_n_0,
   S(0) => W_34_27_i_9_n_0,
   S(1) => W_34_27_i_8_n_0,
   S(2) => W_34_27_i_7_n_0,
   S(3) => W_34_27_i_6_n_0,
   CO(0) => W_reg_34_27_i_1_n_3,
   CO(1) => W_reg_34_27_i_1_n_2,
   CO(2) => W_reg_34_27_i_1_n_1,
   CO(3) => W_reg_34_27_i_1_n_0,
   O(0) => x86_out_24,
   O(1) => x86_out_25,
   O(2) => x86_out_26,
   O(3) => x86_out_27
);
W_reg_34_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x86_out_28,
   R => '0',
   Q => W_reg_34_28
);
W_reg_34_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x86_out_29,
   R => '0',
   Q => W_reg_34_29
);
W_reg_34_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x86_out_2,
   R => '0',
   Q => W_reg_34_2
);
W_reg_34_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x86_out_30,
   R => '0',
   Q => W_reg_34_30
);
W_reg_34_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x86_out_31,
   R => '0',
   Q => W_reg_34_31
);
W_reg_34_31_i_1 : CARRY4
 port map (
   CI => W_reg_34_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_34_31_i_4_n_0,
   DI(1) => W_34_31_i_3_n_0,
   DI(2) => W_34_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_34_31_i_8_n_0,
   S(1) => W_34_31_i_7_n_0,
   S(2) => W_34_31_i_6_n_0,
   S(3) => W_34_31_i_5_n_0,
   CO(0) => W_reg_34_31_i_1_n_3,
   CO(1) => W_reg_34_31_i_1_n_2,
   CO(2) => W_reg_34_31_i_1_n_1,
   CO(3) => NLW_W_reg_34_31_i_1_CO_UNCONNECTED_3,
   O(0) => x86_out_28,
   O(1) => x86_out_29,
   O(2) => x86_out_30,
   O(3) => x86_out_31
);
W_reg_34_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x86_out_3,
   R => '0',
   Q => W_reg_34_3
);
W_reg_34_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_34_3_i_5_n_0,
   DI(1) => W_34_3_i_4_n_0,
   DI(2) => W_34_3_i_3_n_0,
   DI(3) => W_34_3_i_2_n_0,
   S(0) => W_34_3_i_9_n_0,
   S(1) => W_34_3_i_8_n_0,
   S(2) => W_34_3_i_7_n_0,
   S(3) => W_34_3_i_6_n_0,
   CO(0) => W_reg_34_3_i_1_n_3,
   CO(1) => W_reg_34_3_i_1_n_2,
   CO(2) => W_reg_34_3_i_1_n_1,
   CO(3) => W_reg_34_3_i_1_n_0,
   O(0) => x86_out_0,
   O(1) => x86_out_1,
   O(2) => x86_out_2,
   O(3) => x86_out_3
);
W_reg_34_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x86_out_4,
   R => '0',
   Q => W_reg_34_4
);
W_reg_34_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x86_out_5,
   R => '0',
   Q => W_reg_34_5
);
W_reg_34_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x86_out_6,
   R => '0',
   Q => W_reg_34_6
);
W_reg_34_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x86_out_7,
   R => '0',
   Q => W_reg_34_7
);
W_reg_34_7_i_1 : CARRY4
 port map (
   CI => W_reg_34_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_34_7_i_5_n_0,
   DI(1) => W_34_7_i_4_n_0,
   DI(2) => W_34_7_i_3_n_0,
   DI(3) => W_34_7_i_2_n_0,
   S(0) => W_34_7_i_9_n_0,
   S(1) => W_34_7_i_8_n_0,
   S(2) => W_34_7_i_7_n_0,
   S(3) => W_34_7_i_6_n_0,
   CO(0) => W_reg_34_7_i_1_n_3,
   CO(1) => W_reg_34_7_i_1_n_2,
   CO(2) => W_reg_34_7_i_1_n_1,
   CO(3) => W_reg_34_7_i_1_n_0,
   O(0) => x86_out_4,
   O(1) => x86_out_5,
   O(2) => x86_out_6,
   O(3) => x86_out_7
);
W_reg_34_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x86_out_8,
   R => '0',
   Q => W_reg_34_8
);
W_reg_34_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x86_out_9,
   R => '0',
   Q => W_reg_34_9
);
W_reg_35_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x83_out_0,
   R => '0',
   Q => W_reg_35_0
);
W_reg_35_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x83_out_10,
   R => '0',
   Q => W_reg_35_10
);
W_reg_35_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x83_out_11,
   R => '0',
   Q => W_reg_35_11
);
W_reg_35_11_i_1 : CARRY4
 port map (
   CI => W_reg_35_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_35_11_i_5_n_0,
   DI(1) => W_35_11_i_4_n_0,
   DI(2) => W_35_11_i_3_n_0,
   DI(3) => W_35_11_i_2_n_0,
   S(0) => W_35_11_i_9_n_0,
   S(1) => W_35_11_i_8_n_0,
   S(2) => W_35_11_i_7_n_0,
   S(3) => W_35_11_i_6_n_0,
   CO(0) => W_reg_35_11_i_1_n_3,
   CO(1) => W_reg_35_11_i_1_n_2,
   CO(2) => W_reg_35_11_i_1_n_1,
   CO(3) => W_reg_35_11_i_1_n_0,
   O(0) => x83_out_8,
   O(1) => x83_out_9,
   O(2) => x83_out_10,
   O(3) => x83_out_11
);
W_reg_35_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x83_out_12,
   R => '0',
   Q => W_reg_35_12
);
W_reg_35_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x83_out_13,
   R => '0',
   Q => W_reg_35_13
);
W_reg_35_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x83_out_14,
   R => '0',
   Q => W_reg_35_14
);
W_reg_35_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x83_out_15,
   R => '0',
   Q => W_reg_35_15
);
W_reg_35_15_i_1 : CARRY4
 port map (
   CI => W_reg_35_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_35_15_i_5_n_0,
   DI(1) => W_35_15_i_4_n_0,
   DI(2) => W_35_15_i_3_n_0,
   DI(3) => W_35_15_i_2_n_0,
   S(0) => W_35_15_i_9_n_0,
   S(1) => W_35_15_i_8_n_0,
   S(2) => W_35_15_i_7_n_0,
   S(3) => W_35_15_i_6_n_0,
   CO(0) => W_reg_35_15_i_1_n_3,
   CO(1) => W_reg_35_15_i_1_n_2,
   CO(2) => W_reg_35_15_i_1_n_1,
   CO(3) => W_reg_35_15_i_1_n_0,
   O(0) => x83_out_12,
   O(1) => x83_out_13,
   O(2) => x83_out_14,
   O(3) => x83_out_15
);
W_reg_35_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x83_out_16,
   R => '0',
   Q => W_reg_35_16
);
W_reg_35_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x83_out_17,
   R => '0',
   Q => W_reg_35_17
);
W_reg_35_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x83_out_18,
   R => '0',
   Q => W_reg_35_18
);
W_reg_35_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x83_out_19,
   R => '0',
   Q => W_reg_35_19
);
W_reg_35_19_i_1 : CARRY4
 port map (
   CI => W_reg_35_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_35_19_i_5_n_0,
   DI(1) => W_35_19_i_4_n_0,
   DI(2) => W_35_19_i_3_n_0,
   DI(3) => W_35_19_i_2_n_0,
   S(0) => W_35_19_i_9_n_0,
   S(1) => W_35_19_i_8_n_0,
   S(2) => W_35_19_i_7_n_0,
   S(3) => W_35_19_i_6_n_0,
   CO(0) => W_reg_35_19_i_1_n_3,
   CO(1) => W_reg_35_19_i_1_n_2,
   CO(2) => W_reg_35_19_i_1_n_1,
   CO(3) => W_reg_35_19_i_1_n_0,
   O(0) => x83_out_16,
   O(1) => x83_out_17,
   O(2) => x83_out_18,
   O(3) => x83_out_19
);
W_reg_35_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x83_out_1,
   R => '0',
   Q => W_reg_35_1
);
W_reg_35_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x83_out_20,
   R => '0',
   Q => W_reg_35_20
);
W_reg_35_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x83_out_21,
   R => '0',
   Q => W_reg_35_21
);
W_reg_35_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x83_out_22,
   R => '0',
   Q => W_reg_35_22
);
W_reg_35_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x83_out_23,
   R => '0',
   Q => W_reg_35_23
);
W_reg_35_23_i_1 : CARRY4
 port map (
   CI => W_reg_35_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_35_23_i_5_n_0,
   DI(1) => W_35_23_i_4_n_0,
   DI(2) => W_35_23_i_3_n_0,
   DI(3) => W_35_23_i_2_n_0,
   S(0) => W_35_23_i_9_n_0,
   S(1) => W_35_23_i_8_n_0,
   S(2) => W_35_23_i_7_n_0,
   S(3) => W_35_23_i_6_n_0,
   CO(0) => W_reg_35_23_i_1_n_3,
   CO(1) => W_reg_35_23_i_1_n_2,
   CO(2) => W_reg_35_23_i_1_n_1,
   CO(3) => W_reg_35_23_i_1_n_0,
   O(0) => x83_out_20,
   O(1) => x83_out_21,
   O(2) => x83_out_22,
   O(3) => x83_out_23
);
W_reg_35_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x83_out_24,
   R => '0',
   Q => W_reg_35_24
);
W_reg_35_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x83_out_25,
   R => '0',
   Q => W_reg_35_25
);
W_reg_35_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x83_out_26,
   R => '0',
   Q => W_reg_35_26
);
W_reg_35_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x83_out_27,
   R => '0',
   Q => W_reg_35_27
);
W_reg_35_27_i_1 : CARRY4
 port map (
   CI => W_reg_35_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_35_27_i_5_n_0,
   DI(1) => W_35_27_i_4_n_0,
   DI(2) => W_35_27_i_3_n_0,
   DI(3) => W_35_27_i_2_n_0,
   S(0) => W_35_27_i_9_n_0,
   S(1) => W_35_27_i_8_n_0,
   S(2) => W_35_27_i_7_n_0,
   S(3) => W_35_27_i_6_n_0,
   CO(0) => W_reg_35_27_i_1_n_3,
   CO(1) => W_reg_35_27_i_1_n_2,
   CO(2) => W_reg_35_27_i_1_n_1,
   CO(3) => W_reg_35_27_i_1_n_0,
   O(0) => x83_out_24,
   O(1) => x83_out_25,
   O(2) => x83_out_26,
   O(3) => x83_out_27
);
W_reg_35_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x83_out_28,
   R => '0',
   Q => W_reg_35_28
);
W_reg_35_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x83_out_29,
   R => '0',
   Q => W_reg_35_29
);
W_reg_35_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x83_out_2,
   R => '0',
   Q => W_reg_35_2
);
W_reg_35_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x83_out_30,
   R => '0',
   Q => W_reg_35_30
);
W_reg_35_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x83_out_31,
   R => '0',
   Q => W_reg_35_31
);
W_reg_35_31_i_1 : CARRY4
 port map (
   CI => W_reg_35_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_35_31_i_4_n_0,
   DI(1) => W_35_31_i_3_n_0,
   DI(2) => W_35_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_35_31_i_8_n_0,
   S(1) => W_35_31_i_7_n_0,
   S(2) => W_35_31_i_6_n_0,
   S(3) => W_35_31_i_5_n_0,
   CO(0) => W_reg_35_31_i_1_n_3,
   CO(1) => W_reg_35_31_i_1_n_2,
   CO(2) => W_reg_35_31_i_1_n_1,
   CO(3) => NLW_W_reg_35_31_i_1_CO_UNCONNECTED_3,
   O(0) => x83_out_28,
   O(1) => x83_out_29,
   O(2) => x83_out_30,
   O(3) => x83_out_31
);
W_reg_35_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x83_out_3,
   R => '0',
   Q => W_reg_35_3
);
W_reg_35_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_35_3_i_5_n_0,
   DI(1) => W_35_3_i_4_n_0,
   DI(2) => W_35_3_i_3_n_0,
   DI(3) => W_35_3_i_2_n_0,
   S(0) => W_35_3_i_9_n_0,
   S(1) => W_35_3_i_8_n_0,
   S(2) => W_35_3_i_7_n_0,
   S(3) => W_35_3_i_6_n_0,
   CO(0) => W_reg_35_3_i_1_n_3,
   CO(1) => W_reg_35_3_i_1_n_2,
   CO(2) => W_reg_35_3_i_1_n_1,
   CO(3) => W_reg_35_3_i_1_n_0,
   O(0) => x83_out_0,
   O(1) => x83_out_1,
   O(2) => x83_out_2,
   O(3) => x83_out_3
);
W_reg_35_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x83_out_4,
   R => '0',
   Q => W_reg_35_4
);
W_reg_35_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x83_out_5,
   R => '0',
   Q => W_reg_35_5
);
W_reg_35_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x83_out_6,
   R => '0',
   Q => W_reg_35_6
);
W_reg_35_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x83_out_7,
   R => '0',
   Q => W_reg_35_7
);
W_reg_35_7_i_1 : CARRY4
 port map (
   CI => W_reg_35_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_35_7_i_5_n_0,
   DI(1) => W_35_7_i_4_n_0,
   DI(2) => W_35_7_i_3_n_0,
   DI(3) => W_35_7_i_2_n_0,
   S(0) => W_35_7_i_9_n_0,
   S(1) => W_35_7_i_8_n_0,
   S(2) => W_35_7_i_7_n_0,
   S(3) => W_35_7_i_6_n_0,
   CO(0) => W_reg_35_7_i_1_n_3,
   CO(1) => W_reg_35_7_i_1_n_2,
   CO(2) => W_reg_35_7_i_1_n_1,
   CO(3) => W_reg_35_7_i_1_n_0,
   O(0) => x83_out_4,
   O(1) => x83_out_5,
   O(2) => x83_out_6,
   O(3) => x83_out_7
);
W_reg_35_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x83_out_8,
   R => '0',
   Q => W_reg_35_8
);
W_reg_35_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x83_out_9,
   R => '0',
   Q => W_reg_35_9
);
W_reg_36_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x80_out_0,
   R => '0',
   Q => W_reg_36_0
);
W_reg_36_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x80_out_10,
   R => '0',
   Q => W_reg_36_10
);
W_reg_36_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x80_out_11,
   R => '0',
   Q => W_reg_36_11
);
W_reg_36_11_i_1 : CARRY4
 port map (
   CI => W_reg_36_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_36_11_i_5_n_0,
   DI(1) => W_36_11_i_4_n_0,
   DI(2) => W_36_11_i_3_n_0,
   DI(3) => W_36_11_i_2_n_0,
   S(0) => W_36_11_i_9_n_0,
   S(1) => W_36_11_i_8_n_0,
   S(2) => W_36_11_i_7_n_0,
   S(3) => W_36_11_i_6_n_0,
   CO(0) => W_reg_36_11_i_1_n_3,
   CO(1) => W_reg_36_11_i_1_n_2,
   CO(2) => W_reg_36_11_i_1_n_1,
   CO(3) => W_reg_36_11_i_1_n_0,
   O(0) => x80_out_8,
   O(1) => x80_out_9,
   O(2) => x80_out_10,
   O(3) => x80_out_11
);
W_reg_36_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x80_out_12,
   R => '0',
   Q => W_reg_36_12
);
W_reg_36_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x80_out_13,
   R => '0',
   Q => W_reg_36_13
);
W_reg_36_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x80_out_14,
   R => '0',
   Q => W_reg_36_14
);
W_reg_36_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x80_out_15,
   R => '0',
   Q => W_reg_36_15
);
W_reg_36_15_i_1 : CARRY4
 port map (
   CI => W_reg_36_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_36_15_i_5_n_0,
   DI(1) => W_36_15_i_4_n_0,
   DI(2) => W_36_15_i_3_n_0,
   DI(3) => W_36_15_i_2_n_0,
   S(0) => W_36_15_i_9_n_0,
   S(1) => W_36_15_i_8_n_0,
   S(2) => W_36_15_i_7_n_0,
   S(3) => W_36_15_i_6_n_0,
   CO(0) => W_reg_36_15_i_1_n_3,
   CO(1) => W_reg_36_15_i_1_n_2,
   CO(2) => W_reg_36_15_i_1_n_1,
   CO(3) => W_reg_36_15_i_1_n_0,
   O(0) => x80_out_12,
   O(1) => x80_out_13,
   O(2) => x80_out_14,
   O(3) => x80_out_15
);
W_reg_36_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x80_out_16,
   R => '0',
   Q => W_reg_36_16
);
W_reg_36_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x80_out_17,
   R => '0',
   Q => W_reg_36_17
);
W_reg_36_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x80_out_18,
   R => '0',
   Q => W_reg_36_18
);
W_reg_36_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x80_out_19,
   R => '0',
   Q => W_reg_36_19
);
W_reg_36_19_i_1 : CARRY4
 port map (
   CI => W_reg_36_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_36_19_i_5_n_0,
   DI(1) => W_36_19_i_4_n_0,
   DI(2) => W_36_19_i_3_n_0,
   DI(3) => W_36_19_i_2_n_0,
   S(0) => W_36_19_i_9_n_0,
   S(1) => W_36_19_i_8_n_0,
   S(2) => W_36_19_i_7_n_0,
   S(3) => W_36_19_i_6_n_0,
   CO(0) => W_reg_36_19_i_1_n_3,
   CO(1) => W_reg_36_19_i_1_n_2,
   CO(2) => W_reg_36_19_i_1_n_1,
   CO(3) => W_reg_36_19_i_1_n_0,
   O(0) => x80_out_16,
   O(1) => x80_out_17,
   O(2) => x80_out_18,
   O(3) => x80_out_19
);
W_reg_36_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x80_out_1,
   R => '0',
   Q => W_reg_36_1
);
W_reg_36_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x80_out_20,
   R => '0',
   Q => W_reg_36_20
);
W_reg_36_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x80_out_21,
   R => '0',
   Q => W_reg_36_21
);
W_reg_36_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x80_out_22,
   R => '0',
   Q => W_reg_36_22
);
W_reg_36_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x80_out_23,
   R => '0',
   Q => W_reg_36_23
);
W_reg_36_23_i_1 : CARRY4
 port map (
   CI => W_reg_36_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_36_23_i_5_n_0,
   DI(1) => W_36_23_i_4_n_0,
   DI(2) => W_36_23_i_3_n_0,
   DI(3) => W_36_23_i_2_n_0,
   S(0) => W_36_23_i_9_n_0,
   S(1) => W_36_23_i_8_n_0,
   S(2) => W_36_23_i_7_n_0,
   S(3) => W_36_23_i_6_n_0,
   CO(0) => W_reg_36_23_i_1_n_3,
   CO(1) => W_reg_36_23_i_1_n_2,
   CO(2) => W_reg_36_23_i_1_n_1,
   CO(3) => W_reg_36_23_i_1_n_0,
   O(0) => x80_out_20,
   O(1) => x80_out_21,
   O(2) => x80_out_22,
   O(3) => x80_out_23
);
W_reg_36_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x80_out_24,
   R => '0',
   Q => W_reg_36_24
);
W_reg_36_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x80_out_25,
   R => '0',
   Q => W_reg_36_25
);
W_reg_36_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x80_out_26,
   R => '0',
   Q => W_reg_36_26
);
W_reg_36_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x80_out_27,
   R => '0',
   Q => W_reg_36_27
);
W_reg_36_27_i_1 : CARRY4
 port map (
   CI => W_reg_36_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_36_27_i_5_n_0,
   DI(1) => W_36_27_i_4_n_0,
   DI(2) => W_36_27_i_3_n_0,
   DI(3) => W_36_27_i_2_n_0,
   S(0) => W_36_27_i_9_n_0,
   S(1) => W_36_27_i_8_n_0,
   S(2) => W_36_27_i_7_n_0,
   S(3) => W_36_27_i_6_n_0,
   CO(0) => W_reg_36_27_i_1_n_3,
   CO(1) => W_reg_36_27_i_1_n_2,
   CO(2) => W_reg_36_27_i_1_n_1,
   CO(3) => W_reg_36_27_i_1_n_0,
   O(0) => x80_out_24,
   O(1) => x80_out_25,
   O(2) => x80_out_26,
   O(3) => x80_out_27
);
W_reg_36_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x80_out_28,
   R => '0',
   Q => W_reg_36_28
);
W_reg_36_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x80_out_29,
   R => '0',
   Q => W_reg_36_29
);
W_reg_36_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x80_out_2,
   R => '0',
   Q => W_reg_36_2
);
W_reg_36_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x80_out_30,
   R => '0',
   Q => W_reg_36_30
);
W_reg_36_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x80_out_31,
   R => '0',
   Q => W_reg_36_31
);
W_reg_36_31_i_1 : CARRY4
 port map (
   CI => W_reg_36_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_36_31_i_4_n_0,
   DI(1) => W_36_31_i_3_n_0,
   DI(2) => W_36_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_36_31_i_8_n_0,
   S(1) => W_36_31_i_7_n_0,
   S(2) => W_36_31_i_6_n_0,
   S(3) => W_36_31_i_5_n_0,
   CO(0) => W_reg_36_31_i_1_n_3,
   CO(1) => W_reg_36_31_i_1_n_2,
   CO(2) => W_reg_36_31_i_1_n_1,
   CO(3) => NLW_W_reg_36_31_i_1_CO_UNCONNECTED_3,
   O(0) => x80_out_28,
   O(1) => x80_out_29,
   O(2) => x80_out_30,
   O(3) => x80_out_31
);
W_reg_36_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x80_out_3,
   R => '0',
   Q => W_reg_36_3
);
W_reg_36_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_36_3_i_5_n_0,
   DI(1) => W_36_3_i_4_n_0,
   DI(2) => W_36_3_i_3_n_0,
   DI(3) => W_36_3_i_2_n_0,
   S(0) => W_36_3_i_9_n_0,
   S(1) => W_36_3_i_8_n_0,
   S(2) => W_36_3_i_7_n_0,
   S(3) => W_36_3_i_6_n_0,
   CO(0) => W_reg_36_3_i_1_n_3,
   CO(1) => W_reg_36_3_i_1_n_2,
   CO(2) => W_reg_36_3_i_1_n_1,
   CO(3) => W_reg_36_3_i_1_n_0,
   O(0) => x80_out_0,
   O(1) => x80_out_1,
   O(2) => x80_out_2,
   O(3) => x80_out_3
);
W_reg_36_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x80_out_4,
   R => '0',
   Q => W_reg_36_4
);
W_reg_36_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x80_out_5,
   R => '0',
   Q => W_reg_36_5
);
W_reg_36_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x80_out_6,
   R => '0',
   Q => W_reg_36_6
);
W_reg_36_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x80_out_7,
   R => '0',
   Q => W_reg_36_7
);
W_reg_36_7_i_1 : CARRY4
 port map (
   CI => W_reg_36_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_36_7_i_5_n_0,
   DI(1) => W_36_7_i_4_n_0,
   DI(2) => W_36_7_i_3_n_0,
   DI(3) => W_36_7_i_2_n_0,
   S(0) => W_36_7_i_9_n_0,
   S(1) => W_36_7_i_8_n_0,
   S(2) => W_36_7_i_7_n_0,
   S(3) => W_36_7_i_6_n_0,
   CO(0) => W_reg_36_7_i_1_n_3,
   CO(1) => W_reg_36_7_i_1_n_2,
   CO(2) => W_reg_36_7_i_1_n_1,
   CO(3) => W_reg_36_7_i_1_n_0,
   O(0) => x80_out_4,
   O(1) => x80_out_5,
   O(2) => x80_out_6,
   O(3) => x80_out_7
);
W_reg_36_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x80_out_8,
   R => '0',
   Q => W_reg_36_8
);
W_reg_36_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x80_out_9,
   R => '0',
   Q => W_reg_36_9
);
W_reg_37_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x77_out_0,
   R => '0',
   Q => W_reg_37_0
);
W_reg_37_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x77_out_10,
   R => '0',
   Q => W_reg_37_10
);
W_reg_37_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x77_out_11,
   R => '0',
   Q => W_reg_37_11
);
W_reg_37_11_i_1 : CARRY4
 port map (
   CI => W_reg_37_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_37_11_i_5_n_0,
   DI(1) => W_37_11_i_4_n_0,
   DI(2) => W_37_11_i_3_n_0,
   DI(3) => W_37_11_i_2_n_0,
   S(0) => W_37_11_i_9_n_0,
   S(1) => W_37_11_i_8_n_0,
   S(2) => W_37_11_i_7_n_0,
   S(3) => W_37_11_i_6_n_0,
   CO(0) => W_reg_37_11_i_1_n_3,
   CO(1) => W_reg_37_11_i_1_n_2,
   CO(2) => W_reg_37_11_i_1_n_1,
   CO(3) => W_reg_37_11_i_1_n_0,
   O(0) => x77_out_8,
   O(1) => x77_out_9,
   O(2) => x77_out_10,
   O(3) => x77_out_11
);
W_reg_37_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x77_out_12,
   R => '0',
   Q => W_reg_37_12
);
W_reg_37_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x77_out_13,
   R => '0',
   Q => W_reg_37_13
);
W_reg_37_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x77_out_14,
   R => '0',
   Q => W_reg_37_14
);
W_reg_37_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x77_out_15,
   R => '0',
   Q => W_reg_37_15
);
W_reg_37_15_i_1 : CARRY4
 port map (
   CI => W_reg_37_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_37_15_i_5_n_0,
   DI(1) => W_37_15_i_4_n_0,
   DI(2) => W_37_15_i_3_n_0,
   DI(3) => W_37_15_i_2_n_0,
   S(0) => W_37_15_i_9_n_0,
   S(1) => W_37_15_i_8_n_0,
   S(2) => W_37_15_i_7_n_0,
   S(3) => W_37_15_i_6_n_0,
   CO(0) => W_reg_37_15_i_1_n_3,
   CO(1) => W_reg_37_15_i_1_n_2,
   CO(2) => W_reg_37_15_i_1_n_1,
   CO(3) => W_reg_37_15_i_1_n_0,
   O(0) => x77_out_12,
   O(1) => x77_out_13,
   O(2) => x77_out_14,
   O(3) => x77_out_15
);
W_reg_37_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x77_out_16,
   R => '0',
   Q => W_reg_37_16
);
W_reg_37_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x77_out_17,
   R => '0',
   Q => W_reg_37_17
);
W_reg_37_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x77_out_18,
   R => '0',
   Q => W_reg_37_18
);
W_reg_37_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x77_out_19,
   R => '0',
   Q => W_reg_37_19
);
W_reg_37_19_i_1 : CARRY4
 port map (
   CI => W_reg_37_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_37_19_i_5_n_0,
   DI(1) => W_37_19_i_4_n_0,
   DI(2) => W_37_19_i_3_n_0,
   DI(3) => W_37_19_i_2_n_0,
   S(0) => W_37_19_i_9_n_0,
   S(1) => W_37_19_i_8_n_0,
   S(2) => W_37_19_i_7_n_0,
   S(3) => W_37_19_i_6_n_0,
   CO(0) => W_reg_37_19_i_1_n_3,
   CO(1) => W_reg_37_19_i_1_n_2,
   CO(2) => W_reg_37_19_i_1_n_1,
   CO(3) => W_reg_37_19_i_1_n_0,
   O(0) => x77_out_16,
   O(1) => x77_out_17,
   O(2) => x77_out_18,
   O(3) => x77_out_19
);
W_reg_37_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x77_out_1,
   R => '0',
   Q => W_reg_37_1
);
W_reg_37_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x77_out_20,
   R => '0',
   Q => W_reg_37_20
);
W_reg_37_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x77_out_21,
   R => '0',
   Q => W_reg_37_21
);
W_reg_37_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x77_out_22,
   R => '0',
   Q => W_reg_37_22
);
W_reg_37_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x77_out_23,
   R => '0',
   Q => W_reg_37_23
);
W_reg_37_23_i_1 : CARRY4
 port map (
   CI => W_reg_37_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_37_23_i_5_n_0,
   DI(1) => W_37_23_i_4_n_0,
   DI(2) => W_37_23_i_3_n_0,
   DI(3) => W_37_23_i_2_n_0,
   S(0) => W_37_23_i_9_n_0,
   S(1) => W_37_23_i_8_n_0,
   S(2) => W_37_23_i_7_n_0,
   S(3) => W_37_23_i_6_n_0,
   CO(0) => W_reg_37_23_i_1_n_3,
   CO(1) => W_reg_37_23_i_1_n_2,
   CO(2) => W_reg_37_23_i_1_n_1,
   CO(3) => W_reg_37_23_i_1_n_0,
   O(0) => x77_out_20,
   O(1) => x77_out_21,
   O(2) => x77_out_22,
   O(3) => x77_out_23
);
W_reg_37_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x77_out_24,
   R => '0',
   Q => W_reg_37_24
);
W_reg_37_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x77_out_25,
   R => '0',
   Q => W_reg_37_25
);
W_reg_37_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x77_out_26,
   R => '0',
   Q => W_reg_37_26
);
W_reg_37_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x77_out_27,
   R => '0',
   Q => W_reg_37_27
);
W_reg_37_27_i_1 : CARRY4
 port map (
   CI => W_reg_37_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_37_27_i_5_n_0,
   DI(1) => W_37_27_i_4_n_0,
   DI(2) => W_37_27_i_3_n_0,
   DI(3) => W_37_27_i_2_n_0,
   S(0) => W_37_27_i_9_n_0,
   S(1) => W_37_27_i_8_n_0,
   S(2) => W_37_27_i_7_n_0,
   S(3) => W_37_27_i_6_n_0,
   CO(0) => W_reg_37_27_i_1_n_3,
   CO(1) => W_reg_37_27_i_1_n_2,
   CO(2) => W_reg_37_27_i_1_n_1,
   CO(3) => W_reg_37_27_i_1_n_0,
   O(0) => x77_out_24,
   O(1) => x77_out_25,
   O(2) => x77_out_26,
   O(3) => x77_out_27
);
W_reg_37_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x77_out_28,
   R => '0',
   Q => W_reg_37_28
);
W_reg_37_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x77_out_29,
   R => '0',
   Q => W_reg_37_29
);
W_reg_37_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x77_out_2,
   R => '0',
   Q => W_reg_37_2
);
W_reg_37_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x77_out_30,
   R => '0',
   Q => W_reg_37_30
);
W_reg_37_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x77_out_31,
   R => '0',
   Q => W_reg_37_31
);
W_reg_37_31_i_1 : CARRY4
 port map (
   CI => W_reg_37_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_37_31_i_4_n_0,
   DI(1) => W_37_31_i_3_n_0,
   DI(2) => W_37_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_37_31_i_8_n_0,
   S(1) => W_37_31_i_7_n_0,
   S(2) => W_37_31_i_6_n_0,
   S(3) => W_37_31_i_5_n_0,
   CO(0) => W_reg_37_31_i_1_n_3,
   CO(1) => W_reg_37_31_i_1_n_2,
   CO(2) => W_reg_37_31_i_1_n_1,
   CO(3) => NLW_W_reg_37_31_i_1_CO_UNCONNECTED_3,
   O(0) => x77_out_28,
   O(1) => x77_out_29,
   O(2) => x77_out_30,
   O(3) => x77_out_31
);
W_reg_37_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x77_out_3,
   R => '0',
   Q => W_reg_37_3
);
W_reg_37_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_37_3_i_5_n_0,
   DI(1) => W_37_3_i_4_n_0,
   DI(2) => W_37_3_i_3_n_0,
   DI(3) => W_37_3_i_2_n_0,
   S(0) => W_37_3_i_9_n_0,
   S(1) => W_37_3_i_8_n_0,
   S(2) => W_37_3_i_7_n_0,
   S(3) => W_37_3_i_6_n_0,
   CO(0) => W_reg_37_3_i_1_n_3,
   CO(1) => W_reg_37_3_i_1_n_2,
   CO(2) => W_reg_37_3_i_1_n_1,
   CO(3) => W_reg_37_3_i_1_n_0,
   O(0) => x77_out_0,
   O(1) => x77_out_1,
   O(2) => x77_out_2,
   O(3) => x77_out_3
);
W_reg_37_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x77_out_4,
   R => '0',
   Q => W_reg_37_4
);
W_reg_37_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x77_out_5,
   R => '0',
   Q => W_reg_37_5
);
W_reg_37_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x77_out_6,
   R => '0',
   Q => W_reg_37_6
);
W_reg_37_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x77_out_7,
   R => '0',
   Q => W_reg_37_7
);
W_reg_37_7_i_1 : CARRY4
 port map (
   CI => W_reg_37_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_37_7_i_5_n_0,
   DI(1) => W_37_7_i_4_n_0,
   DI(2) => W_37_7_i_3_n_0,
   DI(3) => W_37_7_i_2_n_0,
   S(0) => W_37_7_i_9_n_0,
   S(1) => W_37_7_i_8_n_0,
   S(2) => W_37_7_i_7_n_0,
   S(3) => W_37_7_i_6_n_0,
   CO(0) => W_reg_37_7_i_1_n_3,
   CO(1) => W_reg_37_7_i_1_n_2,
   CO(2) => W_reg_37_7_i_1_n_1,
   CO(3) => W_reg_37_7_i_1_n_0,
   O(0) => x77_out_4,
   O(1) => x77_out_5,
   O(2) => x77_out_6,
   O(3) => x77_out_7
);
W_reg_37_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x77_out_8,
   R => '0',
   Q => W_reg_37_8
);
W_reg_37_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x77_out_9,
   R => '0',
   Q => W_reg_37_9
);
W_reg_38_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x74_out_0,
   R => '0',
   Q => W_reg_38_0
);
W_reg_38_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x74_out_10,
   R => '0',
   Q => W_reg_38_10
);
W_reg_38_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x74_out_11,
   R => '0',
   Q => W_reg_38_11
);
W_reg_38_11_i_1 : CARRY4
 port map (
   CI => W_reg_38_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_38_11_i_5_n_0,
   DI(1) => W_38_11_i_4_n_0,
   DI(2) => W_38_11_i_3_n_0,
   DI(3) => W_38_11_i_2_n_0,
   S(0) => W_38_11_i_9_n_0,
   S(1) => W_38_11_i_8_n_0,
   S(2) => W_38_11_i_7_n_0,
   S(3) => W_38_11_i_6_n_0,
   CO(0) => W_reg_38_11_i_1_n_3,
   CO(1) => W_reg_38_11_i_1_n_2,
   CO(2) => W_reg_38_11_i_1_n_1,
   CO(3) => W_reg_38_11_i_1_n_0,
   O(0) => x74_out_8,
   O(1) => x74_out_9,
   O(2) => x74_out_10,
   O(3) => x74_out_11
);
W_reg_38_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x74_out_12,
   R => '0',
   Q => W_reg_38_12
);
W_reg_38_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x74_out_13,
   R => '0',
   Q => W_reg_38_13
);
W_reg_38_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x74_out_14,
   R => '0',
   Q => W_reg_38_14
);
W_reg_38_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x74_out_15,
   R => '0',
   Q => W_reg_38_15
);
W_reg_38_15_i_1 : CARRY4
 port map (
   CI => W_reg_38_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_38_15_i_5_n_0,
   DI(1) => W_38_15_i_4_n_0,
   DI(2) => W_38_15_i_3_n_0,
   DI(3) => W_38_15_i_2_n_0,
   S(0) => W_38_15_i_9_n_0,
   S(1) => W_38_15_i_8_n_0,
   S(2) => W_38_15_i_7_n_0,
   S(3) => W_38_15_i_6_n_0,
   CO(0) => W_reg_38_15_i_1_n_3,
   CO(1) => W_reg_38_15_i_1_n_2,
   CO(2) => W_reg_38_15_i_1_n_1,
   CO(3) => W_reg_38_15_i_1_n_0,
   O(0) => x74_out_12,
   O(1) => x74_out_13,
   O(2) => x74_out_14,
   O(3) => x74_out_15
);
W_reg_38_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x74_out_16,
   R => '0',
   Q => W_reg_38_16
);
W_reg_38_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x74_out_17,
   R => '0',
   Q => W_reg_38_17
);
W_reg_38_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x74_out_18,
   R => '0',
   Q => W_reg_38_18
);
W_reg_38_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x74_out_19,
   R => '0',
   Q => W_reg_38_19
);
W_reg_38_19_i_1 : CARRY4
 port map (
   CI => W_reg_38_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_38_19_i_5_n_0,
   DI(1) => W_38_19_i_4_n_0,
   DI(2) => W_38_19_i_3_n_0,
   DI(3) => W_38_19_i_2_n_0,
   S(0) => W_38_19_i_9_n_0,
   S(1) => W_38_19_i_8_n_0,
   S(2) => W_38_19_i_7_n_0,
   S(3) => W_38_19_i_6_n_0,
   CO(0) => W_reg_38_19_i_1_n_3,
   CO(1) => W_reg_38_19_i_1_n_2,
   CO(2) => W_reg_38_19_i_1_n_1,
   CO(3) => W_reg_38_19_i_1_n_0,
   O(0) => x74_out_16,
   O(1) => x74_out_17,
   O(2) => x74_out_18,
   O(3) => x74_out_19
);
W_reg_38_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x74_out_1,
   R => '0',
   Q => W_reg_38_1
);
W_reg_38_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x74_out_20,
   R => '0',
   Q => W_reg_38_20
);
W_reg_38_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x74_out_21,
   R => '0',
   Q => W_reg_38_21
);
W_reg_38_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x74_out_22,
   R => '0',
   Q => W_reg_38_22
);
W_reg_38_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x74_out_23,
   R => '0',
   Q => W_reg_38_23
);
W_reg_38_23_i_1 : CARRY4
 port map (
   CI => W_reg_38_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_38_23_i_5_n_0,
   DI(1) => W_38_23_i_4_n_0,
   DI(2) => W_38_23_i_3_n_0,
   DI(3) => W_38_23_i_2_n_0,
   S(0) => W_38_23_i_9_n_0,
   S(1) => W_38_23_i_8_n_0,
   S(2) => W_38_23_i_7_n_0,
   S(3) => W_38_23_i_6_n_0,
   CO(0) => W_reg_38_23_i_1_n_3,
   CO(1) => W_reg_38_23_i_1_n_2,
   CO(2) => W_reg_38_23_i_1_n_1,
   CO(3) => W_reg_38_23_i_1_n_0,
   O(0) => x74_out_20,
   O(1) => x74_out_21,
   O(2) => x74_out_22,
   O(3) => x74_out_23
);
W_reg_38_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x74_out_24,
   R => '0',
   Q => W_reg_38_24
);
W_reg_38_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x74_out_25,
   R => '0',
   Q => W_reg_38_25
);
W_reg_38_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x74_out_26,
   R => '0',
   Q => W_reg_38_26
);
W_reg_38_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x74_out_27,
   R => '0',
   Q => W_reg_38_27
);
W_reg_38_27_i_1 : CARRY4
 port map (
   CI => W_reg_38_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_38_27_i_5_n_0,
   DI(1) => W_38_27_i_4_n_0,
   DI(2) => W_38_27_i_3_n_0,
   DI(3) => W_38_27_i_2_n_0,
   S(0) => W_38_27_i_9_n_0,
   S(1) => W_38_27_i_8_n_0,
   S(2) => W_38_27_i_7_n_0,
   S(3) => W_38_27_i_6_n_0,
   CO(0) => W_reg_38_27_i_1_n_3,
   CO(1) => W_reg_38_27_i_1_n_2,
   CO(2) => W_reg_38_27_i_1_n_1,
   CO(3) => W_reg_38_27_i_1_n_0,
   O(0) => x74_out_24,
   O(1) => x74_out_25,
   O(2) => x74_out_26,
   O(3) => x74_out_27
);
W_reg_38_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x74_out_28,
   R => '0',
   Q => W_reg_38_28
);
W_reg_38_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x74_out_29,
   R => '0',
   Q => W_reg_38_29
);
W_reg_38_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x74_out_2,
   R => '0',
   Q => W_reg_38_2
);
W_reg_38_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x74_out_30,
   R => '0',
   Q => W_reg_38_30
);
W_reg_38_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x74_out_31,
   R => '0',
   Q => W_reg_38_31
);
W_reg_38_31_i_1 : CARRY4
 port map (
   CI => W_reg_38_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_38_31_i_4_n_0,
   DI(1) => W_38_31_i_3_n_0,
   DI(2) => W_38_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_38_31_i_8_n_0,
   S(1) => W_38_31_i_7_n_0,
   S(2) => W_38_31_i_6_n_0,
   S(3) => W_38_31_i_5_n_0,
   CO(0) => W_reg_38_31_i_1_n_3,
   CO(1) => W_reg_38_31_i_1_n_2,
   CO(2) => W_reg_38_31_i_1_n_1,
   CO(3) => NLW_W_reg_38_31_i_1_CO_UNCONNECTED_3,
   O(0) => x74_out_28,
   O(1) => x74_out_29,
   O(2) => x74_out_30,
   O(3) => x74_out_31
);
W_reg_38_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x74_out_3,
   R => '0',
   Q => W_reg_38_3
);
W_reg_38_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_38_3_i_5_n_0,
   DI(1) => W_38_3_i_4_n_0,
   DI(2) => W_38_3_i_3_n_0,
   DI(3) => W_38_3_i_2_n_0,
   S(0) => W_38_3_i_9_n_0,
   S(1) => W_38_3_i_8_n_0,
   S(2) => W_38_3_i_7_n_0,
   S(3) => W_38_3_i_6_n_0,
   CO(0) => W_reg_38_3_i_1_n_3,
   CO(1) => W_reg_38_3_i_1_n_2,
   CO(2) => W_reg_38_3_i_1_n_1,
   CO(3) => W_reg_38_3_i_1_n_0,
   O(0) => x74_out_0,
   O(1) => x74_out_1,
   O(2) => x74_out_2,
   O(3) => x74_out_3
);
W_reg_38_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x74_out_4,
   R => '0',
   Q => W_reg_38_4
);
W_reg_38_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x74_out_5,
   R => '0',
   Q => W_reg_38_5
);
W_reg_38_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x74_out_6,
   R => '0',
   Q => W_reg_38_6
);
W_reg_38_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x74_out_7,
   R => '0',
   Q => W_reg_38_7
);
W_reg_38_7_i_1 : CARRY4
 port map (
   CI => W_reg_38_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_38_7_i_5_n_0,
   DI(1) => W_38_7_i_4_n_0,
   DI(2) => W_38_7_i_3_n_0,
   DI(3) => W_38_7_i_2_n_0,
   S(0) => W_38_7_i_9_n_0,
   S(1) => W_38_7_i_8_n_0,
   S(2) => W_38_7_i_7_n_0,
   S(3) => W_38_7_i_6_n_0,
   CO(0) => W_reg_38_7_i_1_n_3,
   CO(1) => W_reg_38_7_i_1_n_2,
   CO(2) => W_reg_38_7_i_1_n_1,
   CO(3) => W_reg_38_7_i_1_n_0,
   O(0) => x74_out_4,
   O(1) => x74_out_5,
   O(2) => x74_out_6,
   O(3) => x74_out_7
);
W_reg_38_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x74_out_8,
   R => '0',
   Q => W_reg_38_8
);
W_reg_38_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x74_out_9,
   R => '0',
   Q => W_reg_38_9
);
W_reg_39_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x71_out_0,
   R => '0',
   Q => W_reg_39_0
);
W_reg_39_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x71_out_10,
   R => '0',
   Q => W_reg_39_10
);
W_reg_39_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x71_out_11,
   R => '0',
   Q => W_reg_39_11
);
W_reg_39_11_i_1 : CARRY4
 port map (
   CI => W_reg_39_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_39_11_i_5_n_0,
   DI(1) => W_39_11_i_4_n_0,
   DI(2) => W_39_11_i_3_n_0,
   DI(3) => W_39_11_i_2_n_0,
   S(0) => W_39_11_i_9_n_0,
   S(1) => W_39_11_i_8_n_0,
   S(2) => W_39_11_i_7_n_0,
   S(3) => W_39_11_i_6_n_0,
   CO(0) => W_reg_39_11_i_1_n_3,
   CO(1) => W_reg_39_11_i_1_n_2,
   CO(2) => W_reg_39_11_i_1_n_1,
   CO(3) => W_reg_39_11_i_1_n_0,
   O(0) => x71_out_8,
   O(1) => x71_out_9,
   O(2) => x71_out_10,
   O(3) => x71_out_11
);
W_reg_39_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x71_out_12,
   R => '0',
   Q => W_reg_39_12
);
W_reg_39_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x71_out_13,
   R => '0',
   Q => W_reg_39_13
);
W_reg_39_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x71_out_14,
   R => '0',
   Q => W_reg_39_14
);
W_reg_39_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x71_out_15,
   R => '0',
   Q => W_reg_39_15
);
W_reg_39_15_i_1 : CARRY4
 port map (
   CI => W_reg_39_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_39_15_i_5_n_0,
   DI(1) => W_39_15_i_4_n_0,
   DI(2) => W_39_15_i_3_n_0,
   DI(3) => W_39_15_i_2_n_0,
   S(0) => W_39_15_i_9_n_0,
   S(1) => W_39_15_i_8_n_0,
   S(2) => W_39_15_i_7_n_0,
   S(3) => W_39_15_i_6_n_0,
   CO(0) => W_reg_39_15_i_1_n_3,
   CO(1) => W_reg_39_15_i_1_n_2,
   CO(2) => W_reg_39_15_i_1_n_1,
   CO(3) => W_reg_39_15_i_1_n_0,
   O(0) => x71_out_12,
   O(1) => x71_out_13,
   O(2) => x71_out_14,
   O(3) => x71_out_15
);
W_reg_39_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x71_out_16,
   R => '0',
   Q => W_reg_39_16
);
W_reg_39_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x71_out_17,
   R => '0',
   Q => W_reg_39_17
);
W_reg_39_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x71_out_18,
   R => '0',
   Q => W_reg_39_18
);
W_reg_39_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x71_out_19,
   R => '0',
   Q => W_reg_39_19
);
W_reg_39_19_i_1 : CARRY4
 port map (
   CI => W_reg_39_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_39_19_i_5_n_0,
   DI(1) => W_39_19_i_4_n_0,
   DI(2) => W_39_19_i_3_n_0,
   DI(3) => W_39_19_i_2_n_0,
   S(0) => W_39_19_i_9_n_0,
   S(1) => W_39_19_i_8_n_0,
   S(2) => W_39_19_i_7_n_0,
   S(3) => W_39_19_i_6_n_0,
   CO(0) => W_reg_39_19_i_1_n_3,
   CO(1) => W_reg_39_19_i_1_n_2,
   CO(2) => W_reg_39_19_i_1_n_1,
   CO(3) => W_reg_39_19_i_1_n_0,
   O(0) => x71_out_16,
   O(1) => x71_out_17,
   O(2) => x71_out_18,
   O(3) => x71_out_19
);
W_reg_39_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x71_out_1,
   R => '0',
   Q => W_reg_39_1
);
W_reg_39_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x71_out_20,
   R => '0',
   Q => W_reg_39_20
);
W_reg_39_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x71_out_21,
   R => '0',
   Q => W_reg_39_21
);
W_reg_39_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x71_out_22,
   R => '0',
   Q => W_reg_39_22
);
W_reg_39_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x71_out_23,
   R => '0',
   Q => W_reg_39_23
);
W_reg_39_23_i_1 : CARRY4
 port map (
   CI => W_reg_39_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_39_23_i_5_n_0,
   DI(1) => W_39_23_i_4_n_0,
   DI(2) => W_39_23_i_3_n_0,
   DI(3) => W_39_23_i_2_n_0,
   S(0) => W_39_23_i_9_n_0,
   S(1) => W_39_23_i_8_n_0,
   S(2) => W_39_23_i_7_n_0,
   S(3) => W_39_23_i_6_n_0,
   CO(0) => W_reg_39_23_i_1_n_3,
   CO(1) => W_reg_39_23_i_1_n_2,
   CO(2) => W_reg_39_23_i_1_n_1,
   CO(3) => W_reg_39_23_i_1_n_0,
   O(0) => x71_out_20,
   O(1) => x71_out_21,
   O(2) => x71_out_22,
   O(3) => x71_out_23
);
W_reg_39_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x71_out_24,
   R => '0',
   Q => W_reg_39_24
);
W_reg_39_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x71_out_25,
   R => '0',
   Q => W_reg_39_25
);
W_reg_39_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x71_out_26,
   R => '0',
   Q => W_reg_39_26
);
W_reg_39_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x71_out_27,
   R => '0',
   Q => W_reg_39_27
);
W_reg_39_27_i_1 : CARRY4
 port map (
   CI => W_reg_39_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_39_27_i_5_n_0,
   DI(1) => W_39_27_i_4_n_0,
   DI(2) => W_39_27_i_3_n_0,
   DI(3) => W_39_27_i_2_n_0,
   S(0) => W_39_27_i_9_n_0,
   S(1) => W_39_27_i_8_n_0,
   S(2) => W_39_27_i_7_n_0,
   S(3) => W_39_27_i_6_n_0,
   CO(0) => W_reg_39_27_i_1_n_3,
   CO(1) => W_reg_39_27_i_1_n_2,
   CO(2) => W_reg_39_27_i_1_n_1,
   CO(3) => W_reg_39_27_i_1_n_0,
   O(0) => x71_out_24,
   O(1) => x71_out_25,
   O(2) => x71_out_26,
   O(3) => x71_out_27
);
W_reg_39_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x71_out_28,
   R => '0',
   Q => W_reg_39_28
);
W_reg_39_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x71_out_29,
   R => '0',
   Q => W_reg_39_29
);
W_reg_39_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x71_out_2,
   R => '0',
   Q => W_reg_39_2
);
W_reg_39_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x71_out_30,
   R => '0',
   Q => W_reg_39_30
);
W_reg_39_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x71_out_31,
   R => '0',
   Q => W_reg_39_31
);
W_reg_39_31_i_1 : CARRY4
 port map (
   CI => W_reg_39_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_39_31_i_4_n_0,
   DI(1) => W_39_31_i_3_n_0,
   DI(2) => W_39_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_39_31_i_8_n_0,
   S(1) => W_39_31_i_7_n_0,
   S(2) => W_39_31_i_6_n_0,
   S(3) => W_39_31_i_5_n_0,
   CO(0) => W_reg_39_31_i_1_n_3,
   CO(1) => W_reg_39_31_i_1_n_2,
   CO(2) => W_reg_39_31_i_1_n_1,
   CO(3) => NLW_W_reg_39_31_i_1_CO_UNCONNECTED_3,
   O(0) => x71_out_28,
   O(1) => x71_out_29,
   O(2) => x71_out_30,
   O(3) => x71_out_31
);
W_reg_39_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x71_out_3,
   R => '0',
   Q => W_reg_39_3
);
W_reg_39_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_39_3_i_5_n_0,
   DI(1) => W_39_3_i_4_n_0,
   DI(2) => W_39_3_i_3_n_0,
   DI(3) => W_39_3_i_2_n_0,
   S(0) => W_39_3_i_9_n_0,
   S(1) => W_39_3_i_8_n_0,
   S(2) => W_39_3_i_7_n_0,
   S(3) => W_39_3_i_6_n_0,
   CO(0) => W_reg_39_3_i_1_n_3,
   CO(1) => W_reg_39_3_i_1_n_2,
   CO(2) => W_reg_39_3_i_1_n_1,
   CO(3) => W_reg_39_3_i_1_n_0,
   O(0) => x71_out_0,
   O(1) => x71_out_1,
   O(2) => x71_out_2,
   O(3) => x71_out_3
);
W_reg_39_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x71_out_4,
   R => '0',
   Q => W_reg_39_4
);
W_reg_39_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x71_out_5,
   R => '0',
   Q => W_reg_39_5
);
W_reg_39_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x71_out_6,
   R => '0',
   Q => W_reg_39_6
);
W_reg_39_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x71_out_7,
   R => '0',
   Q => W_reg_39_7
);
W_reg_39_7_i_1 : CARRY4
 port map (
   CI => W_reg_39_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_39_7_i_5_n_0,
   DI(1) => W_39_7_i_4_n_0,
   DI(2) => W_39_7_i_3_n_0,
   DI(3) => W_39_7_i_2_n_0,
   S(0) => W_39_7_i_9_n_0,
   S(1) => W_39_7_i_8_n_0,
   S(2) => W_39_7_i_7_n_0,
   S(3) => W_39_7_i_6_n_0,
   CO(0) => W_reg_39_7_i_1_n_3,
   CO(1) => W_reg_39_7_i_1_n_2,
   CO(2) => W_reg_39_7_i_1_n_1,
   CO(3) => W_reg_39_7_i_1_n_0,
   O(0) => x71_out_4,
   O(1) => x71_out_5,
   O(2) => x71_out_6,
   O(3) => x71_out_7
);
W_reg_39_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x71_out_8,
   R => '0',
   Q => W_reg_39_8
);
W_reg_39_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x71_out_9,
   R => '0',
   Q => W_reg_39_9
);
W_reg_3_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_3_0,
   R => '0',
   Q => W_reg_3_0
);
W_reg_3_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_3_10,
   R => '0',
   Q => W_reg_3_10
);
W_reg_3_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_3_11,
   R => '0',
   Q => W_reg_3_11
);
W_reg_3_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_3_12,
   R => '0',
   Q => W_reg_3_12
);
W_reg_3_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_3_13,
   R => '0',
   Q => W_reg_3_13
);
W_reg_3_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_3_14,
   R => '0',
   Q => W_reg_3_14
);
W_reg_3_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_3_15,
   R => '0',
   Q => W_reg_3_15
);
W_reg_3_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_3_16,
   R => '0',
   Q => W_reg_3_16
);
W_reg_3_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_3_17,
   R => '0',
   Q => W_reg_3_17
);
W_reg_3_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_3_18,
   R => '0',
   Q => W_reg_3_18
);
W_reg_3_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_3_19,
   R => '0',
   Q => W_reg_3_19
);
W_reg_3_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_3_1,
   R => '0',
   Q => W_reg_3_1
);
W_reg_3_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_3_20,
   R => '0',
   Q => W_reg_3_20
);
W_reg_3_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_3_21,
   R => '0',
   Q => W_reg_3_21
);
W_reg_3_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_3_22,
   R => '0',
   Q => W_reg_3_22
);
W_reg_3_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_3_23,
   R => '0',
   Q => W_reg_3_23
);
W_reg_3_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_3_24,
   R => '0',
   Q => W_reg_3_24
);
W_reg_3_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_3_25,
   R => '0',
   Q => W_reg_3_25
);
W_reg_3_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_3_26,
   R => '0',
   Q => W_reg_3_26
);
W_reg_3_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_3_27,
   R => '0',
   Q => W_reg_3_27
);
W_reg_3_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_3_28,
   R => '0',
   Q => W_reg_3_28
);
W_reg_3_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_3_29,
   R => '0',
   Q => W_reg_3_29
);
W_reg_3_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_3_2,
   R => '0',
   Q => W_reg_3_2
);
W_reg_3_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_3_30,
   R => '0',
   Q => W_reg_3_30
);
W_reg_3_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_3_31,
   R => '0',
   Q => W_reg_3_31
);
W_reg_3_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_3_3,
   R => '0',
   Q => W_reg_3_3
);
W_reg_3_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_3_4,
   R => '0',
   Q => W_reg_3_4
);
W_reg_3_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_3_5,
   R => '0',
   Q => W_reg_3_5
);
W_reg_3_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_3_6,
   R => '0',
   Q => W_reg_3_6
);
W_reg_3_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_3_7,
   R => '0',
   Q => W_reg_3_7
);
W_reg_3_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_3_8,
   R => '0',
   Q => W_reg_3_8
);
W_reg_3_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_3_9,
   R => '0',
   Q => W_reg_3_9
);
W_reg_40_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x68_out_0,
   R => '0',
   Q => W_reg_40_0
);
W_reg_40_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x68_out_10,
   R => '0',
   Q => W_reg_40_10
);
W_reg_40_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x68_out_11,
   R => '0',
   Q => W_reg_40_11
);
W_reg_40_11_i_1 : CARRY4
 port map (
   CI => W_reg_40_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_40_11_i_5_n_0,
   DI(1) => W_40_11_i_4_n_0,
   DI(2) => W_40_11_i_3_n_0,
   DI(3) => W_40_11_i_2_n_0,
   S(0) => W_40_11_i_9_n_0,
   S(1) => W_40_11_i_8_n_0,
   S(2) => W_40_11_i_7_n_0,
   S(3) => W_40_11_i_6_n_0,
   CO(0) => W_reg_40_11_i_1_n_3,
   CO(1) => W_reg_40_11_i_1_n_2,
   CO(2) => W_reg_40_11_i_1_n_1,
   CO(3) => W_reg_40_11_i_1_n_0,
   O(0) => x68_out_8,
   O(1) => x68_out_9,
   O(2) => x68_out_10,
   O(3) => x68_out_11
);
W_reg_40_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x68_out_12,
   R => '0',
   Q => W_reg_40_12
);
W_reg_40_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x68_out_13,
   R => '0',
   Q => W_reg_40_13
);
W_reg_40_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x68_out_14,
   R => '0',
   Q => W_reg_40_14
);
W_reg_40_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x68_out_15,
   R => '0',
   Q => W_reg_40_15
);
W_reg_40_15_i_1 : CARRY4
 port map (
   CI => W_reg_40_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_40_15_i_5_n_0,
   DI(1) => W_40_15_i_4_n_0,
   DI(2) => W_40_15_i_3_n_0,
   DI(3) => W_40_15_i_2_n_0,
   S(0) => W_40_15_i_9_n_0,
   S(1) => W_40_15_i_8_n_0,
   S(2) => W_40_15_i_7_n_0,
   S(3) => W_40_15_i_6_n_0,
   CO(0) => W_reg_40_15_i_1_n_3,
   CO(1) => W_reg_40_15_i_1_n_2,
   CO(2) => W_reg_40_15_i_1_n_1,
   CO(3) => W_reg_40_15_i_1_n_0,
   O(0) => x68_out_12,
   O(1) => x68_out_13,
   O(2) => x68_out_14,
   O(3) => x68_out_15
);
W_reg_40_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x68_out_16,
   R => '0',
   Q => W_reg_40_16
);
W_reg_40_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x68_out_17,
   R => '0',
   Q => W_reg_40_17
);
W_reg_40_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x68_out_18,
   R => '0',
   Q => W_reg_40_18
);
W_reg_40_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x68_out_19,
   R => '0',
   Q => W_reg_40_19
);
W_reg_40_19_i_1 : CARRY4
 port map (
   CI => W_reg_40_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_40_19_i_5_n_0,
   DI(1) => W_40_19_i_4_n_0,
   DI(2) => W_40_19_i_3_n_0,
   DI(3) => W_40_19_i_2_n_0,
   S(0) => W_40_19_i_9_n_0,
   S(1) => W_40_19_i_8_n_0,
   S(2) => W_40_19_i_7_n_0,
   S(3) => W_40_19_i_6_n_0,
   CO(0) => W_reg_40_19_i_1_n_3,
   CO(1) => W_reg_40_19_i_1_n_2,
   CO(2) => W_reg_40_19_i_1_n_1,
   CO(3) => W_reg_40_19_i_1_n_0,
   O(0) => x68_out_16,
   O(1) => x68_out_17,
   O(2) => x68_out_18,
   O(3) => x68_out_19
);
W_reg_40_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x68_out_1,
   R => '0',
   Q => W_reg_40_1
);
W_reg_40_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x68_out_20,
   R => '0',
   Q => W_reg_40_20
);
W_reg_40_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x68_out_21,
   R => '0',
   Q => W_reg_40_21
);
W_reg_40_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x68_out_22,
   R => '0',
   Q => W_reg_40_22
);
W_reg_40_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x68_out_23,
   R => '0',
   Q => W_reg_40_23
);
W_reg_40_23_i_1 : CARRY4
 port map (
   CI => W_reg_40_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_40_23_i_5_n_0,
   DI(1) => W_40_23_i_4_n_0,
   DI(2) => W_40_23_i_3_n_0,
   DI(3) => W_40_23_i_2_n_0,
   S(0) => W_40_23_i_9_n_0,
   S(1) => W_40_23_i_8_n_0,
   S(2) => W_40_23_i_7_n_0,
   S(3) => W_40_23_i_6_n_0,
   CO(0) => W_reg_40_23_i_1_n_3,
   CO(1) => W_reg_40_23_i_1_n_2,
   CO(2) => W_reg_40_23_i_1_n_1,
   CO(3) => W_reg_40_23_i_1_n_0,
   O(0) => x68_out_20,
   O(1) => x68_out_21,
   O(2) => x68_out_22,
   O(3) => x68_out_23
);
W_reg_40_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x68_out_24,
   R => '0',
   Q => W_reg_40_24
);
W_reg_40_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x68_out_25,
   R => '0',
   Q => W_reg_40_25
);
W_reg_40_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x68_out_26,
   R => '0',
   Q => W_reg_40_26
);
W_reg_40_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x68_out_27,
   R => '0',
   Q => W_reg_40_27
);
W_reg_40_27_i_1 : CARRY4
 port map (
   CI => W_reg_40_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_40_27_i_5_n_0,
   DI(1) => W_40_27_i_4_n_0,
   DI(2) => W_40_27_i_3_n_0,
   DI(3) => W_40_27_i_2_n_0,
   S(0) => W_40_27_i_9_n_0,
   S(1) => W_40_27_i_8_n_0,
   S(2) => W_40_27_i_7_n_0,
   S(3) => W_40_27_i_6_n_0,
   CO(0) => W_reg_40_27_i_1_n_3,
   CO(1) => W_reg_40_27_i_1_n_2,
   CO(2) => W_reg_40_27_i_1_n_1,
   CO(3) => W_reg_40_27_i_1_n_0,
   O(0) => x68_out_24,
   O(1) => x68_out_25,
   O(2) => x68_out_26,
   O(3) => x68_out_27
);
W_reg_40_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x68_out_28,
   R => '0',
   Q => W_reg_40_28
);
W_reg_40_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x68_out_29,
   R => '0',
   Q => W_reg_40_29
);
W_reg_40_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x68_out_2,
   R => '0',
   Q => W_reg_40_2
);
W_reg_40_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x68_out_30,
   R => '0',
   Q => W_reg_40_30
);
W_reg_40_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x68_out_31,
   R => '0',
   Q => W_reg_40_31
);
W_reg_40_31_i_1 : CARRY4
 port map (
   CI => W_reg_40_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_40_31_i_4_n_0,
   DI(1) => W_40_31_i_3_n_0,
   DI(2) => W_40_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_40_31_i_8_n_0,
   S(1) => W_40_31_i_7_n_0,
   S(2) => W_40_31_i_6_n_0,
   S(3) => W_40_31_i_5_n_0,
   CO(0) => W_reg_40_31_i_1_n_3,
   CO(1) => W_reg_40_31_i_1_n_2,
   CO(2) => W_reg_40_31_i_1_n_1,
   CO(3) => NLW_W_reg_40_31_i_1_CO_UNCONNECTED_3,
   O(0) => x68_out_28,
   O(1) => x68_out_29,
   O(2) => x68_out_30,
   O(3) => x68_out_31
);
W_reg_40_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x68_out_3,
   R => '0',
   Q => W_reg_40_3
);
W_reg_40_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_40_3_i_5_n_0,
   DI(1) => W_40_3_i_4_n_0,
   DI(2) => W_40_3_i_3_n_0,
   DI(3) => W_40_3_i_2_n_0,
   S(0) => W_40_3_i_9_n_0,
   S(1) => W_40_3_i_8_n_0,
   S(2) => W_40_3_i_7_n_0,
   S(3) => W_40_3_i_6_n_0,
   CO(0) => W_reg_40_3_i_1_n_3,
   CO(1) => W_reg_40_3_i_1_n_2,
   CO(2) => W_reg_40_3_i_1_n_1,
   CO(3) => W_reg_40_3_i_1_n_0,
   O(0) => x68_out_0,
   O(1) => x68_out_1,
   O(2) => x68_out_2,
   O(3) => x68_out_3
);
W_reg_40_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x68_out_4,
   R => '0',
   Q => W_reg_40_4
);
W_reg_40_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x68_out_5,
   R => '0',
   Q => W_reg_40_5
);
W_reg_40_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x68_out_6,
   R => '0',
   Q => W_reg_40_6
);
W_reg_40_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x68_out_7,
   R => '0',
   Q => W_reg_40_7
);
W_reg_40_7_i_1 : CARRY4
 port map (
   CI => W_reg_40_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_40_7_i_5_n_0,
   DI(1) => W_40_7_i_4_n_0,
   DI(2) => W_40_7_i_3_n_0,
   DI(3) => W_40_7_i_2_n_0,
   S(0) => W_40_7_i_9_n_0,
   S(1) => W_40_7_i_8_n_0,
   S(2) => W_40_7_i_7_n_0,
   S(3) => W_40_7_i_6_n_0,
   CO(0) => W_reg_40_7_i_1_n_3,
   CO(1) => W_reg_40_7_i_1_n_2,
   CO(2) => W_reg_40_7_i_1_n_1,
   CO(3) => W_reg_40_7_i_1_n_0,
   O(0) => x68_out_4,
   O(1) => x68_out_5,
   O(2) => x68_out_6,
   O(3) => x68_out_7
);
W_reg_40_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x68_out_8,
   R => '0',
   Q => W_reg_40_8
);
W_reg_40_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x68_out_9,
   R => '0',
   Q => W_reg_40_9
);
W_reg_41_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x65_out_0,
   R => '0',
   Q => W_reg_41_0
);
W_reg_41_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x65_out_10,
   R => '0',
   Q => W_reg_41_10
);
W_reg_41_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x65_out_11,
   R => '0',
   Q => W_reg_41_11
);
W_reg_41_11_i_1 : CARRY4
 port map (
   CI => W_reg_41_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_41_11_i_5_n_0,
   DI(1) => W_41_11_i_4_n_0,
   DI(2) => W_41_11_i_3_n_0,
   DI(3) => W_41_11_i_2_n_0,
   S(0) => W_41_11_i_9_n_0,
   S(1) => W_41_11_i_8_n_0,
   S(2) => W_41_11_i_7_n_0,
   S(3) => W_41_11_i_6_n_0,
   CO(0) => W_reg_41_11_i_1_n_3,
   CO(1) => W_reg_41_11_i_1_n_2,
   CO(2) => W_reg_41_11_i_1_n_1,
   CO(3) => W_reg_41_11_i_1_n_0,
   O(0) => x65_out_8,
   O(1) => x65_out_9,
   O(2) => x65_out_10,
   O(3) => x65_out_11
);
W_reg_41_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x65_out_12,
   R => '0',
   Q => W_reg_41_12
);
W_reg_41_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x65_out_13,
   R => '0',
   Q => W_reg_41_13
);
W_reg_41_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x65_out_14,
   R => '0',
   Q => W_reg_41_14
);
W_reg_41_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x65_out_15,
   R => '0',
   Q => W_reg_41_15
);
W_reg_41_15_i_1 : CARRY4
 port map (
   CI => W_reg_41_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_41_15_i_5_n_0,
   DI(1) => W_41_15_i_4_n_0,
   DI(2) => W_41_15_i_3_n_0,
   DI(3) => W_41_15_i_2_n_0,
   S(0) => W_41_15_i_9_n_0,
   S(1) => W_41_15_i_8_n_0,
   S(2) => W_41_15_i_7_n_0,
   S(3) => W_41_15_i_6_n_0,
   CO(0) => W_reg_41_15_i_1_n_3,
   CO(1) => W_reg_41_15_i_1_n_2,
   CO(2) => W_reg_41_15_i_1_n_1,
   CO(3) => W_reg_41_15_i_1_n_0,
   O(0) => x65_out_12,
   O(1) => x65_out_13,
   O(2) => x65_out_14,
   O(3) => x65_out_15
);
W_reg_41_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x65_out_16,
   R => '0',
   Q => W_reg_41_16
);
W_reg_41_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x65_out_17,
   R => '0',
   Q => W_reg_41_17
);
W_reg_41_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x65_out_18,
   R => '0',
   Q => W_reg_41_18
);
W_reg_41_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x65_out_19,
   R => '0',
   Q => W_reg_41_19
);
W_reg_41_19_i_1 : CARRY4
 port map (
   CI => W_reg_41_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_41_19_i_5_n_0,
   DI(1) => W_41_19_i_4_n_0,
   DI(2) => W_41_19_i_3_n_0,
   DI(3) => W_41_19_i_2_n_0,
   S(0) => W_41_19_i_9_n_0,
   S(1) => W_41_19_i_8_n_0,
   S(2) => W_41_19_i_7_n_0,
   S(3) => W_41_19_i_6_n_0,
   CO(0) => W_reg_41_19_i_1_n_3,
   CO(1) => W_reg_41_19_i_1_n_2,
   CO(2) => W_reg_41_19_i_1_n_1,
   CO(3) => W_reg_41_19_i_1_n_0,
   O(0) => x65_out_16,
   O(1) => x65_out_17,
   O(2) => x65_out_18,
   O(3) => x65_out_19
);
W_reg_41_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x65_out_1,
   R => '0',
   Q => W_reg_41_1
);
W_reg_41_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x65_out_20,
   R => '0',
   Q => W_reg_41_20
);
W_reg_41_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x65_out_21,
   R => '0',
   Q => W_reg_41_21
);
W_reg_41_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x65_out_22,
   R => '0',
   Q => W_reg_41_22
);
W_reg_41_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x65_out_23,
   R => '0',
   Q => W_reg_41_23
);
W_reg_41_23_i_1 : CARRY4
 port map (
   CI => W_reg_41_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_41_23_i_5_n_0,
   DI(1) => W_41_23_i_4_n_0,
   DI(2) => W_41_23_i_3_n_0,
   DI(3) => W_41_23_i_2_n_0,
   S(0) => W_41_23_i_9_n_0,
   S(1) => W_41_23_i_8_n_0,
   S(2) => W_41_23_i_7_n_0,
   S(3) => W_41_23_i_6_n_0,
   CO(0) => W_reg_41_23_i_1_n_3,
   CO(1) => W_reg_41_23_i_1_n_2,
   CO(2) => W_reg_41_23_i_1_n_1,
   CO(3) => W_reg_41_23_i_1_n_0,
   O(0) => x65_out_20,
   O(1) => x65_out_21,
   O(2) => x65_out_22,
   O(3) => x65_out_23
);
W_reg_41_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x65_out_24,
   R => '0',
   Q => W_reg_41_24
);
W_reg_41_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x65_out_25,
   R => '0',
   Q => W_reg_41_25
);
W_reg_41_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x65_out_26,
   R => '0',
   Q => W_reg_41_26
);
W_reg_41_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x65_out_27,
   R => '0',
   Q => W_reg_41_27
);
W_reg_41_27_i_1 : CARRY4
 port map (
   CI => W_reg_41_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_41_27_i_5_n_0,
   DI(1) => W_41_27_i_4_n_0,
   DI(2) => W_41_27_i_3_n_0,
   DI(3) => W_41_27_i_2_n_0,
   S(0) => W_41_27_i_9_n_0,
   S(1) => W_41_27_i_8_n_0,
   S(2) => W_41_27_i_7_n_0,
   S(3) => W_41_27_i_6_n_0,
   CO(0) => W_reg_41_27_i_1_n_3,
   CO(1) => W_reg_41_27_i_1_n_2,
   CO(2) => W_reg_41_27_i_1_n_1,
   CO(3) => W_reg_41_27_i_1_n_0,
   O(0) => x65_out_24,
   O(1) => x65_out_25,
   O(2) => x65_out_26,
   O(3) => x65_out_27
);
W_reg_41_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x65_out_28,
   R => '0',
   Q => W_reg_41_28
);
W_reg_41_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x65_out_29,
   R => '0',
   Q => W_reg_41_29
);
W_reg_41_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x65_out_2,
   R => '0',
   Q => W_reg_41_2
);
W_reg_41_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x65_out_30,
   R => '0',
   Q => W_reg_41_30
);
W_reg_41_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x65_out_31,
   R => '0',
   Q => W_reg_41_31
);
W_reg_41_31_i_1 : CARRY4
 port map (
   CI => W_reg_41_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_41_31_i_4_n_0,
   DI(1) => W_41_31_i_3_n_0,
   DI(2) => W_41_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_41_31_i_8_n_0,
   S(1) => W_41_31_i_7_n_0,
   S(2) => W_41_31_i_6_n_0,
   S(3) => W_41_31_i_5_n_0,
   CO(0) => W_reg_41_31_i_1_n_3,
   CO(1) => W_reg_41_31_i_1_n_2,
   CO(2) => W_reg_41_31_i_1_n_1,
   CO(3) => NLW_W_reg_41_31_i_1_CO_UNCONNECTED_3,
   O(0) => x65_out_28,
   O(1) => x65_out_29,
   O(2) => x65_out_30,
   O(3) => x65_out_31
);
W_reg_41_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x65_out_3,
   R => '0',
   Q => W_reg_41_3
);
W_reg_41_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_41_3_i_5_n_0,
   DI(1) => W_41_3_i_4_n_0,
   DI(2) => W_41_3_i_3_n_0,
   DI(3) => W_41_3_i_2_n_0,
   S(0) => W_41_3_i_9_n_0,
   S(1) => W_41_3_i_8_n_0,
   S(2) => W_41_3_i_7_n_0,
   S(3) => W_41_3_i_6_n_0,
   CO(0) => W_reg_41_3_i_1_n_3,
   CO(1) => W_reg_41_3_i_1_n_2,
   CO(2) => W_reg_41_3_i_1_n_1,
   CO(3) => W_reg_41_3_i_1_n_0,
   O(0) => x65_out_0,
   O(1) => x65_out_1,
   O(2) => x65_out_2,
   O(3) => x65_out_3
);
W_reg_41_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x65_out_4,
   R => '0',
   Q => W_reg_41_4
);
W_reg_41_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x65_out_5,
   R => '0',
   Q => W_reg_41_5
);
W_reg_41_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x65_out_6,
   R => '0',
   Q => W_reg_41_6
);
W_reg_41_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x65_out_7,
   R => '0',
   Q => W_reg_41_7
);
W_reg_41_7_i_1 : CARRY4
 port map (
   CI => W_reg_41_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_41_7_i_5_n_0,
   DI(1) => W_41_7_i_4_n_0,
   DI(2) => W_41_7_i_3_n_0,
   DI(3) => W_41_7_i_2_n_0,
   S(0) => W_41_7_i_9_n_0,
   S(1) => W_41_7_i_8_n_0,
   S(2) => W_41_7_i_7_n_0,
   S(3) => W_41_7_i_6_n_0,
   CO(0) => W_reg_41_7_i_1_n_3,
   CO(1) => W_reg_41_7_i_1_n_2,
   CO(2) => W_reg_41_7_i_1_n_1,
   CO(3) => W_reg_41_7_i_1_n_0,
   O(0) => x65_out_4,
   O(1) => x65_out_5,
   O(2) => x65_out_6,
   O(3) => x65_out_7
);
W_reg_41_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x65_out_8,
   R => '0',
   Q => W_reg_41_8
);
W_reg_41_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x65_out_9,
   R => '0',
   Q => W_reg_41_9
);
W_reg_42_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x62_out_0,
   R => '0',
   Q => W_reg_42_0
);
W_reg_42_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x62_out_10,
   R => '0',
   Q => W_reg_42_10
);
W_reg_42_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x62_out_11,
   R => '0',
   Q => W_reg_42_11
);
W_reg_42_11_i_1 : CARRY4
 port map (
   CI => W_reg_42_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_42_11_i_5_n_0,
   DI(1) => W_42_11_i_4_n_0,
   DI(2) => W_42_11_i_3_n_0,
   DI(3) => W_42_11_i_2_n_0,
   S(0) => W_42_11_i_9_n_0,
   S(1) => W_42_11_i_8_n_0,
   S(2) => W_42_11_i_7_n_0,
   S(3) => W_42_11_i_6_n_0,
   CO(0) => W_reg_42_11_i_1_n_3,
   CO(1) => W_reg_42_11_i_1_n_2,
   CO(2) => W_reg_42_11_i_1_n_1,
   CO(3) => W_reg_42_11_i_1_n_0,
   O(0) => x62_out_8,
   O(1) => x62_out_9,
   O(2) => x62_out_10,
   O(3) => x62_out_11
);
W_reg_42_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x62_out_12,
   R => '0',
   Q => W_reg_42_12
);
W_reg_42_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x62_out_13,
   R => '0',
   Q => W_reg_42_13
);
W_reg_42_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x62_out_14,
   R => '0',
   Q => W_reg_42_14
);
W_reg_42_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x62_out_15,
   R => '0',
   Q => W_reg_42_15
);
W_reg_42_15_i_1 : CARRY4
 port map (
   CI => W_reg_42_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_42_15_i_5_n_0,
   DI(1) => W_42_15_i_4_n_0,
   DI(2) => W_42_15_i_3_n_0,
   DI(3) => W_42_15_i_2_n_0,
   S(0) => W_42_15_i_9_n_0,
   S(1) => W_42_15_i_8_n_0,
   S(2) => W_42_15_i_7_n_0,
   S(3) => W_42_15_i_6_n_0,
   CO(0) => W_reg_42_15_i_1_n_3,
   CO(1) => W_reg_42_15_i_1_n_2,
   CO(2) => W_reg_42_15_i_1_n_1,
   CO(3) => W_reg_42_15_i_1_n_0,
   O(0) => x62_out_12,
   O(1) => x62_out_13,
   O(2) => x62_out_14,
   O(3) => x62_out_15
);
W_reg_42_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x62_out_16,
   R => '0',
   Q => W_reg_42_16
);
W_reg_42_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x62_out_17,
   R => '0',
   Q => W_reg_42_17
);
W_reg_42_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x62_out_18,
   R => '0',
   Q => W_reg_42_18
);
W_reg_42_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x62_out_19,
   R => '0',
   Q => W_reg_42_19
);
W_reg_42_19_i_1 : CARRY4
 port map (
   CI => W_reg_42_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_42_19_i_5_n_0,
   DI(1) => W_42_19_i_4_n_0,
   DI(2) => W_42_19_i_3_n_0,
   DI(3) => W_42_19_i_2_n_0,
   S(0) => W_42_19_i_9_n_0,
   S(1) => W_42_19_i_8_n_0,
   S(2) => W_42_19_i_7_n_0,
   S(3) => W_42_19_i_6_n_0,
   CO(0) => W_reg_42_19_i_1_n_3,
   CO(1) => W_reg_42_19_i_1_n_2,
   CO(2) => W_reg_42_19_i_1_n_1,
   CO(3) => W_reg_42_19_i_1_n_0,
   O(0) => x62_out_16,
   O(1) => x62_out_17,
   O(2) => x62_out_18,
   O(3) => x62_out_19
);
W_reg_42_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x62_out_1,
   R => '0',
   Q => W_reg_42_1
);
W_reg_42_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x62_out_20,
   R => '0',
   Q => W_reg_42_20
);
W_reg_42_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x62_out_21,
   R => '0',
   Q => W_reg_42_21
);
W_reg_42_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x62_out_22,
   R => '0',
   Q => W_reg_42_22
);
W_reg_42_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x62_out_23,
   R => '0',
   Q => W_reg_42_23
);
W_reg_42_23_i_1 : CARRY4
 port map (
   CI => W_reg_42_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_42_23_i_5_n_0,
   DI(1) => W_42_23_i_4_n_0,
   DI(2) => W_42_23_i_3_n_0,
   DI(3) => W_42_23_i_2_n_0,
   S(0) => W_42_23_i_9_n_0,
   S(1) => W_42_23_i_8_n_0,
   S(2) => W_42_23_i_7_n_0,
   S(3) => W_42_23_i_6_n_0,
   CO(0) => W_reg_42_23_i_1_n_3,
   CO(1) => W_reg_42_23_i_1_n_2,
   CO(2) => W_reg_42_23_i_1_n_1,
   CO(3) => W_reg_42_23_i_1_n_0,
   O(0) => x62_out_20,
   O(1) => x62_out_21,
   O(2) => x62_out_22,
   O(3) => x62_out_23
);
W_reg_42_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x62_out_24,
   R => '0',
   Q => W_reg_42_24
);
W_reg_42_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x62_out_25,
   R => '0',
   Q => W_reg_42_25
);
W_reg_42_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x62_out_26,
   R => '0',
   Q => W_reg_42_26
);
W_reg_42_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x62_out_27,
   R => '0',
   Q => W_reg_42_27
);
W_reg_42_27_i_1 : CARRY4
 port map (
   CI => W_reg_42_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_42_27_i_5_n_0,
   DI(1) => W_42_27_i_4_n_0,
   DI(2) => W_42_27_i_3_n_0,
   DI(3) => W_42_27_i_2_n_0,
   S(0) => W_42_27_i_9_n_0,
   S(1) => W_42_27_i_8_n_0,
   S(2) => W_42_27_i_7_n_0,
   S(3) => W_42_27_i_6_n_0,
   CO(0) => W_reg_42_27_i_1_n_3,
   CO(1) => W_reg_42_27_i_1_n_2,
   CO(2) => W_reg_42_27_i_1_n_1,
   CO(3) => W_reg_42_27_i_1_n_0,
   O(0) => x62_out_24,
   O(1) => x62_out_25,
   O(2) => x62_out_26,
   O(3) => x62_out_27
);
W_reg_42_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x62_out_28,
   R => '0',
   Q => W_reg_42_28
);
W_reg_42_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x62_out_29,
   R => '0',
   Q => W_reg_42_29
);
W_reg_42_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x62_out_2,
   R => '0',
   Q => W_reg_42_2
);
W_reg_42_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x62_out_30,
   R => '0',
   Q => W_reg_42_30
);
W_reg_42_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x62_out_31,
   R => '0',
   Q => W_reg_42_31
);
W_reg_42_31_i_1 : CARRY4
 port map (
   CI => W_reg_42_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_42_31_i_4_n_0,
   DI(1) => W_42_31_i_3_n_0,
   DI(2) => W_42_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_42_31_i_8_n_0,
   S(1) => W_42_31_i_7_n_0,
   S(2) => W_42_31_i_6_n_0,
   S(3) => W_42_31_i_5_n_0,
   CO(0) => W_reg_42_31_i_1_n_3,
   CO(1) => W_reg_42_31_i_1_n_2,
   CO(2) => W_reg_42_31_i_1_n_1,
   CO(3) => NLW_W_reg_42_31_i_1_CO_UNCONNECTED_3,
   O(0) => x62_out_28,
   O(1) => x62_out_29,
   O(2) => x62_out_30,
   O(3) => x62_out_31
);
W_reg_42_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x62_out_3,
   R => '0',
   Q => W_reg_42_3
);
W_reg_42_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_42_3_i_5_n_0,
   DI(1) => W_42_3_i_4_n_0,
   DI(2) => W_42_3_i_3_n_0,
   DI(3) => W_42_3_i_2_n_0,
   S(0) => W_42_3_i_9_n_0,
   S(1) => W_42_3_i_8_n_0,
   S(2) => W_42_3_i_7_n_0,
   S(3) => W_42_3_i_6_n_0,
   CO(0) => W_reg_42_3_i_1_n_3,
   CO(1) => W_reg_42_3_i_1_n_2,
   CO(2) => W_reg_42_3_i_1_n_1,
   CO(3) => W_reg_42_3_i_1_n_0,
   O(0) => x62_out_0,
   O(1) => x62_out_1,
   O(2) => x62_out_2,
   O(3) => x62_out_3
);
W_reg_42_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x62_out_4,
   R => '0',
   Q => W_reg_42_4
);
W_reg_42_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x62_out_5,
   R => '0',
   Q => W_reg_42_5
);
W_reg_42_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x62_out_6,
   R => '0',
   Q => W_reg_42_6
);
W_reg_42_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x62_out_7,
   R => '0',
   Q => W_reg_42_7
);
W_reg_42_7_i_1 : CARRY4
 port map (
   CI => W_reg_42_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_42_7_i_5_n_0,
   DI(1) => W_42_7_i_4_n_0,
   DI(2) => W_42_7_i_3_n_0,
   DI(3) => W_42_7_i_2_n_0,
   S(0) => W_42_7_i_9_n_0,
   S(1) => W_42_7_i_8_n_0,
   S(2) => W_42_7_i_7_n_0,
   S(3) => W_42_7_i_6_n_0,
   CO(0) => W_reg_42_7_i_1_n_3,
   CO(1) => W_reg_42_7_i_1_n_2,
   CO(2) => W_reg_42_7_i_1_n_1,
   CO(3) => W_reg_42_7_i_1_n_0,
   O(0) => x62_out_4,
   O(1) => x62_out_5,
   O(2) => x62_out_6,
   O(3) => x62_out_7
);
W_reg_42_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x62_out_8,
   R => '0',
   Q => W_reg_42_8
);
W_reg_42_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x62_out_9,
   R => '0',
   Q => W_reg_42_9
);
W_reg_43_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x59_out_0,
   R => '0',
   Q => W_reg_43_0
);
W_reg_43_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x59_out_10,
   R => '0',
   Q => W_reg_43_10
);
W_reg_43_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x59_out_11,
   R => '0',
   Q => W_reg_43_11
);
W_reg_43_11_i_1 : CARRY4
 port map (
   CI => W_reg_43_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_43_11_i_5_n_0,
   DI(1) => W_43_11_i_4_n_0,
   DI(2) => W_43_11_i_3_n_0,
   DI(3) => W_43_11_i_2_n_0,
   S(0) => W_43_11_i_9_n_0,
   S(1) => W_43_11_i_8_n_0,
   S(2) => W_43_11_i_7_n_0,
   S(3) => W_43_11_i_6_n_0,
   CO(0) => W_reg_43_11_i_1_n_3,
   CO(1) => W_reg_43_11_i_1_n_2,
   CO(2) => W_reg_43_11_i_1_n_1,
   CO(3) => W_reg_43_11_i_1_n_0,
   O(0) => x59_out_8,
   O(1) => x59_out_9,
   O(2) => x59_out_10,
   O(3) => x59_out_11
);
W_reg_43_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x59_out_12,
   R => '0',
   Q => W_reg_43_12
);
W_reg_43_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x59_out_13,
   R => '0',
   Q => W_reg_43_13
);
W_reg_43_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x59_out_14,
   R => '0',
   Q => W_reg_43_14
);
W_reg_43_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x59_out_15,
   R => '0',
   Q => W_reg_43_15
);
W_reg_43_15_i_1 : CARRY4
 port map (
   CI => W_reg_43_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_43_15_i_5_n_0,
   DI(1) => W_43_15_i_4_n_0,
   DI(2) => W_43_15_i_3_n_0,
   DI(3) => W_43_15_i_2_n_0,
   S(0) => W_43_15_i_9_n_0,
   S(1) => W_43_15_i_8_n_0,
   S(2) => W_43_15_i_7_n_0,
   S(3) => W_43_15_i_6_n_0,
   CO(0) => W_reg_43_15_i_1_n_3,
   CO(1) => W_reg_43_15_i_1_n_2,
   CO(2) => W_reg_43_15_i_1_n_1,
   CO(3) => W_reg_43_15_i_1_n_0,
   O(0) => x59_out_12,
   O(1) => x59_out_13,
   O(2) => x59_out_14,
   O(3) => x59_out_15
);
W_reg_43_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x59_out_16,
   R => '0',
   Q => W_reg_43_16
);
W_reg_43_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x59_out_17,
   R => '0',
   Q => W_reg_43_17
);
W_reg_43_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x59_out_18,
   R => '0',
   Q => W_reg_43_18
);
W_reg_43_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x59_out_19,
   R => '0',
   Q => W_reg_43_19
);
W_reg_43_19_i_1 : CARRY4
 port map (
   CI => W_reg_43_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_43_19_i_5_n_0,
   DI(1) => W_43_19_i_4_n_0,
   DI(2) => W_43_19_i_3_n_0,
   DI(3) => W_43_19_i_2_n_0,
   S(0) => W_43_19_i_9_n_0,
   S(1) => W_43_19_i_8_n_0,
   S(2) => W_43_19_i_7_n_0,
   S(3) => W_43_19_i_6_n_0,
   CO(0) => W_reg_43_19_i_1_n_3,
   CO(1) => W_reg_43_19_i_1_n_2,
   CO(2) => W_reg_43_19_i_1_n_1,
   CO(3) => W_reg_43_19_i_1_n_0,
   O(0) => x59_out_16,
   O(1) => x59_out_17,
   O(2) => x59_out_18,
   O(3) => x59_out_19
);
W_reg_43_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x59_out_1,
   R => '0',
   Q => W_reg_43_1
);
W_reg_43_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x59_out_20,
   R => '0',
   Q => W_reg_43_20
);
W_reg_43_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x59_out_21,
   R => '0',
   Q => W_reg_43_21
);
W_reg_43_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x59_out_22,
   R => '0',
   Q => W_reg_43_22
);
W_reg_43_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x59_out_23,
   R => '0',
   Q => W_reg_43_23
);
W_reg_43_23_i_1 : CARRY4
 port map (
   CI => W_reg_43_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_43_23_i_5_n_0,
   DI(1) => W_43_23_i_4_n_0,
   DI(2) => W_43_23_i_3_n_0,
   DI(3) => W_43_23_i_2_n_0,
   S(0) => W_43_23_i_9_n_0,
   S(1) => W_43_23_i_8_n_0,
   S(2) => W_43_23_i_7_n_0,
   S(3) => W_43_23_i_6_n_0,
   CO(0) => W_reg_43_23_i_1_n_3,
   CO(1) => W_reg_43_23_i_1_n_2,
   CO(2) => W_reg_43_23_i_1_n_1,
   CO(3) => W_reg_43_23_i_1_n_0,
   O(0) => x59_out_20,
   O(1) => x59_out_21,
   O(2) => x59_out_22,
   O(3) => x59_out_23
);
W_reg_43_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x59_out_24,
   R => '0',
   Q => W_reg_43_24
);
W_reg_43_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x59_out_25,
   R => '0',
   Q => W_reg_43_25
);
W_reg_43_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x59_out_26,
   R => '0',
   Q => W_reg_43_26
);
W_reg_43_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x59_out_27,
   R => '0',
   Q => W_reg_43_27
);
W_reg_43_27_i_1 : CARRY4
 port map (
   CI => W_reg_43_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_43_27_i_5_n_0,
   DI(1) => W_43_27_i_4_n_0,
   DI(2) => W_43_27_i_3_n_0,
   DI(3) => W_43_27_i_2_n_0,
   S(0) => W_43_27_i_9_n_0,
   S(1) => W_43_27_i_8_n_0,
   S(2) => W_43_27_i_7_n_0,
   S(3) => W_43_27_i_6_n_0,
   CO(0) => W_reg_43_27_i_1_n_3,
   CO(1) => W_reg_43_27_i_1_n_2,
   CO(2) => W_reg_43_27_i_1_n_1,
   CO(3) => W_reg_43_27_i_1_n_0,
   O(0) => x59_out_24,
   O(1) => x59_out_25,
   O(2) => x59_out_26,
   O(3) => x59_out_27
);
W_reg_43_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x59_out_28,
   R => '0',
   Q => W_reg_43_28
);
W_reg_43_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x59_out_29,
   R => '0',
   Q => W_reg_43_29
);
W_reg_43_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x59_out_2,
   R => '0',
   Q => W_reg_43_2
);
W_reg_43_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x59_out_30,
   R => '0',
   Q => W_reg_43_30
);
W_reg_43_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x59_out_31,
   R => '0',
   Q => W_reg_43_31
);
W_reg_43_31_i_1 : CARRY4
 port map (
   CI => W_reg_43_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_43_31_i_4_n_0,
   DI(1) => W_43_31_i_3_n_0,
   DI(2) => W_43_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_43_31_i_8_n_0,
   S(1) => W_43_31_i_7_n_0,
   S(2) => W_43_31_i_6_n_0,
   S(3) => W_43_31_i_5_n_0,
   CO(0) => W_reg_43_31_i_1_n_3,
   CO(1) => W_reg_43_31_i_1_n_2,
   CO(2) => W_reg_43_31_i_1_n_1,
   CO(3) => NLW_W_reg_43_31_i_1_CO_UNCONNECTED_3,
   O(0) => x59_out_28,
   O(1) => x59_out_29,
   O(2) => x59_out_30,
   O(3) => x59_out_31
);
W_reg_43_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x59_out_3,
   R => '0',
   Q => W_reg_43_3
);
W_reg_43_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_43_3_i_5_n_0,
   DI(1) => W_43_3_i_4_n_0,
   DI(2) => W_43_3_i_3_n_0,
   DI(3) => W_43_3_i_2_n_0,
   S(0) => W_43_3_i_9_n_0,
   S(1) => W_43_3_i_8_n_0,
   S(2) => W_43_3_i_7_n_0,
   S(3) => W_43_3_i_6_n_0,
   CO(0) => W_reg_43_3_i_1_n_3,
   CO(1) => W_reg_43_3_i_1_n_2,
   CO(2) => W_reg_43_3_i_1_n_1,
   CO(3) => W_reg_43_3_i_1_n_0,
   O(0) => x59_out_0,
   O(1) => x59_out_1,
   O(2) => x59_out_2,
   O(3) => x59_out_3
);
W_reg_43_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x59_out_4,
   R => '0',
   Q => W_reg_43_4
);
W_reg_43_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x59_out_5,
   R => '0',
   Q => W_reg_43_5
);
W_reg_43_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x59_out_6,
   R => '0',
   Q => W_reg_43_6
);
W_reg_43_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x59_out_7,
   R => '0',
   Q => W_reg_43_7
);
W_reg_43_7_i_1 : CARRY4
 port map (
   CI => W_reg_43_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_43_7_i_5_n_0,
   DI(1) => W_43_7_i_4_n_0,
   DI(2) => W_43_7_i_3_n_0,
   DI(3) => W_43_7_i_2_n_0,
   S(0) => W_43_7_i_9_n_0,
   S(1) => W_43_7_i_8_n_0,
   S(2) => W_43_7_i_7_n_0,
   S(3) => W_43_7_i_6_n_0,
   CO(0) => W_reg_43_7_i_1_n_3,
   CO(1) => W_reg_43_7_i_1_n_2,
   CO(2) => W_reg_43_7_i_1_n_1,
   CO(3) => W_reg_43_7_i_1_n_0,
   O(0) => x59_out_4,
   O(1) => x59_out_5,
   O(2) => x59_out_6,
   O(3) => x59_out_7
);
W_reg_43_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x59_out_8,
   R => '0',
   Q => W_reg_43_8
);
W_reg_43_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x59_out_9,
   R => '0',
   Q => W_reg_43_9
);
W_reg_44_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x56_out_0,
   R => '0',
   Q => W_reg_44_0
);
W_reg_44_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x56_out_10,
   R => '0',
   Q => W_reg_44_10
);
W_reg_44_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x56_out_11,
   R => '0',
   Q => W_reg_44_11
);
W_reg_44_11_i_1 : CARRY4
 port map (
   CI => W_reg_44_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_44_11_i_5_n_0,
   DI(1) => W_44_11_i_4_n_0,
   DI(2) => W_44_11_i_3_n_0,
   DI(3) => W_44_11_i_2_n_0,
   S(0) => W_44_11_i_9_n_0,
   S(1) => W_44_11_i_8_n_0,
   S(2) => W_44_11_i_7_n_0,
   S(3) => W_44_11_i_6_n_0,
   CO(0) => W_reg_44_11_i_1_n_3,
   CO(1) => W_reg_44_11_i_1_n_2,
   CO(2) => W_reg_44_11_i_1_n_1,
   CO(3) => W_reg_44_11_i_1_n_0,
   O(0) => x56_out_8,
   O(1) => x56_out_9,
   O(2) => x56_out_10,
   O(3) => x56_out_11
);
W_reg_44_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x56_out_12,
   R => '0',
   Q => W_reg_44_12
);
W_reg_44_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x56_out_13,
   R => '0',
   Q => W_reg_44_13
);
W_reg_44_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x56_out_14,
   R => '0',
   Q => W_reg_44_14
);
W_reg_44_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x56_out_15,
   R => '0',
   Q => W_reg_44_15
);
W_reg_44_15_i_1 : CARRY4
 port map (
   CI => W_reg_44_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_44_15_i_5_n_0,
   DI(1) => W_44_15_i_4_n_0,
   DI(2) => W_44_15_i_3_n_0,
   DI(3) => W_44_15_i_2_n_0,
   S(0) => W_44_15_i_9_n_0,
   S(1) => W_44_15_i_8_n_0,
   S(2) => W_44_15_i_7_n_0,
   S(3) => W_44_15_i_6_n_0,
   CO(0) => W_reg_44_15_i_1_n_3,
   CO(1) => W_reg_44_15_i_1_n_2,
   CO(2) => W_reg_44_15_i_1_n_1,
   CO(3) => W_reg_44_15_i_1_n_0,
   O(0) => x56_out_12,
   O(1) => x56_out_13,
   O(2) => x56_out_14,
   O(3) => x56_out_15
);
W_reg_44_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x56_out_16,
   R => '0',
   Q => W_reg_44_16
);
W_reg_44_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x56_out_17,
   R => '0',
   Q => W_reg_44_17
);
W_reg_44_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x56_out_18,
   R => '0',
   Q => W_reg_44_18
);
W_reg_44_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x56_out_19,
   R => '0',
   Q => W_reg_44_19
);
W_reg_44_19_i_1 : CARRY4
 port map (
   CI => W_reg_44_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_44_19_i_5_n_0,
   DI(1) => W_44_19_i_4_n_0,
   DI(2) => W_44_19_i_3_n_0,
   DI(3) => W_44_19_i_2_n_0,
   S(0) => W_44_19_i_9_n_0,
   S(1) => W_44_19_i_8_n_0,
   S(2) => W_44_19_i_7_n_0,
   S(3) => W_44_19_i_6_n_0,
   CO(0) => W_reg_44_19_i_1_n_3,
   CO(1) => W_reg_44_19_i_1_n_2,
   CO(2) => W_reg_44_19_i_1_n_1,
   CO(3) => W_reg_44_19_i_1_n_0,
   O(0) => x56_out_16,
   O(1) => x56_out_17,
   O(2) => x56_out_18,
   O(3) => x56_out_19
);
W_reg_44_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x56_out_1,
   R => '0',
   Q => W_reg_44_1
);
W_reg_44_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x56_out_20,
   R => '0',
   Q => W_reg_44_20
);
W_reg_44_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x56_out_21,
   R => '0',
   Q => W_reg_44_21
);
W_reg_44_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x56_out_22,
   R => '0',
   Q => W_reg_44_22
);
W_reg_44_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x56_out_23,
   R => '0',
   Q => W_reg_44_23
);
W_reg_44_23_i_1 : CARRY4
 port map (
   CI => W_reg_44_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_44_23_i_5_n_0,
   DI(1) => W_44_23_i_4_n_0,
   DI(2) => W_44_23_i_3_n_0,
   DI(3) => W_44_23_i_2_n_0,
   S(0) => W_44_23_i_9_n_0,
   S(1) => W_44_23_i_8_n_0,
   S(2) => W_44_23_i_7_n_0,
   S(3) => W_44_23_i_6_n_0,
   CO(0) => W_reg_44_23_i_1_n_3,
   CO(1) => W_reg_44_23_i_1_n_2,
   CO(2) => W_reg_44_23_i_1_n_1,
   CO(3) => W_reg_44_23_i_1_n_0,
   O(0) => x56_out_20,
   O(1) => x56_out_21,
   O(2) => x56_out_22,
   O(3) => x56_out_23
);
W_reg_44_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x56_out_24,
   R => '0',
   Q => W_reg_44_24
);
W_reg_44_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x56_out_25,
   R => '0',
   Q => W_reg_44_25
);
W_reg_44_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x56_out_26,
   R => '0',
   Q => W_reg_44_26
);
W_reg_44_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x56_out_27,
   R => '0',
   Q => W_reg_44_27
);
W_reg_44_27_i_1 : CARRY4
 port map (
   CI => W_reg_44_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_44_27_i_5_n_0,
   DI(1) => W_44_27_i_4_n_0,
   DI(2) => W_44_27_i_3_n_0,
   DI(3) => W_44_27_i_2_n_0,
   S(0) => W_44_27_i_9_n_0,
   S(1) => W_44_27_i_8_n_0,
   S(2) => W_44_27_i_7_n_0,
   S(3) => W_44_27_i_6_n_0,
   CO(0) => W_reg_44_27_i_1_n_3,
   CO(1) => W_reg_44_27_i_1_n_2,
   CO(2) => W_reg_44_27_i_1_n_1,
   CO(3) => W_reg_44_27_i_1_n_0,
   O(0) => x56_out_24,
   O(1) => x56_out_25,
   O(2) => x56_out_26,
   O(3) => x56_out_27
);
W_reg_44_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x56_out_28,
   R => '0',
   Q => W_reg_44_28
);
W_reg_44_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x56_out_29,
   R => '0',
   Q => W_reg_44_29
);
W_reg_44_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x56_out_2,
   R => '0',
   Q => W_reg_44_2
);
W_reg_44_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x56_out_30,
   R => '0',
   Q => W_reg_44_30
);
W_reg_44_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x56_out_31,
   R => '0',
   Q => W_reg_44_31
);
W_reg_44_31_i_1 : CARRY4
 port map (
   CI => W_reg_44_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_44_31_i_4_n_0,
   DI(1) => W_44_31_i_3_n_0,
   DI(2) => W_44_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_44_31_i_8_n_0,
   S(1) => W_44_31_i_7_n_0,
   S(2) => W_44_31_i_6_n_0,
   S(3) => W_44_31_i_5_n_0,
   CO(0) => W_reg_44_31_i_1_n_3,
   CO(1) => W_reg_44_31_i_1_n_2,
   CO(2) => W_reg_44_31_i_1_n_1,
   CO(3) => NLW_W_reg_44_31_i_1_CO_UNCONNECTED_3,
   O(0) => x56_out_28,
   O(1) => x56_out_29,
   O(2) => x56_out_30,
   O(3) => x56_out_31
);
W_reg_44_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x56_out_3,
   R => '0',
   Q => W_reg_44_3
);
W_reg_44_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_44_3_i_5_n_0,
   DI(1) => W_44_3_i_4_n_0,
   DI(2) => W_44_3_i_3_n_0,
   DI(3) => W_44_3_i_2_n_0,
   S(0) => W_44_3_i_9_n_0,
   S(1) => W_44_3_i_8_n_0,
   S(2) => W_44_3_i_7_n_0,
   S(3) => W_44_3_i_6_n_0,
   CO(0) => W_reg_44_3_i_1_n_3,
   CO(1) => W_reg_44_3_i_1_n_2,
   CO(2) => W_reg_44_3_i_1_n_1,
   CO(3) => W_reg_44_3_i_1_n_0,
   O(0) => x56_out_0,
   O(1) => x56_out_1,
   O(2) => x56_out_2,
   O(3) => x56_out_3
);
W_reg_44_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x56_out_4,
   R => '0',
   Q => W_reg_44_4
);
W_reg_44_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x56_out_5,
   R => '0',
   Q => W_reg_44_5
);
W_reg_44_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x56_out_6,
   R => '0',
   Q => W_reg_44_6
);
W_reg_44_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x56_out_7,
   R => '0',
   Q => W_reg_44_7
);
W_reg_44_7_i_1 : CARRY4
 port map (
   CI => W_reg_44_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_44_7_i_5_n_0,
   DI(1) => W_44_7_i_4_n_0,
   DI(2) => W_44_7_i_3_n_0,
   DI(3) => W_44_7_i_2_n_0,
   S(0) => W_44_7_i_9_n_0,
   S(1) => W_44_7_i_8_n_0,
   S(2) => W_44_7_i_7_n_0,
   S(3) => W_44_7_i_6_n_0,
   CO(0) => W_reg_44_7_i_1_n_3,
   CO(1) => W_reg_44_7_i_1_n_2,
   CO(2) => W_reg_44_7_i_1_n_1,
   CO(3) => W_reg_44_7_i_1_n_0,
   O(0) => x56_out_4,
   O(1) => x56_out_5,
   O(2) => x56_out_6,
   O(3) => x56_out_7
);
W_reg_44_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x56_out_8,
   R => '0',
   Q => W_reg_44_8
);
W_reg_44_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x56_out_9,
   R => '0',
   Q => W_reg_44_9
);
W_reg_45_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x53_out_0,
   R => '0',
   Q => W_reg_45_0
);
W_reg_45_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x53_out_10,
   R => '0',
   Q => W_reg_45_10
);
W_reg_45_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x53_out_11,
   R => '0',
   Q => W_reg_45_11
);
W_reg_45_11_i_1 : CARRY4
 port map (
   CI => W_reg_45_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_45_11_i_5_n_0,
   DI(1) => W_45_11_i_4_n_0,
   DI(2) => W_45_11_i_3_n_0,
   DI(3) => W_45_11_i_2_n_0,
   S(0) => W_45_11_i_9_n_0,
   S(1) => W_45_11_i_8_n_0,
   S(2) => W_45_11_i_7_n_0,
   S(3) => W_45_11_i_6_n_0,
   CO(0) => W_reg_45_11_i_1_n_3,
   CO(1) => W_reg_45_11_i_1_n_2,
   CO(2) => W_reg_45_11_i_1_n_1,
   CO(3) => W_reg_45_11_i_1_n_0,
   O(0) => x53_out_8,
   O(1) => x53_out_9,
   O(2) => x53_out_10,
   O(3) => x53_out_11
);
W_reg_45_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x53_out_12,
   R => '0',
   Q => W_reg_45_12
);
W_reg_45_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x53_out_13,
   R => '0',
   Q => W_reg_45_13
);
W_reg_45_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x53_out_14,
   R => '0',
   Q => W_reg_45_14
);
W_reg_45_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x53_out_15,
   R => '0',
   Q => W_reg_45_15
);
W_reg_45_15_i_1 : CARRY4
 port map (
   CI => W_reg_45_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_45_15_i_5_n_0,
   DI(1) => W_45_15_i_4_n_0,
   DI(2) => W_45_15_i_3_n_0,
   DI(3) => W_45_15_i_2_n_0,
   S(0) => W_45_15_i_9_n_0,
   S(1) => W_45_15_i_8_n_0,
   S(2) => W_45_15_i_7_n_0,
   S(3) => W_45_15_i_6_n_0,
   CO(0) => W_reg_45_15_i_1_n_3,
   CO(1) => W_reg_45_15_i_1_n_2,
   CO(2) => W_reg_45_15_i_1_n_1,
   CO(3) => W_reg_45_15_i_1_n_0,
   O(0) => x53_out_12,
   O(1) => x53_out_13,
   O(2) => x53_out_14,
   O(3) => x53_out_15
);
W_reg_45_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x53_out_16,
   R => '0',
   Q => W_reg_45_16
);
W_reg_45_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x53_out_17,
   R => '0',
   Q => W_reg_45_17
);
W_reg_45_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x53_out_18,
   R => '0',
   Q => W_reg_45_18
);
W_reg_45_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x53_out_19,
   R => '0',
   Q => W_reg_45_19
);
W_reg_45_19_i_1 : CARRY4
 port map (
   CI => W_reg_45_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_45_19_i_5_n_0,
   DI(1) => W_45_19_i_4_n_0,
   DI(2) => W_45_19_i_3_n_0,
   DI(3) => W_45_19_i_2_n_0,
   S(0) => W_45_19_i_9_n_0,
   S(1) => W_45_19_i_8_n_0,
   S(2) => W_45_19_i_7_n_0,
   S(3) => W_45_19_i_6_n_0,
   CO(0) => W_reg_45_19_i_1_n_3,
   CO(1) => W_reg_45_19_i_1_n_2,
   CO(2) => W_reg_45_19_i_1_n_1,
   CO(3) => W_reg_45_19_i_1_n_0,
   O(0) => x53_out_16,
   O(1) => x53_out_17,
   O(2) => x53_out_18,
   O(3) => x53_out_19
);
W_reg_45_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x53_out_1,
   R => '0',
   Q => W_reg_45_1
);
W_reg_45_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x53_out_20,
   R => '0',
   Q => W_reg_45_20
);
W_reg_45_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x53_out_21,
   R => '0',
   Q => W_reg_45_21
);
W_reg_45_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x53_out_22,
   R => '0',
   Q => W_reg_45_22
);
W_reg_45_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x53_out_23,
   R => '0',
   Q => W_reg_45_23
);
W_reg_45_23_i_1 : CARRY4
 port map (
   CI => W_reg_45_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_45_23_i_5_n_0,
   DI(1) => W_45_23_i_4_n_0,
   DI(2) => W_45_23_i_3_n_0,
   DI(3) => W_45_23_i_2_n_0,
   S(0) => W_45_23_i_9_n_0,
   S(1) => W_45_23_i_8_n_0,
   S(2) => W_45_23_i_7_n_0,
   S(3) => W_45_23_i_6_n_0,
   CO(0) => W_reg_45_23_i_1_n_3,
   CO(1) => W_reg_45_23_i_1_n_2,
   CO(2) => W_reg_45_23_i_1_n_1,
   CO(3) => W_reg_45_23_i_1_n_0,
   O(0) => x53_out_20,
   O(1) => x53_out_21,
   O(2) => x53_out_22,
   O(3) => x53_out_23
);
W_reg_45_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x53_out_24,
   R => '0',
   Q => W_reg_45_24
);
W_reg_45_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x53_out_25,
   R => '0',
   Q => W_reg_45_25
);
W_reg_45_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x53_out_26,
   R => '0',
   Q => W_reg_45_26
);
W_reg_45_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x53_out_27,
   R => '0',
   Q => W_reg_45_27
);
W_reg_45_27_i_1 : CARRY4
 port map (
   CI => W_reg_45_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_45_27_i_5_n_0,
   DI(1) => W_45_27_i_4_n_0,
   DI(2) => W_45_27_i_3_n_0,
   DI(3) => W_45_27_i_2_n_0,
   S(0) => W_45_27_i_9_n_0,
   S(1) => W_45_27_i_8_n_0,
   S(2) => W_45_27_i_7_n_0,
   S(3) => W_45_27_i_6_n_0,
   CO(0) => W_reg_45_27_i_1_n_3,
   CO(1) => W_reg_45_27_i_1_n_2,
   CO(2) => W_reg_45_27_i_1_n_1,
   CO(3) => W_reg_45_27_i_1_n_0,
   O(0) => x53_out_24,
   O(1) => x53_out_25,
   O(2) => x53_out_26,
   O(3) => x53_out_27
);
W_reg_45_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x53_out_28,
   R => '0',
   Q => W_reg_45_28
);
W_reg_45_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x53_out_29,
   R => '0',
   Q => W_reg_45_29
);
W_reg_45_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x53_out_2,
   R => '0',
   Q => W_reg_45_2
);
W_reg_45_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x53_out_30,
   R => '0',
   Q => W_reg_45_30
);
W_reg_45_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x53_out_31,
   R => '0',
   Q => W_reg_45_31
);
W_reg_45_31_i_1 : CARRY4
 port map (
   CI => W_reg_45_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_45_31_i_4_n_0,
   DI(1) => W_45_31_i_3_n_0,
   DI(2) => W_45_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_45_31_i_8_n_0,
   S(1) => W_45_31_i_7_n_0,
   S(2) => W_45_31_i_6_n_0,
   S(3) => W_45_31_i_5_n_0,
   CO(0) => W_reg_45_31_i_1_n_3,
   CO(1) => W_reg_45_31_i_1_n_2,
   CO(2) => W_reg_45_31_i_1_n_1,
   CO(3) => NLW_W_reg_45_31_i_1_CO_UNCONNECTED_3,
   O(0) => x53_out_28,
   O(1) => x53_out_29,
   O(2) => x53_out_30,
   O(3) => x53_out_31
);
W_reg_45_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x53_out_3,
   R => '0',
   Q => W_reg_45_3
);
W_reg_45_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_45_3_i_5_n_0,
   DI(1) => W_45_3_i_4_n_0,
   DI(2) => W_45_3_i_3_n_0,
   DI(3) => W_45_3_i_2_n_0,
   S(0) => W_45_3_i_9_n_0,
   S(1) => W_45_3_i_8_n_0,
   S(2) => W_45_3_i_7_n_0,
   S(3) => W_45_3_i_6_n_0,
   CO(0) => W_reg_45_3_i_1_n_3,
   CO(1) => W_reg_45_3_i_1_n_2,
   CO(2) => W_reg_45_3_i_1_n_1,
   CO(3) => W_reg_45_3_i_1_n_0,
   O(0) => x53_out_0,
   O(1) => x53_out_1,
   O(2) => x53_out_2,
   O(3) => x53_out_3
);
W_reg_45_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x53_out_4,
   R => '0',
   Q => W_reg_45_4
);
W_reg_45_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x53_out_5,
   R => '0',
   Q => W_reg_45_5
);
W_reg_45_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x53_out_6,
   R => '0',
   Q => W_reg_45_6
);
W_reg_45_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x53_out_7,
   R => '0',
   Q => W_reg_45_7
);
W_reg_45_7_i_1 : CARRY4
 port map (
   CI => W_reg_45_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_45_7_i_5_n_0,
   DI(1) => W_45_7_i_4_n_0,
   DI(2) => W_45_7_i_3_n_0,
   DI(3) => W_45_7_i_2_n_0,
   S(0) => W_45_7_i_9_n_0,
   S(1) => W_45_7_i_8_n_0,
   S(2) => W_45_7_i_7_n_0,
   S(3) => W_45_7_i_6_n_0,
   CO(0) => W_reg_45_7_i_1_n_3,
   CO(1) => W_reg_45_7_i_1_n_2,
   CO(2) => W_reg_45_7_i_1_n_1,
   CO(3) => W_reg_45_7_i_1_n_0,
   O(0) => x53_out_4,
   O(1) => x53_out_5,
   O(2) => x53_out_6,
   O(3) => x53_out_7
);
W_reg_45_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x53_out_8,
   R => '0',
   Q => W_reg_45_8
);
W_reg_45_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x53_out_9,
   R => '0',
   Q => W_reg_45_9
);
W_reg_46_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x50_out_0,
   R => '0',
   Q => W_reg_46_0
);
W_reg_46_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x50_out_10,
   R => '0',
   Q => W_reg_46_10
);
W_reg_46_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x50_out_11,
   R => '0',
   Q => W_reg_46_11
);
W_reg_46_11_i_1 : CARRY4
 port map (
   CI => W_reg_46_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_46_11_i_5_n_0,
   DI(1) => W_46_11_i_4_n_0,
   DI(2) => W_46_11_i_3_n_0,
   DI(3) => W_46_11_i_2_n_0,
   S(0) => W_46_11_i_9_n_0,
   S(1) => W_46_11_i_8_n_0,
   S(2) => W_46_11_i_7_n_0,
   S(3) => W_46_11_i_6_n_0,
   CO(0) => W_reg_46_11_i_1_n_3,
   CO(1) => W_reg_46_11_i_1_n_2,
   CO(2) => W_reg_46_11_i_1_n_1,
   CO(3) => W_reg_46_11_i_1_n_0,
   O(0) => x50_out_8,
   O(1) => x50_out_9,
   O(2) => x50_out_10,
   O(3) => x50_out_11
);
W_reg_46_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x50_out_12,
   R => '0',
   Q => W_reg_46_12
);
W_reg_46_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x50_out_13,
   R => '0',
   Q => W_reg_46_13
);
W_reg_46_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x50_out_14,
   R => '0',
   Q => W_reg_46_14
);
W_reg_46_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x50_out_15,
   R => '0',
   Q => W_reg_46_15
);
W_reg_46_15_i_1 : CARRY4
 port map (
   CI => W_reg_46_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_46_15_i_5_n_0,
   DI(1) => W_46_15_i_4_n_0,
   DI(2) => W_46_15_i_3_n_0,
   DI(3) => W_46_15_i_2_n_0,
   S(0) => W_46_15_i_9_n_0,
   S(1) => W_46_15_i_8_n_0,
   S(2) => W_46_15_i_7_n_0,
   S(3) => W_46_15_i_6_n_0,
   CO(0) => W_reg_46_15_i_1_n_3,
   CO(1) => W_reg_46_15_i_1_n_2,
   CO(2) => W_reg_46_15_i_1_n_1,
   CO(3) => W_reg_46_15_i_1_n_0,
   O(0) => x50_out_12,
   O(1) => x50_out_13,
   O(2) => x50_out_14,
   O(3) => x50_out_15
);
W_reg_46_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x50_out_16,
   R => '0',
   Q => W_reg_46_16
);
W_reg_46_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x50_out_17,
   R => '0',
   Q => W_reg_46_17
);
W_reg_46_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x50_out_18,
   R => '0',
   Q => W_reg_46_18
);
W_reg_46_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x50_out_19,
   R => '0',
   Q => W_reg_46_19
);
W_reg_46_19_i_1 : CARRY4
 port map (
   CI => W_reg_46_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_46_19_i_5_n_0,
   DI(1) => W_46_19_i_4_n_0,
   DI(2) => W_46_19_i_3_n_0,
   DI(3) => W_46_19_i_2_n_0,
   S(0) => W_46_19_i_9_n_0,
   S(1) => W_46_19_i_8_n_0,
   S(2) => W_46_19_i_7_n_0,
   S(3) => W_46_19_i_6_n_0,
   CO(0) => W_reg_46_19_i_1_n_3,
   CO(1) => W_reg_46_19_i_1_n_2,
   CO(2) => W_reg_46_19_i_1_n_1,
   CO(3) => W_reg_46_19_i_1_n_0,
   O(0) => x50_out_16,
   O(1) => x50_out_17,
   O(2) => x50_out_18,
   O(3) => x50_out_19
);
W_reg_46_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x50_out_1,
   R => '0',
   Q => W_reg_46_1
);
W_reg_46_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x50_out_20,
   R => '0',
   Q => W_reg_46_20
);
W_reg_46_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x50_out_21,
   R => '0',
   Q => W_reg_46_21
);
W_reg_46_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x50_out_22,
   R => '0',
   Q => W_reg_46_22
);
W_reg_46_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x50_out_23,
   R => '0',
   Q => W_reg_46_23
);
W_reg_46_23_i_1 : CARRY4
 port map (
   CI => W_reg_46_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_46_23_i_5_n_0,
   DI(1) => W_46_23_i_4_n_0,
   DI(2) => W_46_23_i_3_n_0,
   DI(3) => W_46_23_i_2_n_0,
   S(0) => W_46_23_i_9_n_0,
   S(1) => W_46_23_i_8_n_0,
   S(2) => W_46_23_i_7_n_0,
   S(3) => W_46_23_i_6_n_0,
   CO(0) => W_reg_46_23_i_1_n_3,
   CO(1) => W_reg_46_23_i_1_n_2,
   CO(2) => W_reg_46_23_i_1_n_1,
   CO(3) => W_reg_46_23_i_1_n_0,
   O(0) => x50_out_20,
   O(1) => x50_out_21,
   O(2) => x50_out_22,
   O(3) => x50_out_23
);
W_reg_46_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x50_out_24,
   R => '0',
   Q => W_reg_46_24
);
W_reg_46_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x50_out_25,
   R => '0',
   Q => W_reg_46_25
);
W_reg_46_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x50_out_26,
   R => '0',
   Q => W_reg_46_26
);
W_reg_46_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x50_out_27,
   R => '0',
   Q => W_reg_46_27
);
W_reg_46_27_i_1 : CARRY4
 port map (
   CI => W_reg_46_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_46_27_i_5_n_0,
   DI(1) => W_46_27_i_4_n_0,
   DI(2) => W_46_27_i_3_n_0,
   DI(3) => W_46_27_i_2_n_0,
   S(0) => W_46_27_i_9_n_0,
   S(1) => W_46_27_i_8_n_0,
   S(2) => W_46_27_i_7_n_0,
   S(3) => W_46_27_i_6_n_0,
   CO(0) => W_reg_46_27_i_1_n_3,
   CO(1) => W_reg_46_27_i_1_n_2,
   CO(2) => W_reg_46_27_i_1_n_1,
   CO(3) => W_reg_46_27_i_1_n_0,
   O(0) => x50_out_24,
   O(1) => x50_out_25,
   O(2) => x50_out_26,
   O(3) => x50_out_27
);
W_reg_46_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x50_out_28,
   R => '0',
   Q => W_reg_46_28
);
W_reg_46_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x50_out_29,
   R => '0',
   Q => W_reg_46_29
);
W_reg_46_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x50_out_2,
   R => '0',
   Q => W_reg_46_2
);
W_reg_46_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x50_out_30,
   R => '0',
   Q => W_reg_46_30
);
W_reg_46_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x50_out_31,
   R => '0',
   Q => W_reg_46_31
);
W_reg_46_31_i_1 : CARRY4
 port map (
   CI => W_reg_46_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_46_31_i_4_n_0,
   DI(1) => W_46_31_i_3_n_0,
   DI(2) => W_46_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_46_31_i_8_n_0,
   S(1) => W_46_31_i_7_n_0,
   S(2) => W_46_31_i_6_n_0,
   S(3) => W_46_31_i_5_n_0,
   CO(0) => W_reg_46_31_i_1_n_3,
   CO(1) => W_reg_46_31_i_1_n_2,
   CO(2) => W_reg_46_31_i_1_n_1,
   CO(3) => NLW_W_reg_46_31_i_1_CO_UNCONNECTED_3,
   O(0) => x50_out_28,
   O(1) => x50_out_29,
   O(2) => x50_out_30,
   O(3) => x50_out_31
);
W_reg_46_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x50_out_3,
   R => '0',
   Q => W_reg_46_3
);
W_reg_46_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_46_3_i_5_n_0,
   DI(1) => W_46_3_i_4_n_0,
   DI(2) => W_46_3_i_3_n_0,
   DI(3) => W_46_3_i_2_n_0,
   S(0) => W_46_3_i_9_n_0,
   S(1) => W_46_3_i_8_n_0,
   S(2) => W_46_3_i_7_n_0,
   S(3) => W_46_3_i_6_n_0,
   CO(0) => W_reg_46_3_i_1_n_3,
   CO(1) => W_reg_46_3_i_1_n_2,
   CO(2) => W_reg_46_3_i_1_n_1,
   CO(3) => W_reg_46_3_i_1_n_0,
   O(0) => x50_out_0,
   O(1) => x50_out_1,
   O(2) => x50_out_2,
   O(3) => x50_out_3
);
W_reg_46_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x50_out_4,
   R => '0',
   Q => W_reg_46_4
);
W_reg_46_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x50_out_5,
   R => '0',
   Q => W_reg_46_5
);
W_reg_46_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x50_out_6,
   R => '0',
   Q => W_reg_46_6
);
W_reg_46_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x50_out_7,
   R => '0',
   Q => W_reg_46_7
);
W_reg_46_7_i_1 : CARRY4
 port map (
   CI => W_reg_46_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_46_7_i_5_n_0,
   DI(1) => W_46_7_i_4_n_0,
   DI(2) => W_46_7_i_3_n_0,
   DI(3) => W_46_7_i_2_n_0,
   S(0) => W_46_7_i_9_n_0,
   S(1) => W_46_7_i_8_n_0,
   S(2) => W_46_7_i_7_n_0,
   S(3) => W_46_7_i_6_n_0,
   CO(0) => W_reg_46_7_i_1_n_3,
   CO(1) => W_reg_46_7_i_1_n_2,
   CO(2) => W_reg_46_7_i_1_n_1,
   CO(3) => W_reg_46_7_i_1_n_0,
   O(0) => x50_out_4,
   O(1) => x50_out_5,
   O(2) => x50_out_6,
   O(3) => x50_out_7
);
W_reg_46_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x50_out_8,
   R => '0',
   Q => W_reg_46_8
);
W_reg_46_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x50_out_9,
   R => '0',
   Q => W_reg_46_9
);
W_reg_47_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x47_out_0,
   R => '0',
   Q => W_reg_47_0
);
W_reg_47_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x47_out_10,
   R => '0',
   Q => W_reg_47_10
);
W_reg_47_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x47_out_11,
   R => '0',
   Q => W_reg_47_11
);
W_reg_47_11_i_1 : CARRY4
 port map (
   CI => W_reg_47_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_47_11_i_5_n_0,
   DI(1) => W_47_11_i_4_n_0,
   DI(2) => W_47_11_i_3_n_0,
   DI(3) => W_47_11_i_2_n_0,
   S(0) => W_47_11_i_9_n_0,
   S(1) => W_47_11_i_8_n_0,
   S(2) => W_47_11_i_7_n_0,
   S(3) => W_47_11_i_6_n_0,
   CO(0) => W_reg_47_11_i_1_n_3,
   CO(1) => W_reg_47_11_i_1_n_2,
   CO(2) => W_reg_47_11_i_1_n_1,
   CO(3) => W_reg_47_11_i_1_n_0,
   O(0) => x47_out_8,
   O(1) => x47_out_9,
   O(2) => x47_out_10,
   O(3) => x47_out_11
);
W_reg_47_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x47_out_12,
   R => '0',
   Q => W_reg_47_12
);
W_reg_47_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x47_out_13,
   R => '0',
   Q => W_reg_47_13
);
W_reg_47_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x47_out_14,
   R => '0',
   Q => W_reg_47_14
);
W_reg_47_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x47_out_15,
   R => '0',
   Q => W_reg_47_15
);
W_reg_47_15_i_1 : CARRY4
 port map (
   CI => W_reg_47_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_47_15_i_5_n_0,
   DI(1) => W_47_15_i_4_n_0,
   DI(2) => W_47_15_i_3_n_0,
   DI(3) => W_47_15_i_2_n_0,
   S(0) => W_47_15_i_9_n_0,
   S(1) => W_47_15_i_8_n_0,
   S(2) => W_47_15_i_7_n_0,
   S(3) => W_47_15_i_6_n_0,
   CO(0) => W_reg_47_15_i_1_n_3,
   CO(1) => W_reg_47_15_i_1_n_2,
   CO(2) => W_reg_47_15_i_1_n_1,
   CO(3) => W_reg_47_15_i_1_n_0,
   O(0) => x47_out_12,
   O(1) => x47_out_13,
   O(2) => x47_out_14,
   O(3) => x47_out_15
);
W_reg_47_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x47_out_16,
   R => '0',
   Q => W_reg_47_16
);
W_reg_47_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x47_out_17,
   R => '0',
   Q => W_reg_47_17
);
W_reg_47_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x47_out_18,
   R => '0',
   Q => W_reg_47_18
);
W_reg_47_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x47_out_19,
   R => '0',
   Q => W_reg_47_19
);
W_reg_47_19_i_1 : CARRY4
 port map (
   CI => W_reg_47_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_47_19_i_5_n_0,
   DI(1) => W_47_19_i_4_n_0,
   DI(2) => W_47_19_i_3_n_0,
   DI(3) => W_47_19_i_2_n_0,
   S(0) => W_47_19_i_9_n_0,
   S(1) => W_47_19_i_8_n_0,
   S(2) => W_47_19_i_7_n_0,
   S(3) => W_47_19_i_6_n_0,
   CO(0) => W_reg_47_19_i_1_n_3,
   CO(1) => W_reg_47_19_i_1_n_2,
   CO(2) => W_reg_47_19_i_1_n_1,
   CO(3) => W_reg_47_19_i_1_n_0,
   O(0) => x47_out_16,
   O(1) => x47_out_17,
   O(2) => x47_out_18,
   O(3) => x47_out_19
);
W_reg_47_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x47_out_1,
   R => '0',
   Q => W_reg_47_1
);
W_reg_47_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x47_out_20,
   R => '0',
   Q => W_reg_47_20
);
W_reg_47_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x47_out_21,
   R => '0',
   Q => W_reg_47_21
);
W_reg_47_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x47_out_22,
   R => '0',
   Q => W_reg_47_22
);
W_reg_47_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x47_out_23,
   R => '0',
   Q => W_reg_47_23
);
W_reg_47_23_i_1 : CARRY4
 port map (
   CI => W_reg_47_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_47_23_i_5_n_0,
   DI(1) => W_47_23_i_4_n_0,
   DI(2) => W_47_23_i_3_n_0,
   DI(3) => W_47_23_i_2_n_0,
   S(0) => W_47_23_i_9_n_0,
   S(1) => W_47_23_i_8_n_0,
   S(2) => W_47_23_i_7_n_0,
   S(3) => W_47_23_i_6_n_0,
   CO(0) => W_reg_47_23_i_1_n_3,
   CO(1) => W_reg_47_23_i_1_n_2,
   CO(2) => W_reg_47_23_i_1_n_1,
   CO(3) => W_reg_47_23_i_1_n_0,
   O(0) => x47_out_20,
   O(1) => x47_out_21,
   O(2) => x47_out_22,
   O(3) => x47_out_23
);
W_reg_47_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x47_out_24,
   R => '0',
   Q => W_reg_47_24
);
W_reg_47_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x47_out_25,
   R => '0',
   Q => W_reg_47_25
);
W_reg_47_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x47_out_26,
   R => '0',
   Q => W_reg_47_26
);
W_reg_47_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x47_out_27,
   R => '0',
   Q => W_reg_47_27
);
W_reg_47_27_i_1 : CARRY4
 port map (
   CI => W_reg_47_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_47_27_i_5_n_0,
   DI(1) => W_47_27_i_4_n_0,
   DI(2) => W_47_27_i_3_n_0,
   DI(3) => W_47_27_i_2_n_0,
   S(0) => W_47_27_i_9_n_0,
   S(1) => W_47_27_i_8_n_0,
   S(2) => W_47_27_i_7_n_0,
   S(3) => W_47_27_i_6_n_0,
   CO(0) => W_reg_47_27_i_1_n_3,
   CO(1) => W_reg_47_27_i_1_n_2,
   CO(2) => W_reg_47_27_i_1_n_1,
   CO(3) => W_reg_47_27_i_1_n_0,
   O(0) => x47_out_24,
   O(1) => x47_out_25,
   O(2) => x47_out_26,
   O(3) => x47_out_27
);
W_reg_47_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x47_out_28,
   R => '0',
   Q => W_reg_47_28
);
W_reg_47_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x47_out_29,
   R => '0',
   Q => W_reg_47_29
);
W_reg_47_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x47_out_2,
   R => '0',
   Q => W_reg_47_2
);
W_reg_47_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x47_out_30,
   R => '0',
   Q => W_reg_47_30
);
W_reg_47_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x47_out_31,
   R => '0',
   Q => W_reg_47_31
);
W_reg_47_31_i_1 : CARRY4
 port map (
   CI => W_reg_47_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_47_31_i_4_n_0,
   DI(1) => W_47_31_i_3_n_0,
   DI(2) => W_47_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_47_31_i_8_n_0,
   S(1) => W_47_31_i_7_n_0,
   S(2) => W_47_31_i_6_n_0,
   S(3) => W_47_31_i_5_n_0,
   CO(0) => W_reg_47_31_i_1_n_3,
   CO(1) => W_reg_47_31_i_1_n_2,
   CO(2) => W_reg_47_31_i_1_n_1,
   CO(3) => NLW_W_reg_47_31_i_1_CO_UNCONNECTED_3,
   O(0) => x47_out_28,
   O(1) => x47_out_29,
   O(2) => x47_out_30,
   O(3) => x47_out_31
);
W_reg_47_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x47_out_3,
   R => '0',
   Q => W_reg_47_3
);
W_reg_47_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_47_3_i_5_n_0,
   DI(1) => W_47_3_i_4_n_0,
   DI(2) => W_47_3_i_3_n_0,
   DI(3) => W_47_3_i_2_n_0,
   S(0) => W_47_3_i_9_n_0,
   S(1) => W_47_3_i_8_n_0,
   S(2) => W_47_3_i_7_n_0,
   S(3) => W_47_3_i_6_n_0,
   CO(0) => W_reg_47_3_i_1_n_3,
   CO(1) => W_reg_47_3_i_1_n_2,
   CO(2) => W_reg_47_3_i_1_n_1,
   CO(3) => W_reg_47_3_i_1_n_0,
   O(0) => x47_out_0,
   O(1) => x47_out_1,
   O(2) => x47_out_2,
   O(3) => x47_out_3
);
W_reg_47_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x47_out_4,
   R => '0',
   Q => W_reg_47_4
);
W_reg_47_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x47_out_5,
   R => '0',
   Q => W_reg_47_5
);
W_reg_47_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x47_out_6,
   R => '0',
   Q => W_reg_47_6
);
W_reg_47_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x47_out_7,
   R => '0',
   Q => W_reg_47_7
);
W_reg_47_7_i_1 : CARRY4
 port map (
   CI => W_reg_47_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_47_7_i_5_n_0,
   DI(1) => W_47_7_i_4_n_0,
   DI(2) => W_47_7_i_3_n_0,
   DI(3) => W_47_7_i_2_n_0,
   S(0) => W_47_7_i_9_n_0,
   S(1) => W_47_7_i_8_n_0,
   S(2) => W_47_7_i_7_n_0,
   S(3) => W_47_7_i_6_n_0,
   CO(0) => W_reg_47_7_i_1_n_3,
   CO(1) => W_reg_47_7_i_1_n_2,
   CO(2) => W_reg_47_7_i_1_n_1,
   CO(3) => W_reg_47_7_i_1_n_0,
   O(0) => x47_out_4,
   O(1) => x47_out_5,
   O(2) => x47_out_6,
   O(3) => x47_out_7
);
W_reg_47_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x47_out_8,
   R => '0',
   Q => W_reg_47_8
);
W_reg_47_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_32_0,
   D => x47_out_9,
   R => '0',
   Q => W_reg_47_9
);
W_reg_48_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x44_out_0,
   R => '0',
   Q => W_reg_48_0
);
W_reg_48_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x44_out_10,
   R => '0',
   Q => W_reg_48_10
);
W_reg_48_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x44_out_11,
   R => '0',
   Q => W_reg_48_11
);
W_reg_48_11_i_1 : CARRY4
 port map (
   CI => W_reg_48_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_48_11_i_5_n_0,
   DI(1) => W_48_11_i_4_n_0,
   DI(2) => W_48_11_i_3_n_0,
   DI(3) => W_48_11_i_2_n_0,
   S(0) => W_48_11_i_9_n_0,
   S(1) => W_48_11_i_8_n_0,
   S(2) => W_48_11_i_7_n_0,
   S(3) => W_48_11_i_6_n_0,
   CO(0) => W_reg_48_11_i_1_n_3,
   CO(1) => W_reg_48_11_i_1_n_2,
   CO(2) => W_reg_48_11_i_1_n_1,
   CO(3) => W_reg_48_11_i_1_n_0,
   O(0) => x44_out_8,
   O(1) => x44_out_9,
   O(2) => x44_out_10,
   O(3) => x44_out_11
);
W_reg_48_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x44_out_12,
   R => '0',
   Q => W_reg_48_12
);
W_reg_48_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x44_out_13,
   R => '0',
   Q => W_reg_48_13
);
W_reg_48_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x44_out_14,
   R => '0',
   Q => W_reg_48_14
);
W_reg_48_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x44_out_15,
   R => '0',
   Q => W_reg_48_15
);
W_reg_48_15_i_1 : CARRY4
 port map (
   CI => W_reg_48_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_48_15_i_5_n_0,
   DI(1) => W_48_15_i_4_n_0,
   DI(2) => W_48_15_i_3_n_0,
   DI(3) => W_48_15_i_2_n_0,
   S(0) => W_48_15_i_9_n_0,
   S(1) => W_48_15_i_8_n_0,
   S(2) => W_48_15_i_7_n_0,
   S(3) => W_48_15_i_6_n_0,
   CO(0) => W_reg_48_15_i_1_n_3,
   CO(1) => W_reg_48_15_i_1_n_2,
   CO(2) => W_reg_48_15_i_1_n_1,
   CO(3) => W_reg_48_15_i_1_n_0,
   O(0) => x44_out_12,
   O(1) => x44_out_13,
   O(2) => x44_out_14,
   O(3) => x44_out_15
);
W_reg_48_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x44_out_16,
   R => '0',
   Q => W_reg_48_16
);
W_reg_48_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x44_out_17,
   R => '0',
   Q => W_reg_48_17
);
W_reg_48_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x44_out_18,
   R => '0',
   Q => W_reg_48_18
);
W_reg_48_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x44_out_19,
   R => '0',
   Q => W_reg_48_19
);
W_reg_48_19_i_1 : CARRY4
 port map (
   CI => W_reg_48_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_48_19_i_5_n_0,
   DI(1) => W_48_19_i_4_n_0,
   DI(2) => W_48_19_i_3_n_0,
   DI(3) => W_48_19_i_2_n_0,
   S(0) => W_48_19_i_9_n_0,
   S(1) => W_48_19_i_8_n_0,
   S(2) => W_48_19_i_7_n_0,
   S(3) => W_48_19_i_6_n_0,
   CO(0) => W_reg_48_19_i_1_n_3,
   CO(1) => W_reg_48_19_i_1_n_2,
   CO(2) => W_reg_48_19_i_1_n_1,
   CO(3) => W_reg_48_19_i_1_n_0,
   O(0) => x44_out_16,
   O(1) => x44_out_17,
   O(2) => x44_out_18,
   O(3) => x44_out_19
);
W_reg_48_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x44_out_1,
   R => '0',
   Q => W_reg_48_1
);
W_reg_48_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x44_out_20,
   R => '0',
   Q => W_reg_48_20
);
W_reg_48_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x44_out_21,
   R => '0',
   Q => W_reg_48_21
);
W_reg_48_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x44_out_22,
   R => '0',
   Q => W_reg_48_22
);
W_reg_48_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x44_out_23,
   R => '0',
   Q => W_reg_48_23
);
W_reg_48_23_i_1 : CARRY4
 port map (
   CI => W_reg_48_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_48_23_i_5_n_0,
   DI(1) => W_48_23_i_4_n_0,
   DI(2) => W_48_23_i_3_n_0,
   DI(3) => W_48_23_i_2_n_0,
   S(0) => W_48_23_i_9_n_0,
   S(1) => W_48_23_i_8_n_0,
   S(2) => W_48_23_i_7_n_0,
   S(3) => W_48_23_i_6_n_0,
   CO(0) => W_reg_48_23_i_1_n_3,
   CO(1) => W_reg_48_23_i_1_n_2,
   CO(2) => W_reg_48_23_i_1_n_1,
   CO(3) => W_reg_48_23_i_1_n_0,
   O(0) => x44_out_20,
   O(1) => x44_out_21,
   O(2) => x44_out_22,
   O(3) => x44_out_23
);
W_reg_48_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x44_out_24,
   R => '0',
   Q => W_reg_48_24
);
W_reg_48_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x44_out_25,
   R => '0',
   Q => W_reg_48_25
);
W_reg_48_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x44_out_26,
   R => '0',
   Q => W_reg_48_26
);
W_reg_48_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x44_out_27,
   R => '0',
   Q => W_reg_48_27
);
W_reg_48_27_i_1 : CARRY4
 port map (
   CI => W_reg_48_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_48_27_i_5_n_0,
   DI(1) => W_48_27_i_4_n_0,
   DI(2) => W_48_27_i_3_n_0,
   DI(3) => W_48_27_i_2_n_0,
   S(0) => W_48_27_i_9_n_0,
   S(1) => W_48_27_i_8_n_0,
   S(2) => W_48_27_i_7_n_0,
   S(3) => W_48_27_i_6_n_0,
   CO(0) => W_reg_48_27_i_1_n_3,
   CO(1) => W_reg_48_27_i_1_n_2,
   CO(2) => W_reg_48_27_i_1_n_1,
   CO(3) => W_reg_48_27_i_1_n_0,
   O(0) => x44_out_24,
   O(1) => x44_out_25,
   O(2) => x44_out_26,
   O(3) => x44_out_27
);
W_reg_48_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x44_out_28,
   R => '0',
   Q => W_reg_48_28
);
W_reg_48_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x44_out_29,
   R => '0',
   Q => W_reg_48_29
);
W_reg_48_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x44_out_2,
   R => '0',
   Q => W_reg_48_2
);
W_reg_48_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x44_out_30,
   R => '0',
   Q => W_reg_48_30
);
W_reg_48_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x44_out_31,
   R => '0',
   Q => W_reg_48_31
);
W_reg_48_31_i_2 : CARRY4
 port map (
   CI => W_reg_48_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_48_31_i_5_n_0,
   DI(1) => W_48_31_i_4_n_0,
   DI(2) => W_48_31_i_3_n_0,
   DI(3) => '0',
   S(0) => W_48_31_i_9_n_0,
   S(1) => W_48_31_i_8_n_0,
   S(2) => W_48_31_i_7_n_0,
   S(3) => W_48_31_i_6_n_0,
   CO(0) => W_reg_48_31_i_2_n_3,
   CO(1) => W_reg_48_31_i_2_n_2,
   CO(2) => W_reg_48_31_i_2_n_1,
   CO(3) => NLW_W_reg_48_31_i_2_CO_UNCONNECTED_3,
   O(0) => x44_out_28,
   O(1) => x44_out_29,
   O(2) => x44_out_30,
   O(3) => x44_out_31
);
W_reg_48_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x44_out_3,
   R => '0',
   Q => W_reg_48_3
);
W_reg_48_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_48_3_i_5_n_0,
   DI(1) => W_48_3_i_4_n_0,
   DI(2) => W_48_3_i_3_n_0,
   DI(3) => W_48_3_i_2_n_0,
   S(0) => W_48_3_i_9_n_0,
   S(1) => W_48_3_i_8_n_0,
   S(2) => W_48_3_i_7_n_0,
   S(3) => W_48_3_i_6_n_0,
   CO(0) => W_reg_48_3_i_1_n_3,
   CO(1) => W_reg_48_3_i_1_n_2,
   CO(2) => W_reg_48_3_i_1_n_1,
   CO(3) => W_reg_48_3_i_1_n_0,
   O(0) => x44_out_0,
   O(1) => x44_out_1,
   O(2) => x44_out_2,
   O(3) => x44_out_3
);
W_reg_48_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x44_out_4,
   R => '0',
   Q => W_reg_48_4
);
W_reg_48_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x44_out_5,
   R => '0',
   Q => W_reg_48_5
);
W_reg_48_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x44_out_6,
   R => '0',
   Q => W_reg_48_6
);
W_reg_48_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x44_out_7,
   R => '0',
   Q => W_reg_48_7
);
W_reg_48_7_i_1 : CARRY4
 port map (
   CI => W_reg_48_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_48_7_i_5_n_0,
   DI(1) => W_48_7_i_4_n_0,
   DI(2) => W_48_7_i_3_n_0,
   DI(3) => W_48_7_i_2_n_0,
   S(0) => W_48_7_i_9_n_0,
   S(1) => W_48_7_i_8_n_0,
   S(2) => W_48_7_i_7_n_0,
   S(3) => W_48_7_i_6_n_0,
   CO(0) => W_reg_48_7_i_1_n_3,
   CO(1) => W_reg_48_7_i_1_n_2,
   CO(2) => W_reg_48_7_i_1_n_1,
   CO(3) => W_reg_48_7_i_1_n_0,
   O(0) => x44_out_4,
   O(1) => x44_out_5,
   O(2) => x44_out_6,
   O(3) => x44_out_7
);
W_reg_48_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x44_out_8,
   R => '0',
   Q => W_reg_48_8
);
W_reg_48_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x44_out_9,
   R => '0',
   Q => W_reg_48_9
);
W_reg_49_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x41_out_0,
   R => '0',
   Q => W_reg_49_0
);
W_reg_49_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x41_out_10,
   R => '0',
   Q => W_reg_49_10
);
W_reg_49_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x41_out_11,
   R => '0',
   Q => W_reg_49_11
);
W_reg_49_11_i_1 : CARRY4
 port map (
   CI => W_reg_49_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_49_11_i_5_n_0,
   DI(1) => W_49_11_i_4_n_0,
   DI(2) => W_49_11_i_3_n_0,
   DI(3) => W_49_11_i_2_n_0,
   S(0) => W_49_11_i_9_n_0,
   S(1) => W_49_11_i_8_n_0,
   S(2) => W_49_11_i_7_n_0,
   S(3) => W_49_11_i_6_n_0,
   CO(0) => W_reg_49_11_i_1_n_3,
   CO(1) => W_reg_49_11_i_1_n_2,
   CO(2) => W_reg_49_11_i_1_n_1,
   CO(3) => W_reg_49_11_i_1_n_0,
   O(0) => x41_out_8,
   O(1) => x41_out_9,
   O(2) => x41_out_10,
   O(3) => x41_out_11
);
W_reg_49_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x41_out_12,
   R => '0',
   Q => W_reg_49_12
);
W_reg_49_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x41_out_13,
   R => '0',
   Q => W_reg_49_13
);
W_reg_49_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x41_out_14,
   R => '0',
   Q => W_reg_49_14
);
W_reg_49_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x41_out_15,
   R => '0',
   Q => W_reg_49_15
);
W_reg_49_15_i_1 : CARRY4
 port map (
   CI => W_reg_49_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_49_15_i_5_n_0,
   DI(1) => W_49_15_i_4_n_0,
   DI(2) => W_49_15_i_3_n_0,
   DI(3) => W_49_15_i_2_n_0,
   S(0) => W_49_15_i_9_n_0,
   S(1) => W_49_15_i_8_n_0,
   S(2) => W_49_15_i_7_n_0,
   S(3) => W_49_15_i_6_n_0,
   CO(0) => W_reg_49_15_i_1_n_3,
   CO(1) => W_reg_49_15_i_1_n_2,
   CO(2) => W_reg_49_15_i_1_n_1,
   CO(3) => W_reg_49_15_i_1_n_0,
   O(0) => x41_out_12,
   O(1) => x41_out_13,
   O(2) => x41_out_14,
   O(3) => x41_out_15
);
W_reg_49_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x41_out_16,
   R => '0',
   Q => W_reg_49_16
);
W_reg_49_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x41_out_17,
   R => '0',
   Q => W_reg_49_17
);
W_reg_49_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x41_out_18,
   R => '0',
   Q => W_reg_49_18
);
W_reg_49_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x41_out_19,
   R => '0',
   Q => W_reg_49_19
);
W_reg_49_19_i_1 : CARRY4
 port map (
   CI => W_reg_49_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_49_19_i_5_n_0,
   DI(1) => W_49_19_i_4_n_0,
   DI(2) => W_49_19_i_3_n_0,
   DI(3) => W_49_19_i_2_n_0,
   S(0) => W_49_19_i_9_n_0,
   S(1) => W_49_19_i_8_n_0,
   S(2) => W_49_19_i_7_n_0,
   S(3) => W_49_19_i_6_n_0,
   CO(0) => W_reg_49_19_i_1_n_3,
   CO(1) => W_reg_49_19_i_1_n_2,
   CO(2) => W_reg_49_19_i_1_n_1,
   CO(3) => W_reg_49_19_i_1_n_0,
   O(0) => x41_out_16,
   O(1) => x41_out_17,
   O(2) => x41_out_18,
   O(3) => x41_out_19
);
W_reg_49_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x41_out_1,
   R => '0',
   Q => W_reg_49_1
);
W_reg_49_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x41_out_20,
   R => '0',
   Q => W_reg_49_20
);
W_reg_49_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x41_out_21,
   R => '0',
   Q => W_reg_49_21
);
W_reg_49_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x41_out_22,
   R => '0',
   Q => W_reg_49_22
);
W_reg_49_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x41_out_23,
   R => '0',
   Q => W_reg_49_23
);
W_reg_49_23_i_1 : CARRY4
 port map (
   CI => W_reg_49_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_49_23_i_5_n_0,
   DI(1) => W_49_23_i_4_n_0,
   DI(2) => W_49_23_i_3_n_0,
   DI(3) => W_49_23_i_2_n_0,
   S(0) => W_49_23_i_9_n_0,
   S(1) => W_49_23_i_8_n_0,
   S(2) => W_49_23_i_7_n_0,
   S(3) => W_49_23_i_6_n_0,
   CO(0) => W_reg_49_23_i_1_n_3,
   CO(1) => W_reg_49_23_i_1_n_2,
   CO(2) => W_reg_49_23_i_1_n_1,
   CO(3) => W_reg_49_23_i_1_n_0,
   O(0) => x41_out_20,
   O(1) => x41_out_21,
   O(2) => x41_out_22,
   O(3) => x41_out_23
);
W_reg_49_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x41_out_24,
   R => '0',
   Q => W_reg_49_24
);
W_reg_49_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x41_out_25,
   R => '0',
   Q => W_reg_49_25
);
W_reg_49_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x41_out_26,
   R => '0',
   Q => W_reg_49_26
);
W_reg_49_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x41_out_27,
   R => '0',
   Q => W_reg_49_27
);
W_reg_49_27_i_1 : CARRY4
 port map (
   CI => W_reg_49_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_49_27_i_5_n_0,
   DI(1) => W_49_27_i_4_n_0,
   DI(2) => W_49_27_i_3_n_0,
   DI(3) => W_49_27_i_2_n_0,
   S(0) => W_49_27_i_9_n_0,
   S(1) => W_49_27_i_8_n_0,
   S(2) => W_49_27_i_7_n_0,
   S(3) => W_49_27_i_6_n_0,
   CO(0) => W_reg_49_27_i_1_n_3,
   CO(1) => W_reg_49_27_i_1_n_2,
   CO(2) => W_reg_49_27_i_1_n_1,
   CO(3) => W_reg_49_27_i_1_n_0,
   O(0) => x41_out_24,
   O(1) => x41_out_25,
   O(2) => x41_out_26,
   O(3) => x41_out_27
);
W_reg_49_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x41_out_28,
   R => '0',
   Q => W_reg_49_28
);
W_reg_49_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x41_out_29,
   R => '0',
   Q => W_reg_49_29
);
W_reg_49_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x41_out_2,
   R => '0',
   Q => W_reg_49_2
);
W_reg_49_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x41_out_30,
   R => '0',
   Q => W_reg_49_30
);
W_reg_49_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x41_out_31,
   R => '0',
   Q => W_reg_49_31
);
W_reg_49_31_i_1 : CARRY4
 port map (
   CI => W_reg_49_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_49_31_i_4_n_0,
   DI(1) => W_49_31_i_3_n_0,
   DI(2) => W_49_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_49_31_i_8_n_0,
   S(1) => W_49_31_i_7_n_0,
   S(2) => W_49_31_i_6_n_0,
   S(3) => W_49_31_i_5_n_0,
   CO(0) => W_reg_49_31_i_1_n_3,
   CO(1) => W_reg_49_31_i_1_n_2,
   CO(2) => W_reg_49_31_i_1_n_1,
   CO(3) => NLW_W_reg_49_31_i_1_CO_UNCONNECTED_3,
   O(0) => x41_out_28,
   O(1) => x41_out_29,
   O(2) => x41_out_30,
   O(3) => x41_out_31
);
W_reg_49_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x41_out_3,
   R => '0',
   Q => W_reg_49_3
);
W_reg_49_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_49_3_i_5_n_0,
   DI(1) => W_49_3_i_4_n_0,
   DI(2) => W_49_3_i_3_n_0,
   DI(3) => W_49_3_i_2_n_0,
   S(0) => W_49_3_i_9_n_0,
   S(1) => W_49_3_i_8_n_0,
   S(2) => W_49_3_i_7_n_0,
   S(3) => W_49_3_i_6_n_0,
   CO(0) => W_reg_49_3_i_1_n_3,
   CO(1) => W_reg_49_3_i_1_n_2,
   CO(2) => W_reg_49_3_i_1_n_1,
   CO(3) => W_reg_49_3_i_1_n_0,
   O(0) => x41_out_0,
   O(1) => x41_out_1,
   O(2) => x41_out_2,
   O(3) => x41_out_3
);
W_reg_49_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x41_out_4,
   R => '0',
   Q => W_reg_49_4
);
W_reg_49_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x41_out_5,
   R => '0',
   Q => W_reg_49_5
);
W_reg_49_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x41_out_6,
   R => '0',
   Q => W_reg_49_6
);
W_reg_49_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x41_out_7,
   R => '0',
   Q => W_reg_49_7
);
W_reg_49_7_i_1 : CARRY4
 port map (
   CI => W_reg_49_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_49_7_i_5_n_0,
   DI(1) => W_49_7_i_4_n_0,
   DI(2) => W_49_7_i_3_n_0,
   DI(3) => W_49_7_i_2_n_0,
   S(0) => W_49_7_i_9_n_0,
   S(1) => W_49_7_i_8_n_0,
   S(2) => W_49_7_i_7_n_0,
   S(3) => W_49_7_i_6_n_0,
   CO(0) => W_reg_49_7_i_1_n_3,
   CO(1) => W_reg_49_7_i_1_n_2,
   CO(2) => W_reg_49_7_i_1_n_1,
   CO(3) => W_reg_49_7_i_1_n_0,
   O(0) => x41_out_4,
   O(1) => x41_out_5,
   O(2) => x41_out_6,
   O(3) => x41_out_7
);
W_reg_49_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x41_out_8,
   R => '0',
   Q => W_reg_49_8
);
W_reg_49_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x41_out_9,
   R => '0',
   Q => W_reg_49_9
);
W_reg_4_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_4_0,
   R => '0',
   Q => W_reg_4_0
);
W_reg_4_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_4_10,
   R => '0',
   Q => W_reg_4_10
);
W_reg_4_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_4_11,
   R => '0',
   Q => W_reg_4_11
);
W_reg_4_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_4_12,
   R => '0',
   Q => W_reg_4_12
);
W_reg_4_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_4_13,
   R => '0',
   Q => W_reg_4_13
);
W_reg_4_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_4_14,
   R => '0',
   Q => W_reg_4_14
);
W_reg_4_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_4_15,
   R => '0',
   Q => W_reg_4_15
);
W_reg_4_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_4_16,
   R => '0',
   Q => W_reg_4_16
);
W_reg_4_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_4_17,
   R => '0',
   Q => W_reg_4_17
);
W_reg_4_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_4_18,
   R => '0',
   Q => W_reg_4_18
);
W_reg_4_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_4_19,
   R => '0',
   Q => W_reg_4_19
);
W_reg_4_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_4_1,
   R => '0',
   Q => W_reg_4_1
);
W_reg_4_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_4_20,
   R => '0',
   Q => W_reg_4_20
);
W_reg_4_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_4_21,
   R => '0',
   Q => W_reg_4_21
);
W_reg_4_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_4_22,
   R => '0',
   Q => W_reg_4_22
);
W_reg_4_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_4_23,
   R => '0',
   Q => W_reg_4_23
);
W_reg_4_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_4_24,
   R => '0',
   Q => W_reg_4_24
);
W_reg_4_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_4_25,
   R => '0',
   Q => W_reg_4_25
);
W_reg_4_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_4_26,
   R => '0',
   Q => W_reg_4_26
);
W_reg_4_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_4_27,
   R => '0',
   Q => W_reg_4_27
);
W_reg_4_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_4_28,
   R => '0',
   Q => W_reg_4_28
);
W_reg_4_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_4_29,
   R => '0',
   Q => W_reg_4_29
);
W_reg_4_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_4_2,
   R => '0',
   Q => W_reg_4_2
);
W_reg_4_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_4_30,
   R => '0',
   Q => W_reg_4_30
);
W_reg_4_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_4_31,
   R => '0',
   Q => W_reg_4_31
);
W_reg_4_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_4_3,
   R => '0',
   Q => W_reg_4_3
);
W_reg_4_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_4_4,
   R => '0',
   Q => W_reg_4_4
);
W_reg_4_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_4_5,
   R => '0',
   Q => W_reg_4_5
);
W_reg_4_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_4_6,
   R => '0',
   Q => W_reg_4_6
);
W_reg_4_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_4_7,
   R => '0',
   Q => W_reg_4_7
);
W_reg_4_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_4_8,
   R => '0',
   Q => W_reg_4_8
);
W_reg_4_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_4_9,
   R => '0',
   Q => W_reg_4_9
);
W_reg_50_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x38_out_0,
   R => '0',
   Q => W_reg_50_0
);
W_reg_50_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x38_out_10,
   R => '0',
   Q => W_reg_50_10
);
W_reg_50_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x38_out_11,
   R => '0',
   Q => W_reg_50_11
);
W_reg_50_11_i_1 : CARRY4
 port map (
   CI => W_reg_50_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_50_11_i_5_n_0,
   DI(1) => W_50_11_i_4_n_0,
   DI(2) => W_50_11_i_3_n_0,
   DI(3) => W_50_11_i_2_n_0,
   S(0) => W_50_11_i_9_n_0,
   S(1) => W_50_11_i_8_n_0,
   S(2) => W_50_11_i_7_n_0,
   S(3) => W_50_11_i_6_n_0,
   CO(0) => W_reg_50_11_i_1_n_3,
   CO(1) => W_reg_50_11_i_1_n_2,
   CO(2) => W_reg_50_11_i_1_n_1,
   CO(3) => W_reg_50_11_i_1_n_0,
   O(0) => x38_out_8,
   O(1) => x38_out_9,
   O(2) => x38_out_10,
   O(3) => x38_out_11
);
W_reg_50_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x38_out_12,
   R => '0',
   Q => W_reg_50_12
);
W_reg_50_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x38_out_13,
   R => '0',
   Q => W_reg_50_13
);
W_reg_50_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x38_out_14,
   R => '0',
   Q => W_reg_50_14
);
W_reg_50_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x38_out_15,
   R => '0',
   Q => W_reg_50_15
);
W_reg_50_15_i_1 : CARRY4
 port map (
   CI => W_reg_50_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_50_15_i_5_n_0,
   DI(1) => W_50_15_i_4_n_0,
   DI(2) => W_50_15_i_3_n_0,
   DI(3) => W_50_15_i_2_n_0,
   S(0) => W_50_15_i_9_n_0,
   S(1) => W_50_15_i_8_n_0,
   S(2) => W_50_15_i_7_n_0,
   S(3) => W_50_15_i_6_n_0,
   CO(0) => W_reg_50_15_i_1_n_3,
   CO(1) => W_reg_50_15_i_1_n_2,
   CO(2) => W_reg_50_15_i_1_n_1,
   CO(3) => W_reg_50_15_i_1_n_0,
   O(0) => x38_out_12,
   O(1) => x38_out_13,
   O(2) => x38_out_14,
   O(3) => x38_out_15
);
W_reg_50_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x38_out_16,
   R => '0',
   Q => W_reg_50_16
);
W_reg_50_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x38_out_17,
   R => '0',
   Q => W_reg_50_17
);
W_reg_50_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x38_out_18,
   R => '0',
   Q => W_reg_50_18
);
W_reg_50_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x38_out_19,
   R => '0',
   Q => W_reg_50_19
);
W_reg_50_19_i_1 : CARRY4
 port map (
   CI => W_reg_50_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_50_19_i_5_n_0,
   DI(1) => W_50_19_i_4_n_0,
   DI(2) => W_50_19_i_3_n_0,
   DI(3) => W_50_19_i_2_n_0,
   S(0) => W_50_19_i_9_n_0,
   S(1) => W_50_19_i_8_n_0,
   S(2) => W_50_19_i_7_n_0,
   S(3) => W_50_19_i_6_n_0,
   CO(0) => W_reg_50_19_i_1_n_3,
   CO(1) => W_reg_50_19_i_1_n_2,
   CO(2) => W_reg_50_19_i_1_n_1,
   CO(3) => W_reg_50_19_i_1_n_0,
   O(0) => x38_out_16,
   O(1) => x38_out_17,
   O(2) => x38_out_18,
   O(3) => x38_out_19
);
W_reg_50_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x38_out_1,
   R => '0',
   Q => W_reg_50_1
);
W_reg_50_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x38_out_20,
   R => '0',
   Q => W_reg_50_20
);
W_reg_50_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x38_out_21,
   R => '0',
   Q => W_reg_50_21
);
W_reg_50_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x38_out_22,
   R => '0',
   Q => W_reg_50_22
);
W_reg_50_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x38_out_23,
   R => '0',
   Q => W_reg_50_23
);
W_reg_50_23_i_1 : CARRY4
 port map (
   CI => W_reg_50_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_50_23_i_5_n_0,
   DI(1) => W_50_23_i_4_n_0,
   DI(2) => W_50_23_i_3_n_0,
   DI(3) => W_50_23_i_2_n_0,
   S(0) => W_50_23_i_9_n_0,
   S(1) => W_50_23_i_8_n_0,
   S(2) => W_50_23_i_7_n_0,
   S(3) => W_50_23_i_6_n_0,
   CO(0) => W_reg_50_23_i_1_n_3,
   CO(1) => W_reg_50_23_i_1_n_2,
   CO(2) => W_reg_50_23_i_1_n_1,
   CO(3) => W_reg_50_23_i_1_n_0,
   O(0) => x38_out_20,
   O(1) => x38_out_21,
   O(2) => x38_out_22,
   O(3) => x38_out_23
);
W_reg_50_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x38_out_24,
   R => '0',
   Q => W_reg_50_24
);
W_reg_50_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x38_out_25,
   R => '0',
   Q => W_reg_50_25
);
W_reg_50_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x38_out_26,
   R => '0',
   Q => W_reg_50_26
);
W_reg_50_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x38_out_27,
   R => '0',
   Q => W_reg_50_27
);
W_reg_50_27_i_1 : CARRY4
 port map (
   CI => W_reg_50_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_50_27_i_5_n_0,
   DI(1) => W_50_27_i_4_n_0,
   DI(2) => W_50_27_i_3_n_0,
   DI(3) => W_50_27_i_2_n_0,
   S(0) => W_50_27_i_9_n_0,
   S(1) => W_50_27_i_8_n_0,
   S(2) => W_50_27_i_7_n_0,
   S(3) => W_50_27_i_6_n_0,
   CO(0) => W_reg_50_27_i_1_n_3,
   CO(1) => W_reg_50_27_i_1_n_2,
   CO(2) => W_reg_50_27_i_1_n_1,
   CO(3) => W_reg_50_27_i_1_n_0,
   O(0) => x38_out_24,
   O(1) => x38_out_25,
   O(2) => x38_out_26,
   O(3) => x38_out_27
);
W_reg_50_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x38_out_28,
   R => '0',
   Q => W_reg_50_28
);
W_reg_50_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x38_out_29,
   R => '0',
   Q => W_reg_50_29
);
W_reg_50_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x38_out_2,
   R => '0',
   Q => W_reg_50_2
);
W_reg_50_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x38_out_30,
   R => '0',
   Q => W_reg_50_30
);
W_reg_50_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x38_out_31,
   R => '0',
   Q => W_reg_50_31
);
W_reg_50_31_i_1 : CARRY4
 port map (
   CI => W_reg_50_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_50_31_i_4_n_0,
   DI(1) => W_50_31_i_3_n_0,
   DI(2) => W_50_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_50_31_i_8_n_0,
   S(1) => W_50_31_i_7_n_0,
   S(2) => W_50_31_i_6_n_0,
   S(3) => W_50_31_i_5_n_0,
   CO(0) => W_reg_50_31_i_1_n_3,
   CO(1) => W_reg_50_31_i_1_n_2,
   CO(2) => W_reg_50_31_i_1_n_1,
   CO(3) => NLW_W_reg_50_31_i_1_CO_UNCONNECTED_3,
   O(0) => x38_out_28,
   O(1) => x38_out_29,
   O(2) => x38_out_30,
   O(3) => x38_out_31
);
W_reg_50_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x38_out_3,
   R => '0',
   Q => W_reg_50_3
);
W_reg_50_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_50_3_i_5_n_0,
   DI(1) => W_50_3_i_4_n_0,
   DI(2) => W_50_3_i_3_n_0,
   DI(3) => W_50_3_i_2_n_0,
   S(0) => W_50_3_i_9_n_0,
   S(1) => W_50_3_i_8_n_0,
   S(2) => W_50_3_i_7_n_0,
   S(3) => W_50_3_i_6_n_0,
   CO(0) => W_reg_50_3_i_1_n_3,
   CO(1) => W_reg_50_3_i_1_n_2,
   CO(2) => W_reg_50_3_i_1_n_1,
   CO(3) => W_reg_50_3_i_1_n_0,
   O(0) => x38_out_0,
   O(1) => x38_out_1,
   O(2) => x38_out_2,
   O(3) => x38_out_3
);
W_reg_50_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x38_out_4,
   R => '0',
   Q => W_reg_50_4
);
W_reg_50_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x38_out_5,
   R => '0',
   Q => W_reg_50_5
);
W_reg_50_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x38_out_6,
   R => '0',
   Q => W_reg_50_6
);
W_reg_50_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x38_out_7,
   R => '0',
   Q => W_reg_50_7
);
W_reg_50_7_i_1 : CARRY4
 port map (
   CI => W_reg_50_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_50_7_i_5_n_0,
   DI(1) => W_50_7_i_4_n_0,
   DI(2) => W_50_7_i_3_n_0,
   DI(3) => W_50_7_i_2_n_0,
   S(0) => W_50_7_i_9_n_0,
   S(1) => W_50_7_i_8_n_0,
   S(2) => W_50_7_i_7_n_0,
   S(3) => W_50_7_i_6_n_0,
   CO(0) => W_reg_50_7_i_1_n_3,
   CO(1) => W_reg_50_7_i_1_n_2,
   CO(2) => W_reg_50_7_i_1_n_1,
   CO(3) => W_reg_50_7_i_1_n_0,
   O(0) => x38_out_4,
   O(1) => x38_out_5,
   O(2) => x38_out_6,
   O(3) => x38_out_7
);
W_reg_50_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x38_out_8,
   R => '0',
   Q => W_reg_50_8
);
W_reg_50_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x38_out_9,
   R => '0',
   Q => W_reg_50_9
);
W_reg_51_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x35_out_0,
   R => '0',
   Q => W_reg_51_0
);
W_reg_51_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x35_out_10,
   R => '0',
   Q => W_reg_51_10
);
W_reg_51_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x35_out_11,
   R => '0',
   Q => W_reg_51_11
);
W_reg_51_11_i_1 : CARRY4
 port map (
   CI => W_reg_51_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_51_11_i_5_n_0,
   DI(1) => W_51_11_i_4_n_0,
   DI(2) => W_51_11_i_3_n_0,
   DI(3) => W_51_11_i_2_n_0,
   S(0) => W_51_11_i_9_n_0,
   S(1) => W_51_11_i_8_n_0,
   S(2) => W_51_11_i_7_n_0,
   S(3) => W_51_11_i_6_n_0,
   CO(0) => W_reg_51_11_i_1_n_3,
   CO(1) => W_reg_51_11_i_1_n_2,
   CO(2) => W_reg_51_11_i_1_n_1,
   CO(3) => W_reg_51_11_i_1_n_0,
   O(0) => x35_out_8,
   O(1) => x35_out_9,
   O(2) => x35_out_10,
   O(3) => x35_out_11
);
W_reg_51_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x35_out_12,
   R => '0',
   Q => W_reg_51_12
);
W_reg_51_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x35_out_13,
   R => '0',
   Q => W_reg_51_13
);
W_reg_51_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x35_out_14,
   R => '0',
   Q => W_reg_51_14
);
W_reg_51_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x35_out_15,
   R => '0',
   Q => W_reg_51_15
);
W_reg_51_15_i_1 : CARRY4
 port map (
   CI => W_reg_51_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_51_15_i_5_n_0,
   DI(1) => W_51_15_i_4_n_0,
   DI(2) => W_51_15_i_3_n_0,
   DI(3) => W_51_15_i_2_n_0,
   S(0) => W_51_15_i_9_n_0,
   S(1) => W_51_15_i_8_n_0,
   S(2) => W_51_15_i_7_n_0,
   S(3) => W_51_15_i_6_n_0,
   CO(0) => W_reg_51_15_i_1_n_3,
   CO(1) => W_reg_51_15_i_1_n_2,
   CO(2) => W_reg_51_15_i_1_n_1,
   CO(3) => W_reg_51_15_i_1_n_0,
   O(0) => x35_out_12,
   O(1) => x35_out_13,
   O(2) => x35_out_14,
   O(3) => x35_out_15
);
W_reg_51_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x35_out_16,
   R => '0',
   Q => W_reg_51_16
);
W_reg_51_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x35_out_17,
   R => '0',
   Q => W_reg_51_17
);
W_reg_51_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x35_out_18,
   R => '0',
   Q => W_reg_51_18
);
W_reg_51_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x35_out_19,
   R => '0',
   Q => W_reg_51_19
);
W_reg_51_19_i_1 : CARRY4
 port map (
   CI => W_reg_51_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_51_19_i_5_n_0,
   DI(1) => W_51_19_i_4_n_0,
   DI(2) => W_51_19_i_3_n_0,
   DI(3) => W_51_19_i_2_n_0,
   S(0) => W_51_19_i_9_n_0,
   S(1) => W_51_19_i_8_n_0,
   S(2) => W_51_19_i_7_n_0,
   S(3) => W_51_19_i_6_n_0,
   CO(0) => W_reg_51_19_i_1_n_3,
   CO(1) => W_reg_51_19_i_1_n_2,
   CO(2) => W_reg_51_19_i_1_n_1,
   CO(3) => W_reg_51_19_i_1_n_0,
   O(0) => x35_out_16,
   O(1) => x35_out_17,
   O(2) => x35_out_18,
   O(3) => x35_out_19
);
W_reg_51_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x35_out_1,
   R => '0',
   Q => W_reg_51_1
);
W_reg_51_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x35_out_20,
   R => '0',
   Q => W_reg_51_20
);
W_reg_51_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x35_out_21,
   R => '0',
   Q => W_reg_51_21
);
W_reg_51_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x35_out_22,
   R => '0',
   Q => W_reg_51_22
);
W_reg_51_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x35_out_23,
   R => '0',
   Q => W_reg_51_23
);
W_reg_51_23_i_1 : CARRY4
 port map (
   CI => W_reg_51_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_51_23_i_5_n_0,
   DI(1) => W_51_23_i_4_n_0,
   DI(2) => W_51_23_i_3_n_0,
   DI(3) => W_51_23_i_2_n_0,
   S(0) => W_51_23_i_9_n_0,
   S(1) => W_51_23_i_8_n_0,
   S(2) => W_51_23_i_7_n_0,
   S(3) => W_51_23_i_6_n_0,
   CO(0) => W_reg_51_23_i_1_n_3,
   CO(1) => W_reg_51_23_i_1_n_2,
   CO(2) => W_reg_51_23_i_1_n_1,
   CO(3) => W_reg_51_23_i_1_n_0,
   O(0) => x35_out_20,
   O(1) => x35_out_21,
   O(2) => x35_out_22,
   O(3) => x35_out_23
);
W_reg_51_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x35_out_24,
   R => '0',
   Q => W_reg_51_24
);
W_reg_51_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x35_out_25,
   R => '0',
   Q => W_reg_51_25
);
W_reg_51_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x35_out_26,
   R => '0',
   Q => W_reg_51_26
);
W_reg_51_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x35_out_27,
   R => '0',
   Q => W_reg_51_27
);
W_reg_51_27_i_1 : CARRY4
 port map (
   CI => W_reg_51_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_51_27_i_5_n_0,
   DI(1) => W_51_27_i_4_n_0,
   DI(2) => W_51_27_i_3_n_0,
   DI(3) => W_51_27_i_2_n_0,
   S(0) => W_51_27_i_9_n_0,
   S(1) => W_51_27_i_8_n_0,
   S(2) => W_51_27_i_7_n_0,
   S(3) => W_51_27_i_6_n_0,
   CO(0) => W_reg_51_27_i_1_n_3,
   CO(1) => W_reg_51_27_i_1_n_2,
   CO(2) => W_reg_51_27_i_1_n_1,
   CO(3) => W_reg_51_27_i_1_n_0,
   O(0) => x35_out_24,
   O(1) => x35_out_25,
   O(2) => x35_out_26,
   O(3) => x35_out_27
);
W_reg_51_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x35_out_28,
   R => '0',
   Q => W_reg_51_28
);
W_reg_51_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x35_out_29,
   R => '0',
   Q => W_reg_51_29
);
W_reg_51_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x35_out_2,
   R => '0',
   Q => W_reg_51_2
);
W_reg_51_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x35_out_30,
   R => '0',
   Q => W_reg_51_30
);
W_reg_51_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x35_out_31,
   R => '0',
   Q => W_reg_51_31
);
W_reg_51_31_i_1 : CARRY4
 port map (
   CI => W_reg_51_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_51_31_i_4_n_0,
   DI(1) => W_51_31_i_3_n_0,
   DI(2) => W_51_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_51_31_i_8_n_0,
   S(1) => W_51_31_i_7_n_0,
   S(2) => W_51_31_i_6_n_0,
   S(3) => W_51_31_i_5_n_0,
   CO(0) => W_reg_51_31_i_1_n_3,
   CO(1) => W_reg_51_31_i_1_n_2,
   CO(2) => W_reg_51_31_i_1_n_1,
   CO(3) => NLW_W_reg_51_31_i_1_CO_UNCONNECTED_3,
   O(0) => x35_out_28,
   O(1) => x35_out_29,
   O(2) => x35_out_30,
   O(3) => x35_out_31
);
W_reg_51_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x35_out_3,
   R => '0',
   Q => W_reg_51_3
);
W_reg_51_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_51_3_i_5_n_0,
   DI(1) => W_51_3_i_4_n_0,
   DI(2) => W_51_3_i_3_n_0,
   DI(3) => W_51_3_i_2_n_0,
   S(0) => W_51_3_i_9_n_0,
   S(1) => W_51_3_i_8_n_0,
   S(2) => W_51_3_i_7_n_0,
   S(3) => W_51_3_i_6_n_0,
   CO(0) => W_reg_51_3_i_1_n_3,
   CO(1) => W_reg_51_3_i_1_n_2,
   CO(2) => W_reg_51_3_i_1_n_1,
   CO(3) => W_reg_51_3_i_1_n_0,
   O(0) => x35_out_0,
   O(1) => x35_out_1,
   O(2) => x35_out_2,
   O(3) => x35_out_3
);
W_reg_51_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x35_out_4,
   R => '0',
   Q => W_reg_51_4
);
W_reg_51_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x35_out_5,
   R => '0',
   Q => W_reg_51_5
);
W_reg_51_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x35_out_6,
   R => '0',
   Q => W_reg_51_6
);
W_reg_51_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x35_out_7,
   R => '0',
   Q => W_reg_51_7
);
W_reg_51_7_i_1 : CARRY4
 port map (
   CI => W_reg_51_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_51_7_i_5_n_0,
   DI(1) => W_51_7_i_4_n_0,
   DI(2) => W_51_7_i_3_n_0,
   DI(3) => W_51_7_i_2_n_0,
   S(0) => W_51_7_i_9_n_0,
   S(1) => W_51_7_i_8_n_0,
   S(2) => W_51_7_i_7_n_0,
   S(3) => W_51_7_i_6_n_0,
   CO(0) => W_reg_51_7_i_1_n_3,
   CO(1) => W_reg_51_7_i_1_n_2,
   CO(2) => W_reg_51_7_i_1_n_1,
   CO(3) => W_reg_51_7_i_1_n_0,
   O(0) => x35_out_4,
   O(1) => x35_out_5,
   O(2) => x35_out_6,
   O(3) => x35_out_7
);
W_reg_51_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x35_out_8,
   R => '0',
   Q => W_reg_51_8
);
W_reg_51_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x35_out_9,
   R => '0',
   Q => W_reg_51_9
);
W_reg_52_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x32_out_0,
   R => '0',
   Q => W_reg_52_0
);
W_reg_52_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x32_out_10,
   R => '0',
   Q => W_reg_52_10
);
W_reg_52_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x32_out_11,
   R => '0',
   Q => W_reg_52_11
);
W_reg_52_11_i_1 : CARRY4
 port map (
   CI => W_reg_52_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_52_11_i_5_n_0,
   DI(1) => W_52_11_i_4_n_0,
   DI(2) => W_52_11_i_3_n_0,
   DI(3) => W_52_11_i_2_n_0,
   S(0) => W_52_11_i_9_n_0,
   S(1) => W_52_11_i_8_n_0,
   S(2) => W_52_11_i_7_n_0,
   S(3) => W_52_11_i_6_n_0,
   CO(0) => W_reg_52_11_i_1_n_3,
   CO(1) => W_reg_52_11_i_1_n_2,
   CO(2) => W_reg_52_11_i_1_n_1,
   CO(3) => W_reg_52_11_i_1_n_0,
   O(0) => x32_out_8,
   O(1) => x32_out_9,
   O(2) => x32_out_10,
   O(3) => x32_out_11
);
W_reg_52_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x32_out_12,
   R => '0',
   Q => W_reg_52_12
);
W_reg_52_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x32_out_13,
   R => '0',
   Q => W_reg_52_13
);
W_reg_52_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x32_out_14,
   R => '0',
   Q => W_reg_52_14
);
W_reg_52_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x32_out_15,
   R => '0',
   Q => W_reg_52_15
);
W_reg_52_15_i_1 : CARRY4
 port map (
   CI => W_reg_52_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_52_15_i_5_n_0,
   DI(1) => W_52_15_i_4_n_0,
   DI(2) => W_52_15_i_3_n_0,
   DI(3) => W_52_15_i_2_n_0,
   S(0) => W_52_15_i_9_n_0,
   S(1) => W_52_15_i_8_n_0,
   S(2) => W_52_15_i_7_n_0,
   S(3) => W_52_15_i_6_n_0,
   CO(0) => W_reg_52_15_i_1_n_3,
   CO(1) => W_reg_52_15_i_1_n_2,
   CO(2) => W_reg_52_15_i_1_n_1,
   CO(3) => W_reg_52_15_i_1_n_0,
   O(0) => x32_out_12,
   O(1) => x32_out_13,
   O(2) => x32_out_14,
   O(3) => x32_out_15
);
W_reg_52_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x32_out_16,
   R => '0',
   Q => W_reg_52_16
);
W_reg_52_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x32_out_17,
   R => '0',
   Q => W_reg_52_17
);
W_reg_52_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x32_out_18,
   R => '0',
   Q => W_reg_52_18
);
W_reg_52_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x32_out_19,
   R => '0',
   Q => W_reg_52_19
);
W_reg_52_19_i_1 : CARRY4
 port map (
   CI => W_reg_52_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_52_19_i_5_n_0,
   DI(1) => W_52_19_i_4_n_0,
   DI(2) => W_52_19_i_3_n_0,
   DI(3) => W_52_19_i_2_n_0,
   S(0) => W_52_19_i_9_n_0,
   S(1) => W_52_19_i_8_n_0,
   S(2) => W_52_19_i_7_n_0,
   S(3) => W_52_19_i_6_n_0,
   CO(0) => W_reg_52_19_i_1_n_3,
   CO(1) => W_reg_52_19_i_1_n_2,
   CO(2) => W_reg_52_19_i_1_n_1,
   CO(3) => W_reg_52_19_i_1_n_0,
   O(0) => x32_out_16,
   O(1) => x32_out_17,
   O(2) => x32_out_18,
   O(3) => x32_out_19
);
W_reg_52_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x32_out_1,
   R => '0',
   Q => W_reg_52_1
);
W_reg_52_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x32_out_20,
   R => '0',
   Q => W_reg_52_20
);
W_reg_52_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x32_out_21,
   R => '0',
   Q => W_reg_52_21
);
W_reg_52_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x32_out_22,
   R => '0',
   Q => W_reg_52_22
);
W_reg_52_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x32_out_23,
   R => '0',
   Q => W_reg_52_23
);
W_reg_52_23_i_1 : CARRY4
 port map (
   CI => W_reg_52_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_52_23_i_5_n_0,
   DI(1) => W_52_23_i_4_n_0,
   DI(2) => W_52_23_i_3_n_0,
   DI(3) => W_52_23_i_2_n_0,
   S(0) => W_52_23_i_9_n_0,
   S(1) => W_52_23_i_8_n_0,
   S(2) => W_52_23_i_7_n_0,
   S(3) => W_52_23_i_6_n_0,
   CO(0) => W_reg_52_23_i_1_n_3,
   CO(1) => W_reg_52_23_i_1_n_2,
   CO(2) => W_reg_52_23_i_1_n_1,
   CO(3) => W_reg_52_23_i_1_n_0,
   O(0) => x32_out_20,
   O(1) => x32_out_21,
   O(2) => x32_out_22,
   O(3) => x32_out_23
);
W_reg_52_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x32_out_24,
   R => '0',
   Q => W_reg_52_24
);
W_reg_52_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x32_out_25,
   R => '0',
   Q => W_reg_52_25
);
W_reg_52_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x32_out_26,
   R => '0',
   Q => W_reg_52_26
);
W_reg_52_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x32_out_27,
   R => '0',
   Q => W_reg_52_27
);
W_reg_52_27_i_1 : CARRY4
 port map (
   CI => W_reg_52_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_52_27_i_5_n_0,
   DI(1) => W_52_27_i_4_n_0,
   DI(2) => W_52_27_i_3_n_0,
   DI(3) => W_52_27_i_2_n_0,
   S(0) => W_52_27_i_9_n_0,
   S(1) => W_52_27_i_8_n_0,
   S(2) => W_52_27_i_7_n_0,
   S(3) => W_52_27_i_6_n_0,
   CO(0) => W_reg_52_27_i_1_n_3,
   CO(1) => W_reg_52_27_i_1_n_2,
   CO(2) => W_reg_52_27_i_1_n_1,
   CO(3) => W_reg_52_27_i_1_n_0,
   O(0) => x32_out_24,
   O(1) => x32_out_25,
   O(2) => x32_out_26,
   O(3) => x32_out_27
);
W_reg_52_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x32_out_28,
   R => '0',
   Q => W_reg_52_28
);
W_reg_52_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x32_out_29,
   R => '0',
   Q => W_reg_52_29
);
W_reg_52_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x32_out_2,
   R => '0',
   Q => W_reg_52_2
);
W_reg_52_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x32_out_30,
   R => '0',
   Q => W_reg_52_30
);
W_reg_52_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x32_out_31,
   R => '0',
   Q => W_reg_52_31
);
W_reg_52_31_i_1 : CARRY4
 port map (
   CI => W_reg_52_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_52_31_i_4_n_0,
   DI(1) => W_52_31_i_3_n_0,
   DI(2) => W_52_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_52_31_i_8_n_0,
   S(1) => W_52_31_i_7_n_0,
   S(2) => W_52_31_i_6_n_0,
   S(3) => W_52_31_i_5_n_0,
   CO(0) => W_reg_52_31_i_1_n_3,
   CO(1) => W_reg_52_31_i_1_n_2,
   CO(2) => W_reg_52_31_i_1_n_1,
   CO(3) => NLW_W_reg_52_31_i_1_CO_UNCONNECTED_3,
   O(0) => x32_out_28,
   O(1) => x32_out_29,
   O(2) => x32_out_30,
   O(3) => x32_out_31
);
W_reg_52_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x32_out_3,
   R => '0',
   Q => W_reg_52_3
);
W_reg_52_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_52_3_i_5_n_0,
   DI(1) => W_52_3_i_4_n_0,
   DI(2) => W_52_3_i_3_n_0,
   DI(3) => W_52_3_i_2_n_0,
   S(0) => W_52_3_i_9_n_0,
   S(1) => W_52_3_i_8_n_0,
   S(2) => W_52_3_i_7_n_0,
   S(3) => W_52_3_i_6_n_0,
   CO(0) => W_reg_52_3_i_1_n_3,
   CO(1) => W_reg_52_3_i_1_n_2,
   CO(2) => W_reg_52_3_i_1_n_1,
   CO(3) => W_reg_52_3_i_1_n_0,
   O(0) => x32_out_0,
   O(1) => x32_out_1,
   O(2) => x32_out_2,
   O(3) => x32_out_3
);
W_reg_52_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x32_out_4,
   R => '0',
   Q => W_reg_52_4
);
W_reg_52_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x32_out_5,
   R => '0',
   Q => W_reg_52_5
);
W_reg_52_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x32_out_6,
   R => '0',
   Q => W_reg_52_6
);
W_reg_52_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x32_out_7,
   R => '0',
   Q => W_reg_52_7
);
W_reg_52_7_i_1 : CARRY4
 port map (
   CI => W_reg_52_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_52_7_i_5_n_0,
   DI(1) => W_52_7_i_4_n_0,
   DI(2) => W_52_7_i_3_n_0,
   DI(3) => W_52_7_i_2_n_0,
   S(0) => W_52_7_i_9_n_0,
   S(1) => W_52_7_i_8_n_0,
   S(2) => W_52_7_i_7_n_0,
   S(3) => W_52_7_i_6_n_0,
   CO(0) => W_reg_52_7_i_1_n_3,
   CO(1) => W_reg_52_7_i_1_n_2,
   CO(2) => W_reg_52_7_i_1_n_1,
   CO(3) => W_reg_52_7_i_1_n_0,
   O(0) => x32_out_4,
   O(1) => x32_out_5,
   O(2) => x32_out_6,
   O(3) => x32_out_7
);
W_reg_52_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x32_out_8,
   R => '0',
   Q => W_reg_52_8
);
W_reg_52_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x32_out_9,
   R => '0',
   Q => W_reg_52_9
);
W_reg_53_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x29_out_0,
   R => '0',
   Q => W_reg_53_0
);
W_reg_53_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x29_out_10,
   R => '0',
   Q => W_reg_53_10
);
W_reg_53_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x29_out_11,
   R => '0',
   Q => W_reg_53_11
);
W_reg_53_11_i_1 : CARRY4
 port map (
   CI => W_reg_53_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_53_11_i_5_n_0,
   DI(1) => W_53_11_i_4_n_0,
   DI(2) => W_53_11_i_3_n_0,
   DI(3) => W_53_11_i_2_n_0,
   S(0) => W_53_11_i_9_n_0,
   S(1) => W_53_11_i_8_n_0,
   S(2) => W_53_11_i_7_n_0,
   S(3) => W_53_11_i_6_n_0,
   CO(0) => W_reg_53_11_i_1_n_3,
   CO(1) => W_reg_53_11_i_1_n_2,
   CO(2) => W_reg_53_11_i_1_n_1,
   CO(3) => W_reg_53_11_i_1_n_0,
   O(0) => x29_out_8,
   O(1) => x29_out_9,
   O(2) => x29_out_10,
   O(3) => x29_out_11
);
W_reg_53_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x29_out_12,
   R => '0',
   Q => W_reg_53_12
);
W_reg_53_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x29_out_13,
   R => '0',
   Q => W_reg_53_13
);
W_reg_53_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x29_out_14,
   R => '0',
   Q => W_reg_53_14
);
W_reg_53_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x29_out_15,
   R => '0',
   Q => W_reg_53_15
);
W_reg_53_15_i_1 : CARRY4
 port map (
   CI => W_reg_53_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_53_15_i_5_n_0,
   DI(1) => W_53_15_i_4_n_0,
   DI(2) => W_53_15_i_3_n_0,
   DI(3) => W_53_15_i_2_n_0,
   S(0) => W_53_15_i_9_n_0,
   S(1) => W_53_15_i_8_n_0,
   S(2) => W_53_15_i_7_n_0,
   S(3) => W_53_15_i_6_n_0,
   CO(0) => W_reg_53_15_i_1_n_3,
   CO(1) => W_reg_53_15_i_1_n_2,
   CO(2) => W_reg_53_15_i_1_n_1,
   CO(3) => W_reg_53_15_i_1_n_0,
   O(0) => x29_out_12,
   O(1) => x29_out_13,
   O(2) => x29_out_14,
   O(3) => x29_out_15
);
W_reg_53_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x29_out_16,
   R => '0',
   Q => W_reg_53_16
);
W_reg_53_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x29_out_17,
   R => '0',
   Q => W_reg_53_17
);
W_reg_53_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x29_out_18,
   R => '0',
   Q => W_reg_53_18
);
W_reg_53_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x29_out_19,
   R => '0',
   Q => W_reg_53_19
);
W_reg_53_19_i_1 : CARRY4
 port map (
   CI => W_reg_53_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_53_19_i_5_n_0,
   DI(1) => W_53_19_i_4_n_0,
   DI(2) => W_53_19_i_3_n_0,
   DI(3) => W_53_19_i_2_n_0,
   S(0) => W_53_19_i_9_n_0,
   S(1) => W_53_19_i_8_n_0,
   S(2) => W_53_19_i_7_n_0,
   S(3) => W_53_19_i_6_n_0,
   CO(0) => W_reg_53_19_i_1_n_3,
   CO(1) => W_reg_53_19_i_1_n_2,
   CO(2) => W_reg_53_19_i_1_n_1,
   CO(3) => W_reg_53_19_i_1_n_0,
   O(0) => x29_out_16,
   O(1) => x29_out_17,
   O(2) => x29_out_18,
   O(3) => x29_out_19
);
W_reg_53_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x29_out_1,
   R => '0',
   Q => W_reg_53_1
);
W_reg_53_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x29_out_20,
   R => '0',
   Q => W_reg_53_20
);
W_reg_53_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x29_out_21,
   R => '0',
   Q => W_reg_53_21
);
W_reg_53_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x29_out_22,
   R => '0',
   Q => W_reg_53_22
);
W_reg_53_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x29_out_23,
   R => '0',
   Q => W_reg_53_23
);
W_reg_53_23_i_1 : CARRY4
 port map (
   CI => W_reg_53_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_53_23_i_5_n_0,
   DI(1) => W_53_23_i_4_n_0,
   DI(2) => W_53_23_i_3_n_0,
   DI(3) => W_53_23_i_2_n_0,
   S(0) => W_53_23_i_9_n_0,
   S(1) => W_53_23_i_8_n_0,
   S(2) => W_53_23_i_7_n_0,
   S(3) => W_53_23_i_6_n_0,
   CO(0) => W_reg_53_23_i_1_n_3,
   CO(1) => W_reg_53_23_i_1_n_2,
   CO(2) => W_reg_53_23_i_1_n_1,
   CO(3) => W_reg_53_23_i_1_n_0,
   O(0) => x29_out_20,
   O(1) => x29_out_21,
   O(2) => x29_out_22,
   O(3) => x29_out_23
);
W_reg_53_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x29_out_24,
   R => '0',
   Q => W_reg_53_24
);
W_reg_53_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x29_out_25,
   R => '0',
   Q => W_reg_53_25
);
W_reg_53_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x29_out_26,
   R => '0',
   Q => W_reg_53_26
);
W_reg_53_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x29_out_27,
   R => '0',
   Q => W_reg_53_27
);
W_reg_53_27_i_1 : CARRY4
 port map (
   CI => W_reg_53_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_53_27_i_5_n_0,
   DI(1) => W_53_27_i_4_n_0,
   DI(2) => W_53_27_i_3_n_0,
   DI(3) => W_53_27_i_2_n_0,
   S(0) => W_53_27_i_9_n_0,
   S(1) => W_53_27_i_8_n_0,
   S(2) => W_53_27_i_7_n_0,
   S(3) => W_53_27_i_6_n_0,
   CO(0) => W_reg_53_27_i_1_n_3,
   CO(1) => W_reg_53_27_i_1_n_2,
   CO(2) => W_reg_53_27_i_1_n_1,
   CO(3) => W_reg_53_27_i_1_n_0,
   O(0) => x29_out_24,
   O(1) => x29_out_25,
   O(2) => x29_out_26,
   O(3) => x29_out_27
);
W_reg_53_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x29_out_28,
   R => '0',
   Q => W_reg_53_28
);
W_reg_53_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x29_out_29,
   R => '0',
   Q => W_reg_53_29
);
W_reg_53_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x29_out_2,
   R => '0',
   Q => W_reg_53_2
);
W_reg_53_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x29_out_30,
   R => '0',
   Q => W_reg_53_30
);
W_reg_53_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x29_out_31,
   R => '0',
   Q => W_reg_53_31
);
W_reg_53_31_i_1 : CARRY4
 port map (
   CI => W_reg_53_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_53_31_i_4_n_0,
   DI(1) => W_53_31_i_3_n_0,
   DI(2) => W_53_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_53_31_i_8_n_0,
   S(1) => W_53_31_i_7_n_0,
   S(2) => W_53_31_i_6_n_0,
   S(3) => W_53_31_i_5_n_0,
   CO(0) => W_reg_53_31_i_1_n_3,
   CO(1) => W_reg_53_31_i_1_n_2,
   CO(2) => W_reg_53_31_i_1_n_1,
   CO(3) => NLW_W_reg_53_31_i_1_CO_UNCONNECTED_3,
   O(0) => x29_out_28,
   O(1) => x29_out_29,
   O(2) => x29_out_30,
   O(3) => x29_out_31
);
W_reg_53_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x29_out_3,
   R => '0',
   Q => W_reg_53_3
);
W_reg_53_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_53_3_i_5_n_0,
   DI(1) => W_53_3_i_4_n_0,
   DI(2) => W_53_3_i_3_n_0,
   DI(3) => W_53_3_i_2_n_0,
   S(0) => W_53_3_i_9_n_0,
   S(1) => W_53_3_i_8_n_0,
   S(2) => W_53_3_i_7_n_0,
   S(3) => W_53_3_i_6_n_0,
   CO(0) => W_reg_53_3_i_1_n_3,
   CO(1) => W_reg_53_3_i_1_n_2,
   CO(2) => W_reg_53_3_i_1_n_1,
   CO(3) => W_reg_53_3_i_1_n_0,
   O(0) => x29_out_0,
   O(1) => x29_out_1,
   O(2) => x29_out_2,
   O(3) => x29_out_3
);
W_reg_53_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x29_out_4,
   R => '0',
   Q => W_reg_53_4
);
W_reg_53_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x29_out_5,
   R => '0',
   Q => W_reg_53_5
);
W_reg_53_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x29_out_6,
   R => '0',
   Q => W_reg_53_6
);
W_reg_53_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x29_out_7,
   R => '0',
   Q => W_reg_53_7
);
W_reg_53_7_i_1 : CARRY4
 port map (
   CI => W_reg_53_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_53_7_i_5_n_0,
   DI(1) => W_53_7_i_4_n_0,
   DI(2) => W_53_7_i_3_n_0,
   DI(3) => W_53_7_i_2_n_0,
   S(0) => W_53_7_i_9_n_0,
   S(1) => W_53_7_i_8_n_0,
   S(2) => W_53_7_i_7_n_0,
   S(3) => W_53_7_i_6_n_0,
   CO(0) => W_reg_53_7_i_1_n_3,
   CO(1) => W_reg_53_7_i_1_n_2,
   CO(2) => W_reg_53_7_i_1_n_1,
   CO(3) => W_reg_53_7_i_1_n_0,
   O(0) => x29_out_4,
   O(1) => x29_out_5,
   O(2) => x29_out_6,
   O(3) => x29_out_7
);
W_reg_53_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x29_out_8,
   R => '0',
   Q => W_reg_53_8
);
W_reg_53_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x29_out_9,
   R => '0',
   Q => W_reg_53_9
);
W_reg_54_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x26_out_0,
   R => '0',
   Q => W_reg_54_0
);
W_reg_54_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x26_out_10,
   R => '0',
   Q => W_reg_54_10
);
W_reg_54_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x26_out_11,
   R => '0',
   Q => W_reg_54_11
);
W_reg_54_11_i_1 : CARRY4
 port map (
   CI => W_reg_54_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_54_11_i_5_n_0,
   DI(1) => W_54_11_i_4_n_0,
   DI(2) => W_54_11_i_3_n_0,
   DI(3) => W_54_11_i_2_n_0,
   S(0) => W_54_11_i_9_n_0,
   S(1) => W_54_11_i_8_n_0,
   S(2) => W_54_11_i_7_n_0,
   S(3) => W_54_11_i_6_n_0,
   CO(0) => W_reg_54_11_i_1_n_3,
   CO(1) => W_reg_54_11_i_1_n_2,
   CO(2) => W_reg_54_11_i_1_n_1,
   CO(3) => W_reg_54_11_i_1_n_0,
   O(0) => x26_out_8,
   O(1) => x26_out_9,
   O(2) => x26_out_10,
   O(3) => x26_out_11
);
W_reg_54_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x26_out_12,
   R => '0',
   Q => W_reg_54_12
);
W_reg_54_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x26_out_13,
   R => '0',
   Q => W_reg_54_13
);
W_reg_54_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x26_out_14,
   R => '0',
   Q => W_reg_54_14
);
W_reg_54_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x26_out_15,
   R => '0',
   Q => W_reg_54_15
);
W_reg_54_15_i_1 : CARRY4
 port map (
   CI => W_reg_54_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_54_15_i_5_n_0,
   DI(1) => W_54_15_i_4_n_0,
   DI(2) => W_54_15_i_3_n_0,
   DI(3) => W_54_15_i_2_n_0,
   S(0) => W_54_15_i_9_n_0,
   S(1) => W_54_15_i_8_n_0,
   S(2) => W_54_15_i_7_n_0,
   S(3) => W_54_15_i_6_n_0,
   CO(0) => W_reg_54_15_i_1_n_3,
   CO(1) => W_reg_54_15_i_1_n_2,
   CO(2) => W_reg_54_15_i_1_n_1,
   CO(3) => W_reg_54_15_i_1_n_0,
   O(0) => x26_out_12,
   O(1) => x26_out_13,
   O(2) => x26_out_14,
   O(3) => x26_out_15
);
W_reg_54_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x26_out_16,
   R => '0',
   Q => W_reg_54_16
);
W_reg_54_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x26_out_17,
   R => '0',
   Q => W_reg_54_17
);
W_reg_54_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x26_out_18,
   R => '0',
   Q => W_reg_54_18
);
W_reg_54_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x26_out_19,
   R => '0',
   Q => W_reg_54_19
);
W_reg_54_19_i_1 : CARRY4
 port map (
   CI => W_reg_54_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_54_19_i_5_n_0,
   DI(1) => W_54_19_i_4_n_0,
   DI(2) => W_54_19_i_3_n_0,
   DI(3) => W_54_19_i_2_n_0,
   S(0) => W_54_19_i_9_n_0,
   S(1) => W_54_19_i_8_n_0,
   S(2) => W_54_19_i_7_n_0,
   S(3) => W_54_19_i_6_n_0,
   CO(0) => W_reg_54_19_i_1_n_3,
   CO(1) => W_reg_54_19_i_1_n_2,
   CO(2) => W_reg_54_19_i_1_n_1,
   CO(3) => W_reg_54_19_i_1_n_0,
   O(0) => x26_out_16,
   O(1) => x26_out_17,
   O(2) => x26_out_18,
   O(3) => x26_out_19
);
W_reg_54_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x26_out_1,
   R => '0',
   Q => W_reg_54_1
);
W_reg_54_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x26_out_20,
   R => '0',
   Q => W_reg_54_20
);
W_reg_54_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x26_out_21,
   R => '0',
   Q => W_reg_54_21
);
W_reg_54_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x26_out_22,
   R => '0',
   Q => W_reg_54_22
);
W_reg_54_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x26_out_23,
   R => '0',
   Q => W_reg_54_23
);
W_reg_54_23_i_1 : CARRY4
 port map (
   CI => W_reg_54_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_54_23_i_5_n_0,
   DI(1) => W_54_23_i_4_n_0,
   DI(2) => W_54_23_i_3_n_0,
   DI(3) => W_54_23_i_2_n_0,
   S(0) => W_54_23_i_9_n_0,
   S(1) => W_54_23_i_8_n_0,
   S(2) => W_54_23_i_7_n_0,
   S(3) => W_54_23_i_6_n_0,
   CO(0) => W_reg_54_23_i_1_n_3,
   CO(1) => W_reg_54_23_i_1_n_2,
   CO(2) => W_reg_54_23_i_1_n_1,
   CO(3) => W_reg_54_23_i_1_n_0,
   O(0) => x26_out_20,
   O(1) => x26_out_21,
   O(2) => x26_out_22,
   O(3) => x26_out_23
);
W_reg_54_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x26_out_24,
   R => '0',
   Q => W_reg_54_24
);
W_reg_54_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x26_out_25,
   R => '0',
   Q => W_reg_54_25
);
W_reg_54_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x26_out_26,
   R => '0',
   Q => W_reg_54_26
);
W_reg_54_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x26_out_27,
   R => '0',
   Q => W_reg_54_27
);
W_reg_54_27_i_1 : CARRY4
 port map (
   CI => W_reg_54_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_54_27_i_5_n_0,
   DI(1) => W_54_27_i_4_n_0,
   DI(2) => W_54_27_i_3_n_0,
   DI(3) => W_54_27_i_2_n_0,
   S(0) => W_54_27_i_9_n_0,
   S(1) => W_54_27_i_8_n_0,
   S(2) => W_54_27_i_7_n_0,
   S(3) => W_54_27_i_6_n_0,
   CO(0) => W_reg_54_27_i_1_n_3,
   CO(1) => W_reg_54_27_i_1_n_2,
   CO(2) => W_reg_54_27_i_1_n_1,
   CO(3) => W_reg_54_27_i_1_n_0,
   O(0) => x26_out_24,
   O(1) => x26_out_25,
   O(2) => x26_out_26,
   O(3) => x26_out_27
);
W_reg_54_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x26_out_28,
   R => '0',
   Q => W_reg_54_28
);
W_reg_54_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x26_out_29,
   R => '0',
   Q => W_reg_54_29
);
W_reg_54_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x26_out_2,
   R => '0',
   Q => W_reg_54_2
);
W_reg_54_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x26_out_30,
   R => '0',
   Q => W_reg_54_30
);
W_reg_54_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x26_out_31,
   R => '0',
   Q => W_reg_54_31
);
W_reg_54_31_i_1 : CARRY4
 port map (
   CI => W_reg_54_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_54_31_i_4_n_0,
   DI(1) => W_54_31_i_3_n_0,
   DI(2) => W_54_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_54_31_i_8_n_0,
   S(1) => W_54_31_i_7_n_0,
   S(2) => W_54_31_i_6_n_0,
   S(3) => W_54_31_i_5_n_0,
   CO(0) => W_reg_54_31_i_1_n_3,
   CO(1) => W_reg_54_31_i_1_n_2,
   CO(2) => W_reg_54_31_i_1_n_1,
   CO(3) => NLW_W_reg_54_31_i_1_CO_UNCONNECTED_3,
   O(0) => x26_out_28,
   O(1) => x26_out_29,
   O(2) => x26_out_30,
   O(3) => x26_out_31
);
W_reg_54_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x26_out_3,
   R => '0',
   Q => W_reg_54_3
);
W_reg_54_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_54_3_i_5_n_0,
   DI(1) => W_54_3_i_4_n_0,
   DI(2) => W_54_3_i_3_n_0,
   DI(3) => W_54_3_i_2_n_0,
   S(0) => W_54_3_i_9_n_0,
   S(1) => W_54_3_i_8_n_0,
   S(2) => W_54_3_i_7_n_0,
   S(3) => W_54_3_i_6_n_0,
   CO(0) => W_reg_54_3_i_1_n_3,
   CO(1) => W_reg_54_3_i_1_n_2,
   CO(2) => W_reg_54_3_i_1_n_1,
   CO(3) => W_reg_54_3_i_1_n_0,
   O(0) => x26_out_0,
   O(1) => x26_out_1,
   O(2) => x26_out_2,
   O(3) => x26_out_3
);
W_reg_54_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x26_out_4,
   R => '0',
   Q => W_reg_54_4
);
W_reg_54_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x26_out_5,
   R => '0',
   Q => W_reg_54_5
);
W_reg_54_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x26_out_6,
   R => '0',
   Q => W_reg_54_6
);
W_reg_54_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x26_out_7,
   R => '0',
   Q => W_reg_54_7
);
W_reg_54_7_i_1 : CARRY4
 port map (
   CI => W_reg_54_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_54_7_i_5_n_0,
   DI(1) => W_54_7_i_4_n_0,
   DI(2) => W_54_7_i_3_n_0,
   DI(3) => W_54_7_i_2_n_0,
   S(0) => W_54_7_i_9_n_0,
   S(1) => W_54_7_i_8_n_0,
   S(2) => W_54_7_i_7_n_0,
   S(3) => W_54_7_i_6_n_0,
   CO(0) => W_reg_54_7_i_1_n_3,
   CO(1) => W_reg_54_7_i_1_n_2,
   CO(2) => W_reg_54_7_i_1_n_1,
   CO(3) => W_reg_54_7_i_1_n_0,
   O(0) => x26_out_4,
   O(1) => x26_out_5,
   O(2) => x26_out_6,
   O(3) => x26_out_7
);
W_reg_54_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x26_out_8,
   R => '0',
   Q => W_reg_54_8
);
W_reg_54_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x26_out_9,
   R => '0',
   Q => W_reg_54_9
);
W_reg_55_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x23_out_0,
   R => '0',
   Q => W_reg_55_0
);
W_reg_55_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x23_out_10,
   R => '0',
   Q => W_reg_55_10
);
W_reg_55_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x23_out_11,
   R => '0',
   Q => W_reg_55_11
);
W_reg_55_11_i_1 : CARRY4
 port map (
   CI => W_reg_55_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_55_11_i_5_n_0,
   DI(1) => W_55_11_i_4_n_0,
   DI(2) => W_55_11_i_3_n_0,
   DI(3) => W_55_11_i_2_n_0,
   S(0) => W_55_11_i_9_n_0,
   S(1) => W_55_11_i_8_n_0,
   S(2) => W_55_11_i_7_n_0,
   S(3) => W_55_11_i_6_n_0,
   CO(0) => W_reg_55_11_i_1_n_3,
   CO(1) => W_reg_55_11_i_1_n_2,
   CO(2) => W_reg_55_11_i_1_n_1,
   CO(3) => W_reg_55_11_i_1_n_0,
   O(0) => x23_out_8,
   O(1) => x23_out_9,
   O(2) => x23_out_10,
   O(3) => x23_out_11
);
W_reg_55_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x23_out_12,
   R => '0',
   Q => W_reg_55_12
);
W_reg_55_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x23_out_13,
   R => '0',
   Q => W_reg_55_13
);
W_reg_55_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x23_out_14,
   R => '0',
   Q => W_reg_55_14
);
W_reg_55_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x23_out_15,
   R => '0',
   Q => W_reg_55_15
);
W_reg_55_15_i_1 : CARRY4
 port map (
   CI => W_reg_55_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_55_15_i_5_n_0,
   DI(1) => W_55_15_i_4_n_0,
   DI(2) => W_55_15_i_3_n_0,
   DI(3) => W_55_15_i_2_n_0,
   S(0) => W_55_15_i_9_n_0,
   S(1) => W_55_15_i_8_n_0,
   S(2) => W_55_15_i_7_n_0,
   S(3) => W_55_15_i_6_n_0,
   CO(0) => W_reg_55_15_i_1_n_3,
   CO(1) => W_reg_55_15_i_1_n_2,
   CO(2) => W_reg_55_15_i_1_n_1,
   CO(3) => W_reg_55_15_i_1_n_0,
   O(0) => x23_out_12,
   O(1) => x23_out_13,
   O(2) => x23_out_14,
   O(3) => x23_out_15
);
W_reg_55_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x23_out_16,
   R => '0',
   Q => W_reg_55_16
);
W_reg_55_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x23_out_17,
   R => '0',
   Q => W_reg_55_17
);
W_reg_55_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x23_out_18,
   R => '0',
   Q => W_reg_55_18
);
W_reg_55_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x23_out_19,
   R => '0',
   Q => W_reg_55_19
);
W_reg_55_19_i_1 : CARRY4
 port map (
   CI => W_reg_55_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_55_19_i_5_n_0,
   DI(1) => W_55_19_i_4_n_0,
   DI(2) => W_55_19_i_3_n_0,
   DI(3) => W_55_19_i_2_n_0,
   S(0) => W_55_19_i_9_n_0,
   S(1) => W_55_19_i_8_n_0,
   S(2) => W_55_19_i_7_n_0,
   S(3) => W_55_19_i_6_n_0,
   CO(0) => W_reg_55_19_i_1_n_3,
   CO(1) => W_reg_55_19_i_1_n_2,
   CO(2) => W_reg_55_19_i_1_n_1,
   CO(3) => W_reg_55_19_i_1_n_0,
   O(0) => x23_out_16,
   O(1) => x23_out_17,
   O(2) => x23_out_18,
   O(3) => x23_out_19
);
W_reg_55_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x23_out_1,
   R => '0',
   Q => W_reg_55_1
);
W_reg_55_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x23_out_20,
   R => '0',
   Q => W_reg_55_20
);
W_reg_55_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x23_out_21,
   R => '0',
   Q => W_reg_55_21
);
W_reg_55_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x23_out_22,
   R => '0',
   Q => W_reg_55_22
);
W_reg_55_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x23_out_23,
   R => '0',
   Q => W_reg_55_23
);
W_reg_55_23_i_1 : CARRY4
 port map (
   CI => W_reg_55_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_55_23_i_5_n_0,
   DI(1) => W_55_23_i_4_n_0,
   DI(2) => W_55_23_i_3_n_0,
   DI(3) => W_55_23_i_2_n_0,
   S(0) => W_55_23_i_9_n_0,
   S(1) => W_55_23_i_8_n_0,
   S(2) => W_55_23_i_7_n_0,
   S(3) => W_55_23_i_6_n_0,
   CO(0) => W_reg_55_23_i_1_n_3,
   CO(1) => W_reg_55_23_i_1_n_2,
   CO(2) => W_reg_55_23_i_1_n_1,
   CO(3) => W_reg_55_23_i_1_n_0,
   O(0) => x23_out_20,
   O(1) => x23_out_21,
   O(2) => x23_out_22,
   O(3) => x23_out_23
);
W_reg_55_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x23_out_24,
   R => '0',
   Q => W_reg_55_24
);
W_reg_55_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x23_out_25,
   R => '0',
   Q => W_reg_55_25
);
W_reg_55_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x23_out_26,
   R => '0',
   Q => W_reg_55_26
);
W_reg_55_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x23_out_27,
   R => '0',
   Q => W_reg_55_27
);
W_reg_55_27_i_1 : CARRY4
 port map (
   CI => W_reg_55_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_55_27_i_5_n_0,
   DI(1) => W_55_27_i_4_n_0,
   DI(2) => W_55_27_i_3_n_0,
   DI(3) => W_55_27_i_2_n_0,
   S(0) => W_55_27_i_9_n_0,
   S(1) => W_55_27_i_8_n_0,
   S(2) => W_55_27_i_7_n_0,
   S(3) => W_55_27_i_6_n_0,
   CO(0) => W_reg_55_27_i_1_n_3,
   CO(1) => W_reg_55_27_i_1_n_2,
   CO(2) => W_reg_55_27_i_1_n_1,
   CO(3) => W_reg_55_27_i_1_n_0,
   O(0) => x23_out_24,
   O(1) => x23_out_25,
   O(2) => x23_out_26,
   O(3) => x23_out_27
);
W_reg_55_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x23_out_28,
   R => '0',
   Q => W_reg_55_28
);
W_reg_55_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x23_out_29,
   R => '0',
   Q => W_reg_55_29
);
W_reg_55_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x23_out_2,
   R => '0',
   Q => W_reg_55_2
);
W_reg_55_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x23_out_30,
   R => '0',
   Q => W_reg_55_30
);
W_reg_55_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x23_out_31,
   R => '0',
   Q => W_reg_55_31
);
W_reg_55_31_i_1 : CARRY4
 port map (
   CI => W_reg_55_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_55_31_i_4_n_0,
   DI(1) => W_55_31_i_3_n_0,
   DI(2) => W_55_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_55_31_i_8_n_0,
   S(1) => W_55_31_i_7_n_0,
   S(2) => W_55_31_i_6_n_0,
   S(3) => W_55_31_i_5_n_0,
   CO(0) => W_reg_55_31_i_1_n_3,
   CO(1) => W_reg_55_31_i_1_n_2,
   CO(2) => W_reg_55_31_i_1_n_1,
   CO(3) => NLW_W_reg_55_31_i_1_CO_UNCONNECTED_3,
   O(0) => x23_out_28,
   O(1) => x23_out_29,
   O(2) => x23_out_30,
   O(3) => x23_out_31
);
W_reg_55_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x23_out_3,
   R => '0',
   Q => W_reg_55_3
);
W_reg_55_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_55_3_i_5_n_0,
   DI(1) => W_55_3_i_4_n_0,
   DI(2) => W_55_3_i_3_n_0,
   DI(3) => W_55_3_i_2_n_0,
   S(0) => W_55_3_i_9_n_0,
   S(1) => W_55_3_i_8_n_0,
   S(2) => W_55_3_i_7_n_0,
   S(3) => W_55_3_i_6_n_0,
   CO(0) => W_reg_55_3_i_1_n_3,
   CO(1) => W_reg_55_3_i_1_n_2,
   CO(2) => W_reg_55_3_i_1_n_1,
   CO(3) => W_reg_55_3_i_1_n_0,
   O(0) => x23_out_0,
   O(1) => x23_out_1,
   O(2) => x23_out_2,
   O(3) => x23_out_3
);
W_reg_55_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x23_out_4,
   R => '0',
   Q => W_reg_55_4
);
W_reg_55_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x23_out_5,
   R => '0',
   Q => W_reg_55_5
);
W_reg_55_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x23_out_6,
   R => '0',
   Q => W_reg_55_6
);
W_reg_55_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x23_out_7,
   R => '0',
   Q => W_reg_55_7
);
W_reg_55_7_i_1 : CARRY4
 port map (
   CI => W_reg_55_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_55_7_i_5_n_0,
   DI(1) => W_55_7_i_4_n_0,
   DI(2) => W_55_7_i_3_n_0,
   DI(3) => W_55_7_i_2_n_0,
   S(0) => W_55_7_i_9_n_0,
   S(1) => W_55_7_i_8_n_0,
   S(2) => W_55_7_i_7_n_0,
   S(3) => W_55_7_i_6_n_0,
   CO(0) => W_reg_55_7_i_1_n_3,
   CO(1) => W_reg_55_7_i_1_n_2,
   CO(2) => W_reg_55_7_i_1_n_1,
   CO(3) => W_reg_55_7_i_1_n_0,
   O(0) => x23_out_4,
   O(1) => x23_out_5,
   O(2) => x23_out_6,
   O(3) => x23_out_7
);
W_reg_55_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x23_out_8,
   R => '0',
   Q => W_reg_55_8
);
W_reg_55_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x23_out_9,
   R => '0',
   Q => W_reg_55_9
);
W_reg_56_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x20_out_0,
   R => '0',
   Q => W_reg_56_0
);
W_reg_56_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x20_out_10,
   R => '0',
   Q => W_reg_56_10
);
W_reg_56_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x20_out_11,
   R => '0',
   Q => W_reg_56_11
);
W_reg_56_11_i_1 : CARRY4
 port map (
   CI => W_reg_56_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_56_11_i_5_n_0,
   DI(1) => W_56_11_i_4_n_0,
   DI(2) => W_56_11_i_3_n_0,
   DI(3) => W_56_11_i_2_n_0,
   S(0) => W_56_11_i_9_n_0,
   S(1) => W_56_11_i_8_n_0,
   S(2) => W_56_11_i_7_n_0,
   S(3) => W_56_11_i_6_n_0,
   CO(0) => W_reg_56_11_i_1_n_3,
   CO(1) => W_reg_56_11_i_1_n_2,
   CO(2) => W_reg_56_11_i_1_n_1,
   CO(3) => W_reg_56_11_i_1_n_0,
   O(0) => x20_out_8,
   O(1) => x20_out_9,
   O(2) => x20_out_10,
   O(3) => x20_out_11
);
W_reg_56_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x20_out_12,
   R => '0',
   Q => W_reg_56_12
);
W_reg_56_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x20_out_13,
   R => '0',
   Q => W_reg_56_13
);
W_reg_56_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x20_out_14,
   R => '0',
   Q => W_reg_56_14
);
W_reg_56_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x20_out_15,
   R => '0',
   Q => W_reg_56_15
);
W_reg_56_15_i_1 : CARRY4
 port map (
   CI => W_reg_56_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_56_15_i_5_n_0,
   DI(1) => W_56_15_i_4_n_0,
   DI(2) => W_56_15_i_3_n_0,
   DI(3) => W_56_15_i_2_n_0,
   S(0) => W_56_15_i_9_n_0,
   S(1) => W_56_15_i_8_n_0,
   S(2) => W_56_15_i_7_n_0,
   S(3) => W_56_15_i_6_n_0,
   CO(0) => W_reg_56_15_i_1_n_3,
   CO(1) => W_reg_56_15_i_1_n_2,
   CO(2) => W_reg_56_15_i_1_n_1,
   CO(3) => W_reg_56_15_i_1_n_0,
   O(0) => x20_out_12,
   O(1) => x20_out_13,
   O(2) => x20_out_14,
   O(3) => x20_out_15
);
W_reg_56_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x20_out_16,
   R => '0',
   Q => W_reg_56_16
);
W_reg_56_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x20_out_17,
   R => '0',
   Q => W_reg_56_17
);
W_reg_56_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x20_out_18,
   R => '0',
   Q => W_reg_56_18
);
W_reg_56_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x20_out_19,
   R => '0',
   Q => W_reg_56_19
);
W_reg_56_19_i_1 : CARRY4
 port map (
   CI => W_reg_56_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_56_19_i_5_n_0,
   DI(1) => W_56_19_i_4_n_0,
   DI(2) => W_56_19_i_3_n_0,
   DI(3) => W_56_19_i_2_n_0,
   S(0) => W_56_19_i_9_n_0,
   S(1) => W_56_19_i_8_n_0,
   S(2) => W_56_19_i_7_n_0,
   S(3) => W_56_19_i_6_n_0,
   CO(0) => W_reg_56_19_i_1_n_3,
   CO(1) => W_reg_56_19_i_1_n_2,
   CO(2) => W_reg_56_19_i_1_n_1,
   CO(3) => W_reg_56_19_i_1_n_0,
   O(0) => x20_out_16,
   O(1) => x20_out_17,
   O(2) => x20_out_18,
   O(3) => x20_out_19
);
W_reg_56_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x20_out_1,
   R => '0',
   Q => W_reg_56_1
);
W_reg_56_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x20_out_20,
   R => '0',
   Q => W_reg_56_20
);
W_reg_56_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x20_out_21,
   R => '0',
   Q => W_reg_56_21
);
W_reg_56_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x20_out_22,
   R => '0',
   Q => W_reg_56_22
);
W_reg_56_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x20_out_23,
   R => '0',
   Q => W_reg_56_23
);
W_reg_56_23_i_1 : CARRY4
 port map (
   CI => W_reg_56_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_56_23_i_5_n_0,
   DI(1) => W_56_23_i_4_n_0,
   DI(2) => W_56_23_i_3_n_0,
   DI(3) => W_56_23_i_2_n_0,
   S(0) => W_56_23_i_9_n_0,
   S(1) => W_56_23_i_8_n_0,
   S(2) => W_56_23_i_7_n_0,
   S(3) => W_56_23_i_6_n_0,
   CO(0) => W_reg_56_23_i_1_n_3,
   CO(1) => W_reg_56_23_i_1_n_2,
   CO(2) => W_reg_56_23_i_1_n_1,
   CO(3) => W_reg_56_23_i_1_n_0,
   O(0) => x20_out_20,
   O(1) => x20_out_21,
   O(2) => x20_out_22,
   O(3) => x20_out_23
);
W_reg_56_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x20_out_24,
   R => '0',
   Q => W_reg_56_24
);
W_reg_56_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x20_out_25,
   R => '0',
   Q => W_reg_56_25
);
W_reg_56_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x20_out_26,
   R => '0',
   Q => W_reg_56_26
);
W_reg_56_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x20_out_27,
   R => '0',
   Q => W_reg_56_27
);
W_reg_56_27_i_1 : CARRY4
 port map (
   CI => W_reg_56_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_56_27_i_5_n_0,
   DI(1) => W_56_27_i_4_n_0,
   DI(2) => W_56_27_i_3_n_0,
   DI(3) => W_56_27_i_2_n_0,
   S(0) => W_56_27_i_9_n_0,
   S(1) => W_56_27_i_8_n_0,
   S(2) => W_56_27_i_7_n_0,
   S(3) => W_56_27_i_6_n_0,
   CO(0) => W_reg_56_27_i_1_n_3,
   CO(1) => W_reg_56_27_i_1_n_2,
   CO(2) => W_reg_56_27_i_1_n_1,
   CO(3) => W_reg_56_27_i_1_n_0,
   O(0) => x20_out_24,
   O(1) => x20_out_25,
   O(2) => x20_out_26,
   O(3) => x20_out_27
);
W_reg_56_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x20_out_28,
   R => '0',
   Q => W_reg_56_28
);
W_reg_56_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x20_out_29,
   R => '0',
   Q => W_reg_56_29
);
W_reg_56_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x20_out_2,
   R => '0',
   Q => W_reg_56_2
);
W_reg_56_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x20_out_30,
   R => '0',
   Q => W_reg_56_30
);
W_reg_56_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x20_out_31,
   R => '0',
   Q => W_reg_56_31
);
W_reg_56_31_i_1 : CARRY4
 port map (
   CI => W_reg_56_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_56_31_i_4_n_0,
   DI(1) => W_56_31_i_3_n_0,
   DI(2) => W_56_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_56_31_i_8_n_0,
   S(1) => W_56_31_i_7_n_0,
   S(2) => W_56_31_i_6_n_0,
   S(3) => W_56_31_i_5_n_0,
   CO(0) => W_reg_56_31_i_1_n_3,
   CO(1) => W_reg_56_31_i_1_n_2,
   CO(2) => W_reg_56_31_i_1_n_1,
   CO(3) => NLW_W_reg_56_31_i_1_CO_UNCONNECTED_3,
   O(0) => x20_out_28,
   O(1) => x20_out_29,
   O(2) => x20_out_30,
   O(3) => x20_out_31
);
W_reg_56_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x20_out_3,
   R => '0',
   Q => W_reg_56_3
);
W_reg_56_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_56_3_i_5_n_0,
   DI(1) => W_56_3_i_4_n_0,
   DI(2) => W_56_3_i_3_n_0,
   DI(3) => W_56_3_i_2_n_0,
   S(0) => W_56_3_i_9_n_0,
   S(1) => W_56_3_i_8_n_0,
   S(2) => W_56_3_i_7_n_0,
   S(3) => W_56_3_i_6_n_0,
   CO(0) => W_reg_56_3_i_1_n_3,
   CO(1) => W_reg_56_3_i_1_n_2,
   CO(2) => W_reg_56_3_i_1_n_1,
   CO(3) => W_reg_56_3_i_1_n_0,
   O(0) => x20_out_0,
   O(1) => x20_out_1,
   O(2) => x20_out_2,
   O(3) => x20_out_3
);
W_reg_56_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x20_out_4,
   R => '0',
   Q => W_reg_56_4
);
W_reg_56_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x20_out_5,
   R => '0',
   Q => W_reg_56_5
);
W_reg_56_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x20_out_6,
   R => '0',
   Q => W_reg_56_6
);
W_reg_56_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x20_out_7,
   R => '0',
   Q => W_reg_56_7
);
W_reg_56_7_i_1 : CARRY4
 port map (
   CI => W_reg_56_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_56_7_i_5_n_0,
   DI(1) => W_56_7_i_4_n_0,
   DI(2) => W_56_7_i_3_n_0,
   DI(3) => W_56_7_i_2_n_0,
   S(0) => W_56_7_i_9_n_0,
   S(1) => W_56_7_i_8_n_0,
   S(2) => W_56_7_i_7_n_0,
   S(3) => W_56_7_i_6_n_0,
   CO(0) => W_reg_56_7_i_1_n_3,
   CO(1) => W_reg_56_7_i_1_n_2,
   CO(2) => W_reg_56_7_i_1_n_1,
   CO(3) => W_reg_56_7_i_1_n_0,
   O(0) => x20_out_4,
   O(1) => x20_out_5,
   O(2) => x20_out_6,
   O(3) => x20_out_7
);
W_reg_56_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x20_out_8,
   R => '0',
   Q => W_reg_56_8
);
W_reg_56_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x20_out_9,
   R => '0',
   Q => W_reg_56_9
);
W_reg_57_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x17_out_0,
   R => '0',
   Q => W_reg_57_0
);
W_reg_57_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x17_out_10,
   R => '0',
   Q => W_reg_57_10
);
W_reg_57_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x17_out_11,
   R => '0',
   Q => W_reg_57_11
);
W_reg_57_11_i_1 : CARRY4
 port map (
   CI => W_reg_57_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_57_11_i_5_n_0,
   DI(1) => W_57_11_i_4_n_0,
   DI(2) => W_57_11_i_3_n_0,
   DI(3) => W_57_11_i_2_n_0,
   S(0) => W_57_11_i_9_n_0,
   S(1) => W_57_11_i_8_n_0,
   S(2) => W_57_11_i_7_n_0,
   S(3) => W_57_11_i_6_n_0,
   CO(0) => W_reg_57_11_i_1_n_3,
   CO(1) => W_reg_57_11_i_1_n_2,
   CO(2) => W_reg_57_11_i_1_n_1,
   CO(3) => W_reg_57_11_i_1_n_0,
   O(0) => x17_out_8,
   O(1) => x17_out_9,
   O(2) => x17_out_10,
   O(3) => x17_out_11
);
W_reg_57_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x17_out_12,
   R => '0',
   Q => W_reg_57_12
);
W_reg_57_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x17_out_13,
   R => '0',
   Q => W_reg_57_13
);
W_reg_57_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x17_out_14,
   R => '0',
   Q => W_reg_57_14
);
W_reg_57_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x17_out_15,
   R => '0',
   Q => W_reg_57_15
);
W_reg_57_15_i_1 : CARRY4
 port map (
   CI => W_reg_57_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_57_15_i_5_n_0,
   DI(1) => W_57_15_i_4_n_0,
   DI(2) => W_57_15_i_3_n_0,
   DI(3) => W_57_15_i_2_n_0,
   S(0) => W_57_15_i_9_n_0,
   S(1) => W_57_15_i_8_n_0,
   S(2) => W_57_15_i_7_n_0,
   S(3) => W_57_15_i_6_n_0,
   CO(0) => W_reg_57_15_i_1_n_3,
   CO(1) => W_reg_57_15_i_1_n_2,
   CO(2) => W_reg_57_15_i_1_n_1,
   CO(3) => W_reg_57_15_i_1_n_0,
   O(0) => x17_out_12,
   O(1) => x17_out_13,
   O(2) => x17_out_14,
   O(3) => x17_out_15
);
W_reg_57_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x17_out_16,
   R => '0',
   Q => W_reg_57_16
);
W_reg_57_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x17_out_17,
   R => '0',
   Q => W_reg_57_17
);
W_reg_57_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x17_out_18,
   R => '0',
   Q => W_reg_57_18
);
W_reg_57_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x17_out_19,
   R => '0',
   Q => W_reg_57_19
);
W_reg_57_19_i_1 : CARRY4
 port map (
   CI => W_reg_57_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_57_19_i_5_n_0,
   DI(1) => W_57_19_i_4_n_0,
   DI(2) => W_57_19_i_3_n_0,
   DI(3) => W_57_19_i_2_n_0,
   S(0) => W_57_19_i_9_n_0,
   S(1) => W_57_19_i_8_n_0,
   S(2) => W_57_19_i_7_n_0,
   S(3) => W_57_19_i_6_n_0,
   CO(0) => W_reg_57_19_i_1_n_3,
   CO(1) => W_reg_57_19_i_1_n_2,
   CO(2) => W_reg_57_19_i_1_n_1,
   CO(3) => W_reg_57_19_i_1_n_0,
   O(0) => x17_out_16,
   O(1) => x17_out_17,
   O(2) => x17_out_18,
   O(3) => x17_out_19
);
W_reg_57_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x17_out_1,
   R => '0',
   Q => W_reg_57_1
);
W_reg_57_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x17_out_20,
   R => '0',
   Q => W_reg_57_20
);
W_reg_57_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x17_out_21,
   R => '0',
   Q => W_reg_57_21
);
W_reg_57_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x17_out_22,
   R => '0',
   Q => W_reg_57_22
);
W_reg_57_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x17_out_23,
   R => '0',
   Q => W_reg_57_23
);
W_reg_57_23_i_1 : CARRY4
 port map (
   CI => W_reg_57_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_57_23_i_5_n_0,
   DI(1) => W_57_23_i_4_n_0,
   DI(2) => W_57_23_i_3_n_0,
   DI(3) => W_57_23_i_2_n_0,
   S(0) => W_57_23_i_9_n_0,
   S(1) => W_57_23_i_8_n_0,
   S(2) => W_57_23_i_7_n_0,
   S(3) => W_57_23_i_6_n_0,
   CO(0) => W_reg_57_23_i_1_n_3,
   CO(1) => W_reg_57_23_i_1_n_2,
   CO(2) => W_reg_57_23_i_1_n_1,
   CO(3) => W_reg_57_23_i_1_n_0,
   O(0) => x17_out_20,
   O(1) => x17_out_21,
   O(2) => x17_out_22,
   O(3) => x17_out_23
);
W_reg_57_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x17_out_24,
   R => '0',
   Q => W_reg_57_24
);
W_reg_57_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x17_out_25,
   R => '0',
   Q => W_reg_57_25
);
W_reg_57_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x17_out_26,
   R => '0',
   Q => W_reg_57_26
);
W_reg_57_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x17_out_27,
   R => '0',
   Q => W_reg_57_27
);
W_reg_57_27_i_1 : CARRY4
 port map (
   CI => W_reg_57_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_57_27_i_5_n_0,
   DI(1) => W_57_27_i_4_n_0,
   DI(2) => W_57_27_i_3_n_0,
   DI(3) => W_57_27_i_2_n_0,
   S(0) => W_57_27_i_9_n_0,
   S(1) => W_57_27_i_8_n_0,
   S(2) => W_57_27_i_7_n_0,
   S(3) => W_57_27_i_6_n_0,
   CO(0) => W_reg_57_27_i_1_n_3,
   CO(1) => W_reg_57_27_i_1_n_2,
   CO(2) => W_reg_57_27_i_1_n_1,
   CO(3) => W_reg_57_27_i_1_n_0,
   O(0) => x17_out_24,
   O(1) => x17_out_25,
   O(2) => x17_out_26,
   O(3) => x17_out_27
);
W_reg_57_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x17_out_28,
   R => '0',
   Q => W_reg_57_28
);
W_reg_57_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x17_out_29,
   R => '0',
   Q => W_reg_57_29
);
W_reg_57_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x17_out_2,
   R => '0',
   Q => W_reg_57_2
);
W_reg_57_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x17_out_30,
   R => '0',
   Q => W_reg_57_30
);
W_reg_57_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x17_out_31,
   R => '0',
   Q => W_reg_57_31
);
W_reg_57_31_i_1 : CARRY4
 port map (
   CI => W_reg_57_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_57_31_i_4_n_0,
   DI(1) => W_57_31_i_3_n_0,
   DI(2) => W_57_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_57_31_i_8_n_0,
   S(1) => W_57_31_i_7_n_0,
   S(2) => W_57_31_i_6_n_0,
   S(3) => W_57_31_i_5_n_0,
   CO(0) => W_reg_57_31_i_1_n_3,
   CO(1) => W_reg_57_31_i_1_n_2,
   CO(2) => W_reg_57_31_i_1_n_1,
   CO(3) => NLW_W_reg_57_31_i_1_CO_UNCONNECTED_3,
   O(0) => x17_out_28,
   O(1) => x17_out_29,
   O(2) => x17_out_30,
   O(3) => x17_out_31
);
W_reg_57_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x17_out_3,
   R => '0',
   Q => W_reg_57_3
);
W_reg_57_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_57_3_i_5_n_0,
   DI(1) => W_57_3_i_4_n_0,
   DI(2) => W_57_3_i_3_n_0,
   DI(3) => W_57_3_i_2_n_0,
   S(0) => W_57_3_i_9_n_0,
   S(1) => W_57_3_i_8_n_0,
   S(2) => W_57_3_i_7_n_0,
   S(3) => W_57_3_i_6_n_0,
   CO(0) => W_reg_57_3_i_1_n_3,
   CO(1) => W_reg_57_3_i_1_n_2,
   CO(2) => W_reg_57_3_i_1_n_1,
   CO(3) => W_reg_57_3_i_1_n_0,
   O(0) => x17_out_0,
   O(1) => x17_out_1,
   O(2) => x17_out_2,
   O(3) => x17_out_3
);
W_reg_57_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x17_out_4,
   R => '0',
   Q => W_reg_57_4
);
W_reg_57_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x17_out_5,
   R => '0',
   Q => W_reg_57_5
);
W_reg_57_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x17_out_6,
   R => '0',
   Q => W_reg_57_6
);
W_reg_57_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x17_out_7,
   R => '0',
   Q => W_reg_57_7
);
W_reg_57_7_i_1 : CARRY4
 port map (
   CI => W_reg_57_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_57_7_i_5_n_0,
   DI(1) => W_57_7_i_4_n_0,
   DI(2) => W_57_7_i_3_n_0,
   DI(3) => W_57_7_i_2_n_0,
   S(0) => W_57_7_i_9_n_0,
   S(1) => W_57_7_i_8_n_0,
   S(2) => W_57_7_i_7_n_0,
   S(3) => W_57_7_i_6_n_0,
   CO(0) => W_reg_57_7_i_1_n_3,
   CO(1) => W_reg_57_7_i_1_n_2,
   CO(2) => W_reg_57_7_i_1_n_1,
   CO(3) => W_reg_57_7_i_1_n_0,
   O(0) => x17_out_4,
   O(1) => x17_out_5,
   O(2) => x17_out_6,
   O(3) => x17_out_7
);
W_reg_57_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x17_out_8,
   R => '0',
   Q => W_reg_57_8
);
W_reg_57_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x17_out_9,
   R => '0',
   Q => W_reg_57_9
);
W_reg_58_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x14_out_0,
   R => '0',
   Q => W_reg_58_0
);
W_reg_58_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x14_out_10,
   R => '0',
   Q => W_reg_58_10
);
W_reg_58_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x14_out_11,
   R => '0',
   Q => W_reg_58_11
);
W_reg_58_11_i_1 : CARRY4
 port map (
   CI => W_reg_58_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_58_11_i_5_n_0,
   DI(1) => W_58_11_i_4_n_0,
   DI(2) => W_58_11_i_3_n_0,
   DI(3) => W_58_11_i_2_n_0,
   S(0) => W_58_11_i_9_n_0,
   S(1) => W_58_11_i_8_n_0,
   S(2) => W_58_11_i_7_n_0,
   S(3) => W_58_11_i_6_n_0,
   CO(0) => W_reg_58_11_i_1_n_3,
   CO(1) => W_reg_58_11_i_1_n_2,
   CO(2) => W_reg_58_11_i_1_n_1,
   CO(3) => W_reg_58_11_i_1_n_0,
   O(0) => x14_out_8,
   O(1) => x14_out_9,
   O(2) => x14_out_10,
   O(3) => x14_out_11
);
W_reg_58_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x14_out_12,
   R => '0',
   Q => W_reg_58_12
);
W_reg_58_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x14_out_13,
   R => '0',
   Q => W_reg_58_13
);
W_reg_58_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x14_out_14,
   R => '0',
   Q => W_reg_58_14
);
W_reg_58_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x14_out_15,
   R => '0',
   Q => W_reg_58_15
);
W_reg_58_15_i_1 : CARRY4
 port map (
   CI => W_reg_58_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_58_15_i_5_n_0,
   DI(1) => W_58_15_i_4_n_0,
   DI(2) => W_58_15_i_3_n_0,
   DI(3) => W_58_15_i_2_n_0,
   S(0) => W_58_15_i_9_n_0,
   S(1) => W_58_15_i_8_n_0,
   S(2) => W_58_15_i_7_n_0,
   S(3) => W_58_15_i_6_n_0,
   CO(0) => W_reg_58_15_i_1_n_3,
   CO(1) => W_reg_58_15_i_1_n_2,
   CO(2) => W_reg_58_15_i_1_n_1,
   CO(3) => W_reg_58_15_i_1_n_0,
   O(0) => x14_out_12,
   O(1) => x14_out_13,
   O(2) => x14_out_14,
   O(3) => x14_out_15
);
W_reg_58_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x14_out_16,
   R => '0',
   Q => W_reg_58_16
);
W_reg_58_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x14_out_17,
   R => '0',
   Q => W_reg_58_17
);
W_reg_58_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x14_out_18,
   R => '0',
   Q => W_reg_58_18
);
W_reg_58_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x14_out_19,
   R => '0',
   Q => W_reg_58_19
);
W_reg_58_19_i_1 : CARRY4
 port map (
   CI => W_reg_58_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_58_19_i_5_n_0,
   DI(1) => W_58_19_i_4_n_0,
   DI(2) => W_58_19_i_3_n_0,
   DI(3) => W_58_19_i_2_n_0,
   S(0) => W_58_19_i_9_n_0,
   S(1) => W_58_19_i_8_n_0,
   S(2) => W_58_19_i_7_n_0,
   S(3) => W_58_19_i_6_n_0,
   CO(0) => W_reg_58_19_i_1_n_3,
   CO(1) => W_reg_58_19_i_1_n_2,
   CO(2) => W_reg_58_19_i_1_n_1,
   CO(3) => W_reg_58_19_i_1_n_0,
   O(0) => x14_out_16,
   O(1) => x14_out_17,
   O(2) => x14_out_18,
   O(3) => x14_out_19
);
W_reg_58_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x14_out_1,
   R => '0',
   Q => W_reg_58_1
);
W_reg_58_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x14_out_20,
   R => '0',
   Q => W_reg_58_20
);
W_reg_58_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x14_out_21,
   R => '0',
   Q => W_reg_58_21
);
W_reg_58_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x14_out_22,
   R => '0',
   Q => W_reg_58_22
);
W_reg_58_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x14_out_23,
   R => '0',
   Q => W_reg_58_23
);
W_reg_58_23_i_1 : CARRY4
 port map (
   CI => W_reg_58_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_58_23_i_5_n_0,
   DI(1) => W_58_23_i_4_n_0,
   DI(2) => W_58_23_i_3_n_0,
   DI(3) => W_58_23_i_2_n_0,
   S(0) => W_58_23_i_9_n_0,
   S(1) => W_58_23_i_8_n_0,
   S(2) => W_58_23_i_7_n_0,
   S(3) => W_58_23_i_6_n_0,
   CO(0) => W_reg_58_23_i_1_n_3,
   CO(1) => W_reg_58_23_i_1_n_2,
   CO(2) => W_reg_58_23_i_1_n_1,
   CO(3) => W_reg_58_23_i_1_n_0,
   O(0) => x14_out_20,
   O(1) => x14_out_21,
   O(2) => x14_out_22,
   O(3) => x14_out_23
);
W_reg_58_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x14_out_24,
   R => '0',
   Q => W_reg_58_24
);
W_reg_58_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x14_out_25,
   R => '0',
   Q => W_reg_58_25
);
W_reg_58_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x14_out_26,
   R => '0',
   Q => W_reg_58_26
);
W_reg_58_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x14_out_27,
   R => '0',
   Q => W_reg_58_27
);
W_reg_58_27_i_1 : CARRY4
 port map (
   CI => W_reg_58_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_58_27_i_5_n_0,
   DI(1) => W_58_27_i_4_n_0,
   DI(2) => W_58_27_i_3_n_0,
   DI(3) => W_58_27_i_2_n_0,
   S(0) => W_58_27_i_9_n_0,
   S(1) => W_58_27_i_8_n_0,
   S(2) => W_58_27_i_7_n_0,
   S(3) => W_58_27_i_6_n_0,
   CO(0) => W_reg_58_27_i_1_n_3,
   CO(1) => W_reg_58_27_i_1_n_2,
   CO(2) => W_reg_58_27_i_1_n_1,
   CO(3) => W_reg_58_27_i_1_n_0,
   O(0) => x14_out_24,
   O(1) => x14_out_25,
   O(2) => x14_out_26,
   O(3) => x14_out_27
);
W_reg_58_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x14_out_28,
   R => '0',
   Q => W_reg_58_28
);
W_reg_58_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x14_out_29,
   R => '0',
   Q => W_reg_58_29
);
W_reg_58_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x14_out_2,
   R => '0',
   Q => W_reg_58_2
);
W_reg_58_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x14_out_30,
   R => '0',
   Q => W_reg_58_30
);
W_reg_58_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x14_out_31,
   R => '0',
   Q => W_reg_58_31
);
W_reg_58_31_i_1 : CARRY4
 port map (
   CI => W_reg_58_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_58_31_i_4_n_0,
   DI(1) => W_58_31_i_3_n_0,
   DI(2) => W_58_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_58_31_i_8_n_0,
   S(1) => W_58_31_i_7_n_0,
   S(2) => W_58_31_i_6_n_0,
   S(3) => W_58_31_i_5_n_0,
   CO(0) => W_reg_58_31_i_1_n_3,
   CO(1) => W_reg_58_31_i_1_n_2,
   CO(2) => W_reg_58_31_i_1_n_1,
   CO(3) => NLW_W_reg_58_31_i_1_CO_UNCONNECTED_3,
   O(0) => x14_out_28,
   O(1) => x14_out_29,
   O(2) => x14_out_30,
   O(3) => x14_out_31
);
W_reg_58_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x14_out_3,
   R => '0',
   Q => W_reg_58_3
);
W_reg_58_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_58_3_i_5_n_0,
   DI(1) => W_58_3_i_4_n_0,
   DI(2) => W_58_3_i_3_n_0,
   DI(3) => W_58_3_i_2_n_0,
   S(0) => W_58_3_i_9_n_0,
   S(1) => W_58_3_i_8_n_0,
   S(2) => W_58_3_i_7_n_0,
   S(3) => W_58_3_i_6_n_0,
   CO(0) => W_reg_58_3_i_1_n_3,
   CO(1) => W_reg_58_3_i_1_n_2,
   CO(2) => W_reg_58_3_i_1_n_1,
   CO(3) => W_reg_58_3_i_1_n_0,
   O(0) => x14_out_0,
   O(1) => x14_out_1,
   O(2) => x14_out_2,
   O(3) => x14_out_3
);
W_reg_58_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x14_out_4,
   R => '0',
   Q => W_reg_58_4
);
W_reg_58_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x14_out_5,
   R => '0',
   Q => W_reg_58_5
);
W_reg_58_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x14_out_6,
   R => '0',
   Q => W_reg_58_6
);
W_reg_58_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x14_out_7,
   R => '0',
   Q => W_reg_58_7
);
W_reg_58_7_i_1 : CARRY4
 port map (
   CI => W_reg_58_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_58_7_i_5_n_0,
   DI(1) => W_58_7_i_4_n_0,
   DI(2) => W_58_7_i_3_n_0,
   DI(3) => W_58_7_i_2_n_0,
   S(0) => W_58_7_i_9_n_0,
   S(1) => W_58_7_i_8_n_0,
   S(2) => W_58_7_i_7_n_0,
   S(3) => W_58_7_i_6_n_0,
   CO(0) => W_reg_58_7_i_1_n_3,
   CO(1) => W_reg_58_7_i_1_n_2,
   CO(2) => W_reg_58_7_i_1_n_1,
   CO(3) => W_reg_58_7_i_1_n_0,
   O(0) => x14_out_4,
   O(1) => x14_out_5,
   O(2) => x14_out_6,
   O(3) => x14_out_7
);
W_reg_58_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x14_out_8,
   R => '0',
   Q => W_reg_58_8
);
W_reg_58_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x14_out_9,
   R => '0',
   Q => W_reg_58_9
);
W_reg_59_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x11_out_0,
   R => '0',
   Q => W_reg_59_0
);
W_reg_59_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x11_out_10,
   R => '0',
   Q => W_reg_59_10
);
W_reg_59_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x11_out_11,
   R => '0',
   Q => W_reg_59_11
);
W_reg_59_11_i_1 : CARRY4
 port map (
   CI => W_reg_59_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_59_11_i_5_n_0,
   DI(1) => W_59_11_i_4_n_0,
   DI(2) => W_59_11_i_3_n_0,
   DI(3) => W_59_11_i_2_n_0,
   S(0) => W_59_11_i_9_n_0,
   S(1) => W_59_11_i_8_n_0,
   S(2) => W_59_11_i_7_n_0,
   S(3) => W_59_11_i_6_n_0,
   CO(0) => W_reg_59_11_i_1_n_3,
   CO(1) => W_reg_59_11_i_1_n_2,
   CO(2) => W_reg_59_11_i_1_n_1,
   CO(3) => W_reg_59_11_i_1_n_0,
   O(0) => x11_out_8,
   O(1) => x11_out_9,
   O(2) => x11_out_10,
   O(3) => x11_out_11
);
W_reg_59_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x11_out_12,
   R => '0',
   Q => W_reg_59_12
);
W_reg_59_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x11_out_13,
   R => '0',
   Q => W_reg_59_13
);
W_reg_59_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x11_out_14,
   R => '0',
   Q => W_reg_59_14
);
W_reg_59_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x11_out_15,
   R => '0',
   Q => W_reg_59_15
);
W_reg_59_15_i_1 : CARRY4
 port map (
   CI => W_reg_59_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_59_15_i_5_n_0,
   DI(1) => W_59_15_i_4_n_0,
   DI(2) => W_59_15_i_3_n_0,
   DI(3) => W_59_15_i_2_n_0,
   S(0) => W_59_15_i_9_n_0,
   S(1) => W_59_15_i_8_n_0,
   S(2) => W_59_15_i_7_n_0,
   S(3) => W_59_15_i_6_n_0,
   CO(0) => W_reg_59_15_i_1_n_3,
   CO(1) => W_reg_59_15_i_1_n_2,
   CO(2) => W_reg_59_15_i_1_n_1,
   CO(3) => W_reg_59_15_i_1_n_0,
   O(0) => x11_out_12,
   O(1) => x11_out_13,
   O(2) => x11_out_14,
   O(3) => x11_out_15
);
W_reg_59_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x11_out_16,
   R => '0',
   Q => W_reg_59_16
);
W_reg_59_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x11_out_17,
   R => '0',
   Q => W_reg_59_17
);
W_reg_59_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x11_out_18,
   R => '0',
   Q => W_reg_59_18
);
W_reg_59_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x11_out_19,
   R => '0',
   Q => W_reg_59_19
);
W_reg_59_19_i_1 : CARRY4
 port map (
   CI => W_reg_59_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_59_19_i_5_n_0,
   DI(1) => W_59_19_i_4_n_0,
   DI(2) => W_59_19_i_3_n_0,
   DI(3) => W_59_19_i_2_n_0,
   S(0) => W_59_19_i_9_n_0,
   S(1) => W_59_19_i_8_n_0,
   S(2) => W_59_19_i_7_n_0,
   S(3) => W_59_19_i_6_n_0,
   CO(0) => W_reg_59_19_i_1_n_3,
   CO(1) => W_reg_59_19_i_1_n_2,
   CO(2) => W_reg_59_19_i_1_n_1,
   CO(3) => W_reg_59_19_i_1_n_0,
   O(0) => x11_out_16,
   O(1) => x11_out_17,
   O(2) => x11_out_18,
   O(3) => x11_out_19
);
W_reg_59_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x11_out_1,
   R => '0',
   Q => W_reg_59_1
);
W_reg_59_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x11_out_20,
   R => '0',
   Q => W_reg_59_20
);
W_reg_59_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x11_out_21,
   R => '0',
   Q => W_reg_59_21
);
W_reg_59_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x11_out_22,
   R => '0',
   Q => W_reg_59_22
);
W_reg_59_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x11_out_23,
   R => '0',
   Q => W_reg_59_23
);
W_reg_59_23_i_1 : CARRY4
 port map (
   CI => W_reg_59_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_59_23_i_5_n_0,
   DI(1) => W_59_23_i_4_n_0,
   DI(2) => W_59_23_i_3_n_0,
   DI(3) => W_59_23_i_2_n_0,
   S(0) => W_59_23_i_9_n_0,
   S(1) => W_59_23_i_8_n_0,
   S(2) => W_59_23_i_7_n_0,
   S(3) => W_59_23_i_6_n_0,
   CO(0) => W_reg_59_23_i_1_n_3,
   CO(1) => W_reg_59_23_i_1_n_2,
   CO(2) => W_reg_59_23_i_1_n_1,
   CO(3) => W_reg_59_23_i_1_n_0,
   O(0) => x11_out_20,
   O(1) => x11_out_21,
   O(2) => x11_out_22,
   O(3) => x11_out_23
);
W_reg_59_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x11_out_24,
   R => '0',
   Q => W_reg_59_24
);
W_reg_59_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x11_out_25,
   R => '0',
   Q => W_reg_59_25
);
W_reg_59_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x11_out_26,
   R => '0',
   Q => W_reg_59_26
);
W_reg_59_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x11_out_27,
   R => '0',
   Q => W_reg_59_27
);
W_reg_59_27_i_1 : CARRY4
 port map (
   CI => W_reg_59_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_59_27_i_5_n_0,
   DI(1) => W_59_27_i_4_n_0,
   DI(2) => W_59_27_i_3_n_0,
   DI(3) => W_59_27_i_2_n_0,
   S(0) => W_59_27_i_9_n_0,
   S(1) => W_59_27_i_8_n_0,
   S(2) => W_59_27_i_7_n_0,
   S(3) => W_59_27_i_6_n_0,
   CO(0) => W_reg_59_27_i_1_n_3,
   CO(1) => W_reg_59_27_i_1_n_2,
   CO(2) => W_reg_59_27_i_1_n_1,
   CO(3) => W_reg_59_27_i_1_n_0,
   O(0) => x11_out_24,
   O(1) => x11_out_25,
   O(2) => x11_out_26,
   O(3) => x11_out_27
);
W_reg_59_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x11_out_28,
   R => '0',
   Q => W_reg_59_28
);
W_reg_59_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x11_out_29,
   R => '0',
   Q => W_reg_59_29
);
W_reg_59_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x11_out_2,
   R => '0',
   Q => W_reg_59_2
);
W_reg_59_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x11_out_30,
   R => '0',
   Q => W_reg_59_30
);
W_reg_59_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x11_out_31,
   R => '0',
   Q => W_reg_59_31
);
W_reg_59_31_i_1 : CARRY4
 port map (
   CI => W_reg_59_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_59_31_i_4_n_0,
   DI(1) => W_59_31_i_3_n_0,
   DI(2) => W_59_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_59_31_i_8_n_0,
   S(1) => W_59_31_i_7_n_0,
   S(2) => W_59_31_i_6_n_0,
   S(3) => W_59_31_i_5_n_0,
   CO(0) => W_reg_59_31_i_1_n_3,
   CO(1) => W_reg_59_31_i_1_n_2,
   CO(2) => W_reg_59_31_i_1_n_1,
   CO(3) => NLW_W_reg_59_31_i_1_CO_UNCONNECTED_3,
   O(0) => x11_out_28,
   O(1) => x11_out_29,
   O(2) => x11_out_30,
   O(3) => x11_out_31
);
W_reg_59_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x11_out_3,
   R => '0',
   Q => W_reg_59_3
);
W_reg_59_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_59_3_i_5_n_0,
   DI(1) => W_59_3_i_4_n_0,
   DI(2) => W_59_3_i_3_n_0,
   DI(3) => W_59_3_i_2_n_0,
   S(0) => W_59_3_i_9_n_0,
   S(1) => W_59_3_i_8_n_0,
   S(2) => W_59_3_i_7_n_0,
   S(3) => W_59_3_i_6_n_0,
   CO(0) => W_reg_59_3_i_1_n_3,
   CO(1) => W_reg_59_3_i_1_n_2,
   CO(2) => W_reg_59_3_i_1_n_1,
   CO(3) => W_reg_59_3_i_1_n_0,
   O(0) => x11_out_0,
   O(1) => x11_out_1,
   O(2) => x11_out_2,
   O(3) => x11_out_3
);
W_reg_59_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x11_out_4,
   R => '0',
   Q => W_reg_59_4
);
W_reg_59_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x11_out_5,
   R => '0',
   Q => W_reg_59_5
);
W_reg_59_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x11_out_6,
   R => '0',
   Q => W_reg_59_6
);
W_reg_59_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x11_out_7,
   R => '0',
   Q => W_reg_59_7
);
W_reg_59_7_i_1 : CARRY4
 port map (
   CI => W_reg_59_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_59_7_i_5_n_0,
   DI(1) => W_59_7_i_4_n_0,
   DI(2) => W_59_7_i_3_n_0,
   DI(3) => W_59_7_i_2_n_0,
   S(0) => W_59_7_i_9_n_0,
   S(1) => W_59_7_i_8_n_0,
   S(2) => W_59_7_i_7_n_0,
   S(3) => W_59_7_i_6_n_0,
   CO(0) => W_reg_59_7_i_1_n_3,
   CO(1) => W_reg_59_7_i_1_n_2,
   CO(2) => W_reg_59_7_i_1_n_1,
   CO(3) => W_reg_59_7_i_1_n_0,
   O(0) => x11_out_4,
   O(1) => x11_out_5,
   O(2) => x11_out_6,
   O(3) => x11_out_7
);
W_reg_59_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x11_out_8,
   R => '0',
   Q => W_reg_59_8
);
W_reg_59_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x11_out_9,
   R => '0',
   Q => W_reg_59_9
);
W_reg_5_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_5_0,
   R => '0',
   Q => W_reg_5_0
);
W_reg_5_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_5_10,
   R => '0',
   Q => W_reg_5_10
);
W_reg_5_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_5_11,
   R => '0',
   Q => W_reg_5_11
);
W_reg_5_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_5_12,
   R => '0',
   Q => W_reg_5_12
);
W_reg_5_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_5_13,
   R => '0',
   Q => W_reg_5_13
);
W_reg_5_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_5_14,
   R => '0',
   Q => W_reg_5_14
);
W_reg_5_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_5_15,
   R => '0',
   Q => W_reg_5_15
);
W_reg_5_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_5_16,
   R => '0',
   Q => W_reg_5_16
);
W_reg_5_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_5_17,
   R => '0',
   Q => W_reg_5_17
);
W_reg_5_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_5_18,
   R => '0',
   Q => W_reg_5_18
);
W_reg_5_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_5_19,
   R => '0',
   Q => W_reg_5_19
);
W_reg_5_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_5_1,
   R => '0',
   Q => W_reg_5_1
);
W_reg_5_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_5_20,
   R => '0',
   Q => W_reg_5_20
);
W_reg_5_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_5_21,
   R => '0',
   Q => W_reg_5_21
);
W_reg_5_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_5_22,
   R => '0',
   Q => W_reg_5_22
);
W_reg_5_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_5_23,
   R => '0',
   Q => W_reg_5_23
);
W_reg_5_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_5_24,
   R => '0',
   Q => W_reg_5_24
);
W_reg_5_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_5_25,
   R => '0',
   Q => W_reg_5_25
);
W_reg_5_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_5_26,
   R => '0',
   Q => W_reg_5_26
);
W_reg_5_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_5_27,
   R => '0',
   Q => W_reg_5_27
);
W_reg_5_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_5_28,
   R => '0',
   Q => W_reg_5_28
);
W_reg_5_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_5_29,
   R => '0',
   Q => W_reg_5_29
);
W_reg_5_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_5_2,
   R => '0',
   Q => W_reg_5_2
);
W_reg_5_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_5_30,
   R => '0',
   Q => W_reg_5_30
);
W_reg_5_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_5_31,
   R => '0',
   Q => W_reg_5_31
);
W_reg_5_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_5_3,
   R => '0',
   Q => W_reg_5_3
);
W_reg_5_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_5_4,
   R => '0',
   Q => W_reg_5_4
);
W_reg_5_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_5_5,
   R => '0',
   Q => W_reg_5_5
);
W_reg_5_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_5_6,
   R => '0',
   Q => W_reg_5_6
);
W_reg_5_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_5_7,
   R => '0',
   Q => W_reg_5_7
);
W_reg_5_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_5_8,
   R => '0',
   Q => W_reg_5_8
);
W_reg_5_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_5_9,
   R => '0',
   Q => W_reg_5_9
);
W_reg_60_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x8_out_0,
   R => '0',
   Q => W_reg_60_0
);
W_reg_60_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x8_out_10,
   R => '0',
   Q => W_reg_60_10
);
W_reg_60_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x8_out_11,
   R => '0',
   Q => W_reg_60_11
);
W_reg_60_11_i_1 : CARRY4
 port map (
   CI => W_reg_60_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_60_11_i_5_n_0,
   DI(1) => W_60_11_i_4_n_0,
   DI(2) => W_60_11_i_3_n_0,
   DI(3) => W_60_11_i_2_n_0,
   S(0) => W_60_11_i_9_n_0,
   S(1) => W_60_11_i_8_n_0,
   S(2) => W_60_11_i_7_n_0,
   S(3) => W_60_11_i_6_n_0,
   CO(0) => W_reg_60_11_i_1_n_3,
   CO(1) => W_reg_60_11_i_1_n_2,
   CO(2) => W_reg_60_11_i_1_n_1,
   CO(3) => W_reg_60_11_i_1_n_0,
   O(0) => x8_out_8,
   O(1) => x8_out_9,
   O(2) => x8_out_10,
   O(3) => x8_out_11
);
W_reg_60_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x8_out_12,
   R => '0',
   Q => W_reg_60_12
);
W_reg_60_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x8_out_13,
   R => '0',
   Q => W_reg_60_13
);
W_reg_60_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x8_out_14,
   R => '0',
   Q => W_reg_60_14
);
W_reg_60_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x8_out_15,
   R => '0',
   Q => W_reg_60_15
);
W_reg_60_15_i_1 : CARRY4
 port map (
   CI => W_reg_60_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_60_15_i_5_n_0,
   DI(1) => W_60_15_i_4_n_0,
   DI(2) => W_60_15_i_3_n_0,
   DI(3) => W_60_15_i_2_n_0,
   S(0) => W_60_15_i_9_n_0,
   S(1) => W_60_15_i_8_n_0,
   S(2) => W_60_15_i_7_n_0,
   S(3) => W_60_15_i_6_n_0,
   CO(0) => W_reg_60_15_i_1_n_3,
   CO(1) => W_reg_60_15_i_1_n_2,
   CO(2) => W_reg_60_15_i_1_n_1,
   CO(3) => W_reg_60_15_i_1_n_0,
   O(0) => x8_out_12,
   O(1) => x8_out_13,
   O(2) => x8_out_14,
   O(3) => x8_out_15
);
W_reg_60_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x8_out_16,
   R => '0',
   Q => W_reg_60_16
);
W_reg_60_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x8_out_17,
   R => '0',
   Q => W_reg_60_17
);
W_reg_60_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x8_out_18,
   R => '0',
   Q => W_reg_60_18
);
W_reg_60_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x8_out_19,
   R => '0',
   Q => W_reg_60_19
);
W_reg_60_19_i_1 : CARRY4
 port map (
   CI => W_reg_60_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_60_19_i_5_n_0,
   DI(1) => W_60_19_i_4_n_0,
   DI(2) => W_60_19_i_3_n_0,
   DI(3) => W_60_19_i_2_n_0,
   S(0) => W_60_19_i_9_n_0,
   S(1) => W_60_19_i_8_n_0,
   S(2) => W_60_19_i_7_n_0,
   S(3) => W_60_19_i_6_n_0,
   CO(0) => W_reg_60_19_i_1_n_3,
   CO(1) => W_reg_60_19_i_1_n_2,
   CO(2) => W_reg_60_19_i_1_n_1,
   CO(3) => W_reg_60_19_i_1_n_0,
   O(0) => x8_out_16,
   O(1) => x8_out_17,
   O(2) => x8_out_18,
   O(3) => x8_out_19
);
W_reg_60_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x8_out_1,
   R => '0',
   Q => W_reg_60_1
);
W_reg_60_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x8_out_20,
   R => '0',
   Q => W_reg_60_20
);
W_reg_60_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x8_out_21,
   R => '0',
   Q => W_reg_60_21
);
W_reg_60_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x8_out_22,
   R => '0',
   Q => W_reg_60_22
);
W_reg_60_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x8_out_23,
   R => '0',
   Q => W_reg_60_23
);
W_reg_60_23_i_1 : CARRY4
 port map (
   CI => W_reg_60_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_60_23_i_5_n_0,
   DI(1) => W_60_23_i_4_n_0,
   DI(2) => W_60_23_i_3_n_0,
   DI(3) => W_60_23_i_2_n_0,
   S(0) => W_60_23_i_9_n_0,
   S(1) => W_60_23_i_8_n_0,
   S(2) => W_60_23_i_7_n_0,
   S(3) => W_60_23_i_6_n_0,
   CO(0) => W_reg_60_23_i_1_n_3,
   CO(1) => W_reg_60_23_i_1_n_2,
   CO(2) => W_reg_60_23_i_1_n_1,
   CO(3) => W_reg_60_23_i_1_n_0,
   O(0) => x8_out_20,
   O(1) => x8_out_21,
   O(2) => x8_out_22,
   O(3) => x8_out_23
);
W_reg_60_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x8_out_24,
   R => '0',
   Q => W_reg_60_24
);
W_reg_60_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x8_out_25,
   R => '0',
   Q => W_reg_60_25
);
W_reg_60_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x8_out_26,
   R => '0',
   Q => W_reg_60_26
);
W_reg_60_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x8_out_27,
   R => '0',
   Q => W_reg_60_27
);
W_reg_60_27_i_1 : CARRY4
 port map (
   CI => W_reg_60_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_60_27_i_5_n_0,
   DI(1) => W_60_27_i_4_n_0,
   DI(2) => W_60_27_i_3_n_0,
   DI(3) => W_60_27_i_2_n_0,
   S(0) => W_60_27_i_9_n_0,
   S(1) => W_60_27_i_8_n_0,
   S(2) => W_60_27_i_7_n_0,
   S(3) => W_60_27_i_6_n_0,
   CO(0) => W_reg_60_27_i_1_n_3,
   CO(1) => W_reg_60_27_i_1_n_2,
   CO(2) => W_reg_60_27_i_1_n_1,
   CO(3) => W_reg_60_27_i_1_n_0,
   O(0) => x8_out_24,
   O(1) => x8_out_25,
   O(2) => x8_out_26,
   O(3) => x8_out_27
);
W_reg_60_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x8_out_28,
   R => '0',
   Q => W_reg_60_28
);
W_reg_60_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x8_out_29,
   R => '0',
   Q => W_reg_60_29
);
W_reg_60_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x8_out_2,
   R => '0',
   Q => W_reg_60_2
);
W_reg_60_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x8_out_30,
   R => '0',
   Q => W_reg_60_30
);
W_reg_60_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x8_out_31,
   R => '0',
   Q => W_reg_60_31
);
W_reg_60_31_i_1 : CARRY4
 port map (
   CI => W_reg_60_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_60_31_i_4_n_0,
   DI(1) => W_60_31_i_3_n_0,
   DI(2) => W_60_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_60_31_i_8_n_0,
   S(1) => W_60_31_i_7_n_0,
   S(2) => W_60_31_i_6_n_0,
   S(3) => W_60_31_i_5_n_0,
   CO(0) => W_reg_60_31_i_1_n_3,
   CO(1) => W_reg_60_31_i_1_n_2,
   CO(2) => W_reg_60_31_i_1_n_1,
   CO(3) => NLW_W_reg_60_31_i_1_CO_UNCONNECTED_3,
   O(0) => x8_out_28,
   O(1) => x8_out_29,
   O(2) => x8_out_30,
   O(3) => x8_out_31
);
W_reg_60_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x8_out_3,
   R => '0',
   Q => W_reg_60_3
);
W_reg_60_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_60_3_i_5_n_0,
   DI(1) => W_60_3_i_4_n_0,
   DI(2) => W_60_3_i_3_n_0,
   DI(3) => W_60_3_i_2_n_0,
   S(0) => W_60_3_i_9_n_0,
   S(1) => W_60_3_i_8_n_0,
   S(2) => W_60_3_i_7_n_0,
   S(3) => W_60_3_i_6_n_0,
   CO(0) => W_reg_60_3_i_1_n_3,
   CO(1) => W_reg_60_3_i_1_n_2,
   CO(2) => W_reg_60_3_i_1_n_1,
   CO(3) => W_reg_60_3_i_1_n_0,
   O(0) => x8_out_0,
   O(1) => x8_out_1,
   O(2) => x8_out_2,
   O(3) => x8_out_3
);
W_reg_60_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x8_out_4,
   R => '0',
   Q => W_reg_60_4
);
W_reg_60_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x8_out_5,
   R => '0',
   Q => W_reg_60_5
);
W_reg_60_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x8_out_6,
   R => '0',
   Q => W_reg_60_6
);
W_reg_60_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x8_out_7,
   R => '0',
   Q => W_reg_60_7
);
W_reg_60_7_i_1 : CARRY4
 port map (
   CI => W_reg_60_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_60_7_i_5_n_0,
   DI(1) => W_60_7_i_4_n_0,
   DI(2) => W_60_7_i_3_n_0,
   DI(3) => W_60_7_i_2_n_0,
   S(0) => W_60_7_i_9_n_0,
   S(1) => W_60_7_i_8_n_0,
   S(2) => W_60_7_i_7_n_0,
   S(3) => W_60_7_i_6_n_0,
   CO(0) => W_reg_60_7_i_1_n_3,
   CO(1) => W_reg_60_7_i_1_n_2,
   CO(2) => W_reg_60_7_i_1_n_1,
   CO(3) => W_reg_60_7_i_1_n_0,
   O(0) => x8_out_4,
   O(1) => x8_out_5,
   O(2) => x8_out_6,
   O(3) => x8_out_7
);
W_reg_60_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x8_out_8,
   R => '0',
   Q => W_reg_60_8
);
W_reg_60_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x8_out_9,
   R => '0',
   Q => W_reg_60_9
);
W_reg_61_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x_0,
   R => '0',
   Q => W_reg_61_0
);
W_reg_61_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x_10,
   R => '0',
   Q => W_reg_61_10
);
W_reg_61_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x_11,
   R => '0',
   Q => W_reg_61_11
);
W_reg_61_11_i_1 : CARRY4
 port map (
   CI => W_reg_61_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_61_11_i_5_n_0,
   DI(1) => W_61_11_i_4_n_0,
   DI(2) => W_61_11_i_3_n_0,
   DI(3) => W_61_11_i_2_n_0,
   S(0) => W_61_11_i_9_n_0,
   S(1) => W_61_11_i_8_n_0,
   S(2) => W_61_11_i_7_n_0,
   S(3) => W_61_11_i_6_n_0,
   CO(0) => W_reg_61_11_i_1_n_3,
   CO(1) => W_reg_61_11_i_1_n_2,
   CO(2) => W_reg_61_11_i_1_n_1,
   CO(3) => W_reg_61_11_i_1_n_0,
   O(0) => x_8,
   O(1) => x_9,
   O(2) => x_10,
   O(3) => x_11
);
W_reg_61_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x_12,
   R => '0',
   Q => W_reg_61_12
);
W_reg_61_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x_13,
   R => '0',
   Q => W_reg_61_13
);
W_reg_61_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x_14,
   R => '0',
   Q => W_reg_61_14
);
W_reg_61_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x_15,
   R => '0',
   Q => W_reg_61_15
);
W_reg_61_15_i_1 : CARRY4
 port map (
   CI => W_reg_61_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_61_15_i_5_n_0,
   DI(1) => W_61_15_i_4_n_0,
   DI(2) => W_61_15_i_3_n_0,
   DI(3) => W_61_15_i_2_n_0,
   S(0) => W_61_15_i_9_n_0,
   S(1) => W_61_15_i_8_n_0,
   S(2) => W_61_15_i_7_n_0,
   S(3) => W_61_15_i_6_n_0,
   CO(0) => W_reg_61_15_i_1_n_3,
   CO(1) => W_reg_61_15_i_1_n_2,
   CO(2) => W_reg_61_15_i_1_n_1,
   CO(3) => W_reg_61_15_i_1_n_0,
   O(0) => x_12,
   O(1) => x_13,
   O(2) => x_14,
   O(3) => x_15
);
W_reg_61_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x_16,
   R => '0',
   Q => W_reg_61_16
);
W_reg_61_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x_17,
   R => '0',
   Q => W_reg_61_17
);
W_reg_61_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x_18,
   R => '0',
   Q => W_reg_61_18
);
W_reg_61_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x_19,
   R => '0',
   Q => W_reg_61_19
);
W_reg_61_19_i_1 : CARRY4
 port map (
   CI => W_reg_61_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_61_19_i_5_n_0,
   DI(1) => W_61_19_i_4_n_0,
   DI(2) => W_61_19_i_3_n_0,
   DI(3) => W_61_19_i_2_n_0,
   S(0) => W_61_19_i_9_n_0,
   S(1) => W_61_19_i_8_n_0,
   S(2) => W_61_19_i_7_n_0,
   S(3) => W_61_19_i_6_n_0,
   CO(0) => W_reg_61_19_i_1_n_3,
   CO(1) => W_reg_61_19_i_1_n_2,
   CO(2) => W_reg_61_19_i_1_n_1,
   CO(3) => W_reg_61_19_i_1_n_0,
   O(0) => x_16,
   O(1) => x_17,
   O(2) => x_18,
   O(3) => x_19
);
W_reg_61_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x_1,
   R => '0',
   Q => W_reg_61_1
);
W_reg_61_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x_20,
   R => '0',
   Q => W_reg_61_20
);
W_reg_61_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x_21,
   R => '0',
   Q => W_reg_61_21
);
W_reg_61_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x_22,
   R => '0',
   Q => W_reg_61_22
);
W_reg_61_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x_23,
   R => '0',
   Q => W_reg_61_23
);
W_reg_61_23_i_1 : CARRY4
 port map (
   CI => W_reg_61_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_61_23_i_5_n_0,
   DI(1) => W_61_23_i_4_n_0,
   DI(2) => W_61_23_i_3_n_0,
   DI(3) => W_61_23_i_2_n_0,
   S(0) => W_61_23_i_9_n_0,
   S(1) => W_61_23_i_8_n_0,
   S(2) => W_61_23_i_7_n_0,
   S(3) => W_61_23_i_6_n_0,
   CO(0) => W_reg_61_23_i_1_n_3,
   CO(1) => W_reg_61_23_i_1_n_2,
   CO(2) => W_reg_61_23_i_1_n_1,
   CO(3) => W_reg_61_23_i_1_n_0,
   O(0) => x_20,
   O(1) => x_21,
   O(2) => x_22,
   O(3) => x_23
);
W_reg_61_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x_24,
   R => '0',
   Q => W_reg_61_24
);
W_reg_61_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x_25,
   R => '0',
   Q => W_reg_61_25
);
W_reg_61_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x_26,
   R => '0',
   Q => W_reg_61_26
);
W_reg_61_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x_27,
   R => '0',
   Q => W_reg_61_27
);
W_reg_61_27_i_1 : CARRY4
 port map (
   CI => W_reg_61_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_61_27_i_5_n_0,
   DI(1) => W_61_27_i_4_n_0,
   DI(2) => W_61_27_i_3_n_0,
   DI(3) => W_61_27_i_2_n_0,
   S(0) => W_61_27_i_9_n_0,
   S(1) => W_61_27_i_8_n_0,
   S(2) => W_61_27_i_7_n_0,
   S(3) => W_61_27_i_6_n_0,
   CO(0) => W_reg_61_27_i_1_n_3,
   CO(1) => W_reg_61_27_i_1_n_2,
   CO(2) => W_reg_61_27_i_1_n_1,
   CO(3) => W_reg_61_27_i_1_n_0,
   O(0) => x_24,
   O(1) => x_25,
   O(2) => x_26,
   O(3) => x_27
);
W_reg_61_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x_28,
   R => '0',
   Q => W_reg_61_28
);
W_reg_61_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x_29,
   R => '0',
   Q => W_reg_61_29
);
W_reg_61_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x_2,
   R => '0',
   Q => W_reg_61_2
);
W_reg_61_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x_30,
   R => '0',
   Q => W_reg_61_30
);
W_reg_61_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x_31,
   R => '0',
   Q => W_reg_61_31
);
W_reg_61_31_i_1 : CARRY4
 port map (
   CI => W_reg_61_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_61_31_i_4_n_0,
   DI(1) => W_61_31_i_3_n_0,
   DI(2) => W_61_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_61_31_i_8_n_0,
   S(1) => W_61_31_i_7_n_0,
   S(2) => W_61_31_i_6_n_0,
   S(3) => W_61_31_i_5_n_0,
   CO(0) => W_reg_61_31_i_1_n_3,
   CO(1) => W_reg_61_31_i_1_n_2,
   CO(2) => W_reg_61_31_i_1_n_1,
   CO(3) => NLW_W_reg_61_31_i_1_CO_UNCONNECTED_3,
   O(0) => x_28,
   O(1) => x_29,
   O(2) => x_30,
   O(3) => x_31
);
W_reg_61_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x_3,
   R => '0',
   Q => W_reg_61_3
);
W_reg_61_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_61_3_i_5_n_0,
   DI(1) => W_61_3_i_4_n_0,
   DI(2) => W_61_3_i_3_n_0,
   DI(3) => W_61_3_i_2_n_0,
   S(0) => W_61_3_i_9_n_0,
   S(1) => W_61_3_i_8_n_0,
   S(2) => W_61_3_i_7_n_0,
   S(3) => W_61_3_i_6_n_0,
   CO(0) => W_reg_61_3_i_1_n_3,
   CO(1) => W_reg_61_3_i_1_n_2,
   CO(2) => W_reg_61_3_i_1_n_1,
   CO(3) => W_reg_61_3_i_1_n_0,
   O(0) => x_0,
   O(1) => x_1,
   O(2) => x_2,
   O(3) => x_3
);
W_reg_61_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x_4,
   R => '0',
   Q => W_reg_61_4
);
W_reg_61_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x_5,
   R => '0',
   Q => W_reg_61_5
);
W_reg_61_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x_6,
   R => '0',
   Q => W_reg_61_6
);
W_reg_61_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x_7,
   R => '0',
   Q => W_reg_61_7
);
W_reg_61_7_i_1 : CARRY4
 port map (
   CI => W_reg_61_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_61_7_i_5_n_0,
   DI(1) => W_61_7_i_4_n_0,
   DI(2) => W_61_7_i_3_n_0,
   DI(3) => W_61_7_i_2_n_0,
   S(0) => W_61_7_i_9_n_0,
   S(1) => W_61_7_i_8_n_0,
   S(2) => W_61_7_i_7_n_0,
   S(3) => W_61_7_i_6_n_0,
   CO(0) => W_reg_61_7_i_1_n_3,
   CO(1) => W_reg_61_7_i_1_n_2,
   CO(2) => W_reg_61_7_i_1_n_1,
   CO(3) => W_reg_61_7_i_1_n_0,
   O(0) => x_4,
   O(1) => x_5,
   O(2) => x_6,
   O(3) => x_7
);
W_reg_61_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x_8,
   R => '0',
   Q => W_reg_61_8
);
W_reg_61_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => x_9,
   R => '0',
   Q => W_reg_61_9
);
W_reg_62_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_62_0,
   R => '0',
   Q => W_reg_62_0
);
W_reg_62_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_62_10,
   R => '0',
   Q => W_reg_62_10
);
W_reg_62_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_62_11,
   R => '0',
   Q => W_reg_62_11
);
W_reg_62_11_i_1 : CARRY4
 port map (
   CI => W_reg_62_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_62_11_i_5_n_0,
   DI(1) => W_62_11_i_4_n_0,
   DI(2) => W_62_11_i_3_n_0,
   DI(3) => W_62_11_i_2_n_0,
   S(0) => W_62_11_i_9_n_0,
   S(1) => W_62_11_i_8_n_0,
   S(2) => W_62_11_i_7_n_0,
   S(3) => W_62_11_i_6_n_0,
   CO(0) => W_reg_62_11_i_1_n_3,
   CO(1) => W_reg_62_11_i_1_n_2,
   CO(2) => W_reg_62_11_i_1_n_1,
   CO(3) => W_reg_62_11_i_1_n_0,
   O(0) => W_INT_62_8,
   O(1) => W_INT_62_9,
   O(2) => W_INT_62_10,
   O(3) => W_INT_62_11
);
W_reg_62_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_62_12,
   R => '0',
   Q => W_reg_62_12
);
W_reg_62_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_62_13,
   R => '0',
   Q => W_reg_62_13
);
W_reg_62_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_62_14,
   R => '0',
   Q => W_reg_62_14
);
W_reg_62_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_62_15,
   R => '0',
   Q => W_reg_62_15
);
W_reg_62_15_i_1 : CARRY4
 port map (
   CI => W_reg_62_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_62_15_i_5_n_0,
   DI(1) => W_62_15_i_4_n_0,
   DI(2) => W_62_15_i_3_n_0,
   DI(3) => W_62_15_i_2_n_0,
   S(0) => W_62_15_i_9_n_0,
   S(1) => W_62_15_i_8_n_0,
   S(2) => W_62_15_i_7_n_0,
   S(3) => W_62_15_i_6_n_0,
   CO(0) => W_reg_62_15_i_1_n_3,
   CO(1) => W_reg_62_15_i_1_n_2,
   CO(2) => W_reg_62_15_i_1_n_1,
   CO(3) => W_reg_62_15_i_1_n_0,
   O(0) => W_INT_62_12,
   O(1) => W_INT_62_13,
   O(2) => W_INT_62_14,
   O(3) => W_INT_62_15
);
W_reg_62_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_62_16,
   R => '0',
   Q => W_reg_62_16
);
W_reg_62_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_62_17,
   R => '0',
   Q => W_reg_62_17
);
W_reg_62_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_62_18,
   R => '0',
   Q => W_reg_62_18
);
W_reg_62_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_62_19,
   R => '0',
   Q => W_reg_62_19
);
W_reg_62_19_i_1 : CARRY4
 port map (
   CI => W_reg_62_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_62_19_i_5_n_0,
   DI(1) => W_62_19_i_4_n_0,
   DI(2) => W_62_19_i_3_n_0,
   DI(3) => W_62_19_i_2_n_0,
   S(0) => W_62_19_i_9_n_0,
   S(1) => W_62_19_i_8_n_0,
   S(2) => W_62_19_i_7_n_0,
   S(3) => W_62_19_i_6_n_0,
   CO(0) => W_reg_62_19_i_1_n_3,
   CO(1) => W_reg_62_19_i_1_n_2,
   CO(2) => W_reg_62_19_i_1_n_1,
   CO(3) => W_reg_62_19_i_1_n_0,
   O(0) => W_INT_62_16,
   O(1) => W_INT_62_17,
   O(2) => W_INT_62_18,
   O(3) => W_INT_62_19
);
W_reg_62_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_62_1,
   R => '0',
   Q => W_reg_62_1
);
W_reg_62_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_62_20,
   R => '0',
   Q => W_reg_62_20
);
W_reg_62_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_62_21,
   R => '0',
   Q => W_reg_62_21
);
W_reg_62_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_62_22,
   R => '0',
   Q => W_reg_62_22
);
W_reg_62_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_62_23,
   R => '0',
   Q => W_reg_62_23
);
W_reg_62_23_i_1 : CARRY4
 port map (
   CI => W_reg_62_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_62_23_i_5_n_0,
   DI(1) => W_62_23_i_4_n_0,
   DI(2) => W_62_23_i_3_n_0,
   DI(3) => W_62_23_i_2_n_0,
   S(0) => W_62_23_i_9_n_0,
   S(1) => W_62_23_i_8_n_0,
   S(2) => W_62_23_i_7_n_0,
   S(3) => W_62_23_i_6_n_0,
   CO(0) => W_reg_62_23_i_1_n_3,
   CO(1) => W_reg_62_23_i_1_n_2,
   CO(2) => W_reg_62_23_i_1_n_1,
   CO(3) => W_reg_62_23_i_1_n_0,
   O(0) => W_INT_62_20,
   O(1) => W_INT_62_21,
   O(2) => W_INT_62_22,
   O(3) => W_INT_62_23
);
W_reg_62_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_62_24,
   R => '0',
   Q => W_reg_62_24
);
W_reg_62_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_62_25,
   R => '0',
   Q => W_reg_62_25
);
W_reg_62_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_62_26,
   R => '0',
   Q => W_reg_62_26
);
W_reg_62_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_62_27,
   R => '0',
   Q => W_reg_62_27
);
W_reg_62_27_i_1 : CARRY4
 port map (
   CI => W_reg_62_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_62_27_i_5_n_0,
   DI(1) => W_62_27_i_4_n_0,
   DI(2) => W_62_27_i_3_n_0,
   DI(3) => W_62_27_i_2_n_0,
   S(0) => W_62_27_i_9_n_0,
   S(1) => W_62_27_i_8_n_0,
   S(2) => W_62_27_i_7_n_0,
   S(3) => W_62_27_i_6_n_0,
   CO(0) => W_reg_62_27_i_1_n_3,
   CO(1) => W_reg_62_27_i_1_n_2,
   CO(2) => W_reg_62_27_i_1_n_1,
   CO(3) => W_reg_62_27_i_1_n_0,
   O(0) => W_INT_62_24,
   O(1) => W_INT_62_25,
   O(2) => W_INT_62_26,
   O(3) => W_INT_62_27
);
W_reg_62_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_62_28,
   R => '0',
   Q => W_reg_62_28
);
W_reg_62_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_62_29,
   R => '0',
   Q => W_reg_62_29
);
W_reg_62_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_62_2,
   R => '0',
   Q => W_reg_62_2
);
W_reg_62_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_62_30,
   R => '0',
   Q => W_reg_62_30
);
W_reg_62_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_62_31,
   R => '0',
   Q => W_reg_62_31
);
W_reg_62_31_i_1 : CARRY4
 port map (
   CI => W_reg_62_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_62_31_i_4_n_0,
   DI(1) => W_62_31_i_3_n_0,
   DI(2) => W_62_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_62_31_i_8_n_0,
   S(1) => W_62_31_i_7_n_0,
   S(2) => W_62_31_i_6_n_0,
   S(3) => W_62_31_i_5_n_0,
   CO(0) => W_reg_62_31_i_1_n_3,
   CO(1) => W_reg_62_31_i_1_n_2,
   CO(2) => W_reg_62_31_i_1_n_1,
   CO(3) => NLW_W_reg_62_31_i_1_CO_UNCONNECTED_3,
   O(0) => W_INT_62_28,
   O(1) => W_INT_62_29,
   O(2) => W_INT_62_30,
   O(3) => W_INT_62_31
);
W_reg_62_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_62_3,
   R => '0',
   Q => W_reg_62_3
);
W_reg_62_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_62_3_i_5_n_0,
   DI(1) => W_62_3_i_4_n_0,
   DI(2) => W_62_3_i_3_n_0,
   DI(3) => W_62_3_i_2_n_0,
   S(0) => W_62_3_i_9_n_0,
   S(1) => W_62_3_i_8_n_0,
   S(2) => W_62_3_i_7_n_0,
   S(3) => W_62_3_i_6_n_0,
   CO(0) => W_reg_62_3_i_1_n_3,
   CO(1) => W_reg_62_3_i_1_n_2,
   CO(2) => W_reg_62_3_i_1_n_1,
   CO(3) => W_reg_62_3_i_1_n_0,
   O(0) => W_INT_62_0,
   O(1) => W_INT_62_1,
   O(2) => W_INT_62_2,
   O(3) => W_INT_62_3
);
W_reg_62_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_62_4,
   R => '0',
   Q => W_reg_62_4
);
W_reg_62_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_62_5,
   R => '0',
   Q => W_reg_62_5
);
W_reg_62_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_62_6,
   R => '0',
   Q => W_reg_62_6
);
W_reg_62_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_62_7,
   R => '0',
   Q => W_reg_62_7
);
W_reg_62_7_i_1 : CARRY4
 port map (
   CI => W_reg_62_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_62_7_i_5_n_0,
   DI(1) => W_62_7_i_4_n_0,
   DI(2) => W_62_7_i_3_n_0,
   DI(3) => W_62_7_i_2_n_0,
   S(0) => W_62_7_i_9_n_0,
   S(1) => W_62_7_i_8_n_0,
   S(2) => W_62_7_i_7_n_0,
   S(3) => W_62_7_i_6_n_0,
   CO(0) => W_reg_62_7_i_1_n_3,
   CO(1) => W_reg_62_7_i_1_n_2,
   CO(2) => W_reg_62_7_i_1_n_1,
   CO(3) => W_reg_62_7_i_1_n_0,
   O(0) => W_INT_62_4,
   O(1) => W_INT_62_5,
   O(2) => W_INT_62_6,
   O(3) => W_INT_62_7
);
W_reg_62_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_62_8,
   R => '0',
   Q => W_reg_62_8
);
W_reg_62_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_62_9,
   R => '0',
   Q => W_reg_62_9
);
W_reg_63_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_63_0,
   R => '0',
   Q => W_reg_63_0
);
W_reg_63_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_63_10,
   R => '0',
   Q => W_reg_63_10
);
W_reg_63_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_63_11,
   R => '0',
   Q => W_reg_63_11
);
W_reg_63_11_i_1 : CARRY4
 port map (
   CI => W_reg_63_7_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_63_11_i_5_n_0,
   DI(1) => W_63_11_i_4_n_0,
   DI(2) => W_63_11_i_3_n_0,
   DI(3) => W_63_11_i_2_n_0,
   S(0) => W_63_11_i_9_n_0,
   S(1) => W_63_11_i_8_n_0,
   S(2) => W_63_11_i_7_n_0,
   S(3) => W_63_11_i_6_n_0,
   CO(0) => W_reg_63_11_i_1_n_3,
   CO(1) => W_reg_63_11_i_1_n_2,
   CO(2) => W_reg_63_11_i_1_n_1,
   CO(3) => W_reg_63_11_i_1_n_0,
   O(0) => W_INT_63_8,
   O(1) => W_INT_63_9,
   O(2) => W_INT_63_10,
   O(3) => W_INT_63_11
);
W_reg_63_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_63_12,
   R => '0',
   Q => W_reg_63_12
);
W_reg_63_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_63_13,
   R => '0',
   Q => W_reg_63_13
);
W_reg_63_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_63_14,
   R => '0',
   Q => W_reg_63_14
);
W_reg_63_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_63_15,
   R => '0',
   Q => W_reg_63_15
);
W_reg_63_15_i_1 : CARRY4
 port map (
   CI => W_reg_63_11_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_63_15_i_5_n_0,
   DI(1) => W_63_15_i_4_n_0,
   DI(2) => W_63_15_i_3_n_0,
   DI(3) => W_63_15_i_2_n_0,
   S(0) => W_63_15_i_9_n_0,
   S(1) => W_63_15_i_8_n_0,
   S(2) => W_63_15_i_7_n_0,
   S(3) => W_63_15_i_6_n_0,
   CO(0) => W_reg_63_15_i_1_n_3,
   CO(1) => W_reg_63_15_i_1_n_2,
   CO(2) => W_reg_63_15_i_1_n_1,
   CO(3) => W_reg_63_15_i_1_n_0,
   O(0) => W_INT_63_12,
   O(1) => W_INT_63_13,
   O(2) => W_INT_63_14,
   O(3) => W_INT_63_15
);
W_reg_63_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_63_16,
   R => '0',
   Q => W_reg_63_16
);
W_reg_63_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_63_17,
   R => '0',
   Q => W_reg_63_17
);
W_reg_63_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_63_18,
   R => '0',
   Q => W_reg_63_18
);
W_reg_63_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_63_19,
   R => '0',
   Q => W_reg_63_19
);
W_reg_63_19_i_1 : CARRY4
 port map (
   CI => W_reg_63_15_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_63_19_i_5_n_0,
   DI(1) => W_63_19_i_4_n_0,
   DI(2) => W_63_19_i_3_n_0,
   DI(3) => W_63_19_i_2_n_0,
   S(0) => W_63_19_i_9_n_0,
   S(1) => W_63_19_i_8_n_0,
   S(2) => W_63_19_i_7_n_0,
   S(3) => W_63_19_i_6_n_0,
   CO(0) => W_reg_63_19_i_1_n_3,
   CO(1) => W_reg_63_19_i_1_n_2,
   CO(2) => W_reg_63_19_i_1_n_1,
   CO(3) => W_reg_63_19_i_1_n_0,
   O(0) => W_INT_63_16,
   O(1) => W_INT_63_17,
   O(2) => W_INT_63_18,
   O(3) => W_INT_63_19
);
W_reg_63_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_63_1,
   R => '0',
   Q => W_reg_63_1
);
W_reg_63_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_63_20,
   R => '0',
   Q => W_reg_63_20
);
W_reg_63_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_63_21,
   R => '0',
   Q => W_reg_63_21
);
W_reg_63_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_63_22,
   R => '0',
   Q => W_reg_63_22
);
W_reg_63_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_63_23,
   R => '0',
   Q => W_reg_63_23
);
W_reg_63_23_i_1 : CARRY4
 port map (
   CI => W_reg_63_19_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_63_23_i_5_n_0,
   DI(1) => W_63_23_i_4_n_0,
   DI(2) => W_63_23_i_3_n_0,
   DI(3) => W_63_23_i_2_n_0,
   S(0) => W_63_23_i_9_n_0,
   S(1) => W_63_23_i_8_n_0,
   S(2) => W_63_23_i_7_n_0,
   S(3) => W_63_23_i_6_n_0,
   CO(0) => W_reg_63_23_i_1_n_3,
   CO(1) => W_reg_63_23_i_1_n_2,
   CO(2) => W_reg_63_23_i_1_n_1,
   CO(3) => W_reg_63_23_i_1_n_0,
   O(0) => W_INT_63_20,
   O(1) => W_INT_63_21,
   O(2) => W_INT_63_22,
   O(3) => W_INT_63_23
);
W_reg_63_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_63_24,
   R => '0',
   Q => W_reg_63_24
);
W_reg_63_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_63_25,
   R => '0',
   Q => W_reg_63_25
);
W_reg_63_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_63_26,
   R => '0',
   Q => W_reg_63_26
);
W_reg_63_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_63_27,
   R => '0',
   Q => W_reg_63_27
);
W_reg_63_27_i_1 : CARRY4
 port map (
   CI => W_reg_63_23_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_63_27_i_5_n_0,
   DI(1) => W_63_27_i_4_n_0,
   DI(2) => W_63_27_i_3_n_0,
   DI(3) => W_63_27_i_2_n_0,
   S(0) => W_63_27_i_9_n_0,
   S(1) => W_63_27_i_8_n_0,
   S(2) => W_63_27_i_7_n_0,
   S(3) => W_63_27_i_6_n_0,
   CO(0) => W_reg_63_27_i_1_n_3,
   CO(1) => W_reg_63_27_i_1_n_2,
   CO(2) => W_reg_63_27_i_1_n_1,
   CO(3) => W_reg_63_27_i_1_n_0,
   O(0) => W_INT_63_24,
   O(1) => W_INT_63_25,
   O(2) => W_INT_63_26,
   O(3) => W_INT_63_27
);
W_reg_63_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_63_28,
   R => '0',
   Q => W_reg_63_28
);
W_reg_63_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_63_29,
   R => '0',
   Q => W_reg_63_29
);
W_reg_63_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_63_2,
   R => '0',
   Q => W_reg_63_2
);
W_reg_63_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_63_30,
   R => '0',
   Q => W_reg_63_30
);
W_reg_63_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_63_31,
   R => '0',
   Q => W_reg_63_31
);
W_reg_63_31_i_1 : CARRY4
 port map (
   CI => W_reg_63_27_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_63_31_i_4_n_0,
   DI(1) => W_63_31_i_3_n_0,
   DI(2) => W_63_31_i_2_n_0,
   DI(3) => '0',
   S(0) => W_63_31_i_8_n_0,
   S(1) => W_63_31_i_7_n_0,
   S(2) => W_63_31_i_6_n_0,
   S(3) => W_63_31_i_5_n_0,
   CO(0) => W_reg_63_31_i_1_n_3,
   CO(1) => W_reg_63_31_i_1_n_2,
   CO(2) => W_reg_63_31_i_1_n_1,
   CO(3) => NLW_W_reg_63_31_i_1_CO_UNCONNECTED_3,
   O(0) => W_INT_63_28,
   O(1) => W_INT_63_29,
   O(2) => W_INT_63_30,
   O(3) => W_INT_63_31
);
W_reg_63_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_63_3,
   R => '0',
   Q => W_reg_63_3
);
W_reg_63_3_i_1 : CARRY4
 port map (
   CI => '0',
   CYINIT => '0',
   DI(0) => W_63_3_i_5_n_0,
   DI(1) => W_63_3_i_4_n_0,
   DI(2) => W_63_3_i_3_n_0,
   DI(3) => W_63_3_i_2_n_0,
   S(0) => W_63_3_i_9_n_0,
   S(1) => W_63_3_i_8_n_0,
   S(2) => W_63_3_i_7_n_0,
   S(3) => W_63_3_i_6_n_0,
   CO(0) => W_reg_63_3_i_1_n_3,
   CO(1) => W_reg_63_3_i_1_n_2,
   CO(2) => W_reg_63_3_i_1_n_1,
   CO(3) => W_reg_63_3_i_1_n_0,
   O(0) => W_INT_63_0,
   O(1) => W_INT_63_1,
   O(2) => W_INT_63_2,
   O(3) => W_INT_63_3
);
W_reg_63_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_63_4,
   R => '0',
   Q => W_reg_63_4
);
W_reg_63_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_63_5,
   R => '0',
   Q => W_reg_63_5
);
W_reg_63_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_63_6,
   R => '0',
   Q => W_reg_63_6
);
W_reg_63_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_63_7,
   R => '0',
   Q => W_reg_63_7
);
W_reg_63_7_i_1 : CARRY4
 port map (
   CI => W_reg_63_3_i_1_n_0,
   CYINIT => '0',
   DI(0) => W_63_7_i_5_n_0,
   DI(1) => W_63_7_i_4_n_0,
   DI(2) => W_63_7_i_3_n_0,
   DI(3) => W_63_7_i_2_n_0,
   S(0) => W_63_7_i_9_n_0,
   S(1) => W_63_7_i_8_n_0,
   S(2) => W_63_7_i_7_n_0,
   S(3) => W_63_7_i_6_n_0,
   CO(0) => W_reg_63_7_i_1_n_3,
   CO(1) => W_reg_63_7_i_1_n_2,
   CO(2) => W_reg_63_7_i_1_n_1,
   CO(3) => W_reg_63_7_i_1_n_0,
   O(0) => W_INT_63_4,
   O(1) => W_INT_63_5,
   O(2) => W_INT_63_6,
   O(3) => W_INT_63_7
);
W_reg_63_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_63_8,
   R => '0',
   Q => W_reg_63_8
);
W_reg_63_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_48_0,
   D => W_INT_63_9,
   R => '0',
   Q => W_reg_63_9
);
W_reg_6_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_6_0,
   R => '0',
   Q => W_reg_6_0
);
W_reg_6_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_6_10,
   R => '0',
   Q => W_reg_6_10
);
W_reg_6_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_6_11,
   R => '0',
   Q => W_reg_6_11
);
W_reg_6_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_6_12,
   R => '0',
   Q => W_reg_6_12
);
W_reg_6_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_6_13,
   R => '0',
   Q => W_reg_6_13
);
W_reg_6_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_6_14,
   R => '0',
   Q => W_reg_6_14
);
W_reg_6_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_6_15,
   R => '0',
   Q => W_reg_6_15
);
W_reg_6_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_6_16,
   R => '0',
   Q => W_reg_6_16
);
W_reg_6_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_6_17,
   R => '0',
   Q => W_reg_6_17
);
W_reg_6_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_6_18,
   R => '0',
   Q => W_reg_6_18
);
W_reg_6_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_6_19,
   R => '0',
   Q => W_reg_6_19
);
W_reg_6_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_6_1,
   R => '0',
   Q => W_reg_6_1
);
W_reg_6_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_6_20,
   R => '0',
   Q => W_reg_6_20
);
W_reg_6_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_6_21,
   R => '0',
   Q => W_reg_6_21
);
W_reg_6_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_6_22,
   R => '0',
   Q => W_reg_6_22
);
W_reg_6_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_6_23,
   R => '0',
   Q => W_reg_6_23
);
W_reg_6_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_6_24,
   R => '0',
   Q => W_reg_6_24
);
W_reg_6_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_6_25,
   R => '0',
   Q => W_reg_6_25
);
W_reg_6_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_6_26,
   R => '0',
   Q => W_reg_6_26
);
W_reg_6_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_6_27,
   R => '0',
   Q => W_reg_6_27
);
W_reg_6_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_6_28,
   R => '0',
   Q => W_reg_6_28
);
W_reg_6_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_6_29,
   R => '0',
   Q => W_reg_6_29
);
W_reg_6_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_6_2,
   R => '0',
   Q => W_reg_6_2
);
W_reg_6_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_6_30,
   R => '0',
   Q => W_reg_6_30
);
W_reg_6_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_6_31,
   R => '0',
   Q => W_reg_6_31
);
W_reg_6_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_6_3,
   R => '0',
   Q => W_reg_6_3
);
W_reg_6_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_6_4,
   R => '0',
   Q => W_reg_6_4
);
W_reg_6_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_6_5,
   R => '0',
   Q => W_reg_6_5
);
W_reg_6_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_6_6,
   R => '0',
   Q => W_reg_6_6
);
W_reg_6_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_6_7,
   R => '0',
   Q => W_reg_6_7
);
W_reg_6_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_6_8,
   R => '0',
   Q => W_reg_6_8
);
W_reg_6_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_6_9,
   R => '0',
   Q => W_reg_6_9
);
W_reg_7_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_7_0,
   R => '0',
   Q => W_reg_7_0
);
W_reg_7_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_7_10,
   R => '0',
   Q => W_reg_7_10
);
W_reg_7_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_7_11,
   R => '0',
   Q => W_reg_7_11
);
W_reg_7_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_7_12,
   R => '0',
   Q => W_reg_7_12
);
W_reg_7_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_7_13,
   R => '0',
   Q => W_reg_7_13
);
W_reg_7_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_7_14,
   R => '0',
   Q => W_reg_7_14
);
W_reg_7_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_7_15,
   R => '0',
   Q => W_reg_7_15
);
W_reg_7_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_7_16,
   R => '0',
   Q => W_reg_7_16
);
W_reg_7_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_7_17,
   R => '0',
   Q => W_reg_7_17
);
W_reg_7_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_7_18,
   R => '0',
   Q => W_reg_7_18
);
W_reg_7_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_7_19,
   R => '0',
   Q => W_reg_7_19
);
W_reg_7_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_7_1,
   R => '0',
   Q => W_reg_7_1
);
W_reg_7_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_7_20,
   R => '0',
   Q => W_reg_7_20
);
W_reg_7_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_7_21,
   R => '0',
   Q => W_reg_7_21
);
W_reg_7_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_7_22,
   R => '0',
   Q => W_reg_7_22
);
W_reg_7_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_7_23,
   R => '0',
   Q => W_reg_7_23
);
W_reg_7_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_7_24,
   R => '0',
   Q => W_reg_7_24
);
W_reg_7_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_7_25,
   R => '0',
   Q => W_reg_7_25
);
W_reg_7_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_7_26,
   R => '0',
   Q => W_reg_7_26
);
W_reg_7_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_7_27,
   R => '0',
   Q => W_reg_7_27
);
W_reg_7_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_7_28,
   R => '0',
   Q => W_reg_7_28
);
W_reg_7_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_7_29,
   R => '0',
   Q => W_reg_7_29
);
W_reg_7_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_7_2,
   R => '0',
   Q => W_reg_7_2
);
W_reg_7_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_7_30,
   R => '0',
   Q => W_reg_7_30
);
W_reg_7_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_7_31,
   R => '0',
   Q => W_reg_7_31
);
W_reg_7_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_7_3,
   R => '0',
   Q => W_reg_7_3
);
W_reg_7_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_7_4,
   R => '0',
   Q => W_reg_7_4
);
W_reg_7_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_7_5,
   R => '0',
   Q => W_reg_7_5
);
W_reg_7_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_7_6,
   R => '0',
   Q => W_reg_7_6
);
W_reg_7_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_7_7,
   R => '0',
   Q => W_reg_7_7
);
W_reg_7_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_7_8,
   R => '0',
   Q => W_reg_7_8
);
W_reg_7_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_7_9,
   R => '0',
   Q => W_reg_7_9
);
W_reg_8_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_8_0,
   R => '0',
   Q => W_reg_8_0
);
W_reg_8_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_8_10,
   R => '0',
   Q => W_reg_8_10
);
W_reg_8_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_8_11,
   R => '0',
   Q => W_reg_8_11
);
W_reg_8_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_8_12,
   R => '0',
   Q => W_reg_8_12
);
W_reg_8_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_8_13,
   R => '0',
   Q => W_reg_8_13
);
W_reg_8_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_8_14,
   R => '0',
   Q => W_reg_8_14
);
W_reg_8_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_8_15,
   R => '0',
   Q => W_reg_8_15
);
W_reg_8_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_8_16,
   R => '0',
   Q => W_reg_8_16
);
W_reg_8_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_8_17,
   R => '0',
   Q => W_reg_8_17
);
W_reg_8_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_8_18,
   R => '0',
   Q => W_reg_8_18
);
W_reg_8_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_8_19,
   R => '0',
   Q => W_reg_8_19
);
W_reg_8_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_8_1,
   R => '0',
   Q => W_reg_8_1
);
W_reg_8_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_8_20,
   R => '0',
   Q => W_reg_8_20
);
W_reg_8_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_8_21,
   R => '0',
   Q => W_reg_8_21
);
W_reg_8_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_8_22,
   R => '0',
   Q => W_reg_8_22
);
W_reg_8_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_8_23,
   R => '0',
   Q => W_reg_8_23
);
W_reg_8_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_8_24,
   R => '0',
   Q => W_reg_8_24
);
W_reg_8_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_8_25,
   R => '0',
   Q => W_reg_8_25
);
W_reg_8_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_8_26,
   R => '0',
   Q => W_reg_8_26
);
W_reg_8_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_8_27,
   R => '0',
   Q => W_reg_8_27
);
W_reg_8_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_8_28,
   R => '0',
   Q => W_reg_8_28
);
W_reg_8_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_8_29,
   R => '0',
   Q => W_reg_8_29
);
W_reg_8_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_8_2,
   R => '0',
   Q => W_reg_8_2
);
W_reg_8_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_8_30,
   R => '0',
   Q => W_reg_8_30
);
W_reg_8_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_8_31,
   R => '0',
   Q => W_reg_8_31
);
W_reg_8_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_8_3,
   R => '0',
   Q => W_reg_8_3
);
W_reg_8_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_8_4,
   R => '0',
   Q => W_reg_8_4
);
W_reg_8_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_8_5,
   R => '0',
   Q => W_reg_8_5
);
W_reg_8_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_8_6,
   R => '0',
   Q => W_reg_8_6
);
W_reg_8_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_8_7,
   R => '0',
   Q => W_reg_8_7
);
W_reg_8_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_8_8,
   R => '0',
   Q => W_reg_8_8
);
W_reg_8_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_8_9,
   R => '0',
   Q => W_reg_8_9
);
W_reg_9_0 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_9_0,
   R => '0',
   Q => W_reg_9_0
);
W_reg_9_10 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_9_10,
   R => '0',
   Q => W_reg_9_10
);
W_reg_9_11 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_9_11,
   R => '0',
   Q => W_reg_9_11
);
W_reg_9_12 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_9_12,
   R => '0',
   Q => W_reg_9_12
);
W_reg_9_13 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_9_13,
   R => '0',
   Q => W_reg_9_13
);
W_reg_9_14 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_9_14,
   R => '0',
   Q => W_reg_9_14
);
W_reg_9_15 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_9_15,
   R => '0',
   Q => W_reg_9_15
);
W_reg_9_16 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_9_16,
   R => '0',
   Q => W_reg_9_16
);
W_reg_9_17 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_9_17,
   R => '0',
   Q => W_reg_9_17
);
W_reg_9_18 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_9_18,
   R => '0',
   Q => W_reg_9_18
);
W_reg_9_19 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_9_19,
   R => '0',
   Q => W_reg_9_19
);
W_reg_9_1 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_9_1,
   R => '0',
   Q => W_reg_9_1
);
W_reg_9_20 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_9_20,
   R => '0',
   Q => W_reg_9_20
);
W_reg_9_21 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_9_21,
   R => '0',
   Q => W_reg_9_21
);
W_reg_9_22 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_9_22,
   R => '0',
   Q => W_reg_9_22
);
W_reg_9_23 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_9_23,
   R => '0',
   Q => W_reg_9_23
);
W_reg_9_24 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_9_24,
   R => '0',
   Q => W_reg_9_24
);
W_reg_9_25 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_9_25,
   R => '0',
   Q => W_reg_9_25
);
W_reg_9_26 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_9_26,
   R => '0',
   Q => W_reg_9_26
);
W_reg_9_27 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_9_27,
   R => '0',
   Q => W_reg_9_27
);
W_reg_9_28 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_9_28,
   R => '0',
   Q => W_reg_9_28
);
W_reg_9_29 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_9_29,
   R => '0',
   Q => W_reg_9_29
);
W_reg_9_2 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_9_2,
   R => '0',
   Q => W_reg_9_2
);
W_reg_9_30 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_9_30,
   R => '0',
   Q => W_reg_9_30
);
W_reg_9_31 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_9_31,
   R => '0',
   Q => W_reg_9_31
);
W_reg_9_3 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_9_3,
   R => '0',
   Q => W_reg_9_3
);
W_reg_9_4 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_9_4,
   R => '0',
   Q => W_reg_9_4
);
W_reg_9_5 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_9_5,
   R => '0',
   Q => W_reg_9_5
);
W_reg_9_6 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_9_6,
   R => '0',
   Q => W_reg_9_6
);
W_reg_9_7 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_9_7,
   R => '0',
   Q => W_reg_9_7
);
W_reg_9_8 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_9_8,
   R => '0',
   Q => W_reg_9_8
);
W_reg_9_9 : FDRE
  generic map(
   INIT => '0'
  )
 port map (
   C => clk_IBUF_BUFG,
   CE => W_reg_0_0,
   D => M_reg_9_9,
   R => '0',
   Q => W_reg_9_9
);
global_gnd : GND
 port map (
   G => '0'
);
global_vcc : VCC
 port map (
   P => '1'
);
end STRUCTURE;
