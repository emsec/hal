`timescale 1 ps/1 ps
module top(\simple_cpu_inst/alu_in2(1) ,\simple_cpu_inst/alu_in2(7) ,\simple_cpu_inst/alu_in2(12) ,\simple_cpu_inst/alu_in1_reg_n_0_[10] ,\simple_cpu_inst/alu_in1_reg_n_0_[0] ,\simple_cpu_inst/alu_in1_reg_n_0_[1] ,\simple_cpu_inst/alu_in2(10) ,\simple_cpu_inst/alu_in1_reg_n_0_[9] ,\simple_cpu_inst/alu_in2(20) ,\simple_cpu_inst/alu_in1_reg_n_0_[17] ,\simple_cpu_inst/alu_in1_reg_n_0_[22] ,\simple_cpu_inst/alu_in1_reg_n_0_[25] ,\simple_cpu_inst/alu_in2(18) ,\simple_cpu_inst/alu_in1_reg_n_0_[5] ,\simple_cpu_inst/alu_in2(24) ,\simple_cpu_inst/alu_in2(14) ,\simple_cpu_inst/alu_in1_reg_n_0_[8] ,\simple_cpu_inst/alu_in1_reg_n_0_[20] ,\simple_cpu_inst/alu_in1_reg_n_0_[12] ,\simple_cpu_inst/alu_in1_reg_n_0_[2] ,\simple_cpu_inst/alu_in2(0) ,\simple_cpu_inst/alu_in1_reg_n_0_[21] ,\simple_cpu_inst/alu_in2(19) ,\simple_cpu_inst/alu_in1_reg_n_0_[23] ,\simple_cpu_inst/alu_in1_reg_n_0_[6] ,\simple_cpu_inst/alu_in2(4) ,\simple_cpu_inst/alu_in1_reg_n_0_[18] ,\simple_cpu_inst/alu_in1_reg_n_0_[13] ,\simple_cpu_inst/alu_in1_reg_n_0_[19] ,\simple_cpu_inst/alu_in1_reg_n_0_[29] ,\simple_cpu_inst/alu_in2(23) ,\simple_cpu_inst/alu_in2(22) ,\simple_cpu_inst/alu_in2(31) ,\simple_cpu_inst/alu_in1_reg_n_0_[3] ,\simple_cpu_inst/alu_in2(28) ,\simple_cpu_inst/alu_in2(3) ,\simple_cpu_inst/alu_in1_reg_n_0_[24] ,\simple_cpu_inst/alu_in2(21) ,\simple_cpu_inst/alu_in2(27) ,\simple_cpu_inst/alu_in2(15) ,\simple_cpu_inst/alu_in2(2) ,\simple_cpu_inst/alu_in1_reg_n_0_[11] ,\simple_cpu_inst/alu_in1_reg_n_0_[7] ,\simple_cpu_inst/alu_in1_reg_n_0_[30] ,\simple_cpu_inst/alu_in1_reg_n_0_[28] ,\simple_cpu_inst/alu_in2(29) ,\simple_cpu_inst/alu_in1_reg_n_0_[14] ,\simple_cpu_inst/alu_in2(11) ,\simple_cpu_inst/alu_in1_reg_n_0_[4] ,\simple_cpu_inst/alu_in2(13) ,\simple_cpu_inst/alu_in2(25) ,\simple_cpu_inst/alu_in2(17) ,\simple_cpu_inst/alu_in1_reg_n_0_[15] ,\simple_cpu_inst/alu_in1_reg_n_0_[16] ,\simple_cpu_inst/alu_in2(9) ,\simple_cpu_inst/alu_in2(8) ,\simple_cpu_inst/alu_in2(6) ,\simple_cpu_inst/alu_in2(16) ,\simple_cpu_inst/alu_in1_reg_n_0_[31] ,\simple_cpu_inst/alu_in1_reg_n_0_[27] ,\simple_cpu_inst/alu_in1_reg_n_0_[26] ,\simple_cpu_inst/alu_in2(30) ,\simple_cpu_inst/alu_in2(5) ,\simple_cpu_inst/alu_in2(26) ,\simple_cpu_inst/alu_inst/data5 );
    input \simple_cpu_inst/alu_in2(1) ;
    input \simple_cpu_inst/alu_in2(7) ;
    input \simple_cpu_inst/alu_in2(12) ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[10] ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[0] ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[1] ;
    input \simple_cpu_inst/alu_in2(10) ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[9] ;
    input \simple_cpu_inst/alu_in2(20) ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[17] ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[22] ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[25] ;
    input \simple_cpu_inst/alu_in2(18) ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[5] ;
    input \simple_cpu_inst/alu_in2(24) ;
    input \simple_cpu_inst/alu_in2(14) ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[8] ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[20] ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[12] ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[2] ;
    input \simple_cpu_inst/alu_in2(0) ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[21] ;
    input \simple_cpu_inst/alu_in2(19) ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[23] ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[6] ;
    input \simple_cpu_inst/alu_in2(4) ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[18] ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[13] ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[19] ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[29] ;
    input \simple_cpu_inst/alu_in2(23) ;
    input \simple_cpu_inst/alu_in2(22) ;
    input \simple_cpu_inst/alu_in2(31) ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[3] ;
    input \simple_cpu_inst/alu_in2(28) ;
    input \simple_cpu_inst/alu_in2(3) ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[24] ;
    input \simple_cpu_inst/alu_in2(21) ;
    input \simple_cpu_inst/alu_in2(27) ;
    input \simple_cpu_inst/alu_in2(15) ;
    input \simple_cpu_inst/alu_in2(2) ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[11] ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[7] ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[30] ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[28] ;
    input \simple_cpu_inst/alu_in2(29) ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[14] ;
    input \simple_cpu_inst/alu_in2(11) ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[4] ;
    input \simple_cpu_inst/alu_in2(13) ;
    input \simple_cpu_inst/alu_in2(25) ;
    input \simple_cpu_inst/alu_in2(17) ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[15] ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[16] ;
    input \simple_cpu_inst/alu_in2(9) ;
    input \simple_cpu_inst/alu_in2(8) ;
    input \simple_cpu_inst/alu_in2(6) ;
    input \simple_cpu_inst/alu_in2(16) ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[31] ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[27] ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[26] ;
    input \simple_cpu_inst/alu_in2(30) ;
    input \simple_cpu_inst/alu_in2(5) ;
    input \simple_cpu_inst/alu_in2(26) ;
    output \simple_cpu_inst/alu_inst/data5 ;
    wire i__carry__1_i_2__1_n_0;
    wire \simple_cpu_inst/alu_inst/acc0_inferred__4/i__carry__0_n_3 ;
    wire i__carry__1_i_7_n_0;
    wire i__carry__2_i_4__1_n_0;
    wire i__carry__1_i_6_n_0;
    wire i__carry__1_i_1__1_n_0;
    wire \simple_cpu_inst/alu_inst/acc0_inferred__4/i__carry__1_n_3 ;
    wire i__carry__0_i_2__1_n_0;
    wire i__carry__0_i_1__1_n_0;
    wire i__carry__2_i_7_n_0;
    wire \simple_cpu_inst/alu_inst/acc0_inferred__4/i__carry_n_1 ;
    wire i__carry__2_i_1__2_n_0;
    wire i__carry__2_i_6_n_0;
    wire \simple_cpu_inst/alu_inst/acc0_inferred__4/i__carry__1_n_1 ;
    wire i__carry__1_i_3__1_n_0;
    wire i__carry__2_i_5_n_0;
    wire \simple_cpu_inst/alu_inst/acc0_inferred__4/i__carry__2_n_2 ;
    wire i__carry__0_i_7_n_0;
    wire i__carry__1_i_4__1_n_0;
    wire i__carry_i_8_n_0;
    wire i__carry_i_5_n_0;
    wire \simple_cpu_inst/alu_inst/acc0_inferred__4/i__carry__1_n_2 ;
    wire \simple_cpu_inst/alu_inst/acc0_inferred__4/i__carry__1_n_0 ;
    wire \simple_cpu_inst/alu_inst/acc0_inferred__4/i__carry_n_2 ;
    wire i__carry_i_7_n_0;
    wire i__carry__0_i_8_n_0;
    wire \simple_cpu_inst/alu_inst/acc0_inferred__4/i__carry__0_n_0 ;
    wire i__carry__2_i_2__1_n_0;
    wire i__carry__1_i_5_n_0;
    wire i__carry__2_i_8_n_0;
    wire i__carry_i_1__1_n_0;
    wire i__carry__1_i_8_n_0;
    wire \simple_cpu_inst/alu_inst/acc0_inferred__4/i__carry__0_n_1 ;
    wire \simple_cpu_inst/alu_inst/acc0_inferred__4/i__carry__2_n_3 ;
    wire \simple_cpu_inst/alu_inst/acc0_inferred__4/i__carry_n_0 ;
    wire \simple_cpu_inst/alu_inst/acc0_inferred__4/i__carry_n_3 ;
    wire i__carry_i_6_n_0;
    wire i__carry_i_2__1_n_0;
    wire i__carry_i_4_n_0;
    wire i__carry__0_i_3__1_n_0;
    wire i__carry__0_i_5_n_0;
    wire i__carry__0_i_6_n_0;
    wire i__carry_i_3__0_n_0;
    wire i__carry__2_i_3__1_n_0;
    wire \simple_cpu_inst/alu_inst/acc0_inferred__4/i__carry__0_n_2 ;
    wire i__carry__0_i_4__1_n_0;
    wire \simple_cpu_inst/alu_inst/acc0_inferred__4/i__carry__2_n_1 ;

    CARRY4 \simple_cpu_inst/alu_inst/acc0_inferred__4/i__carry__1  (
        .CI(\simple_cpu_inst/alu_inst/acc0_inferred__4/i__carry__0_n_0 ),
        .CYINIT(1'b0),
        .DI({
            i__carry__1_i_1__1_n_0,
            i__carry__1_i_2__1_n_0,
            i__carry__1_i_3__1_n_0,
            i__carry__1_i_4__1_n_0
        }),
        .S({
            i__carry__1_i_5_n_0,
            i__carry__1_i_6_n_0,
            i__carry__1_i_7_n_0,
            i__carry__1_i_8_n_0
        }),
        .CO({
            \simple_cpu_inst/alu_inst/acc0_inferred__4/i__carry__1_n_0 ,
            \simple_cpu_inst/alu_inst/acc0_inferred__4/i__carry__1_n_1 ,
            \simple_cpu_inst/alu_inst/acc0_inferred__4/i__carry__1_n_2 ,
            \simple_cpu_inst/alu_inst/acc0_inferred__4/i__carry__1_n_3 
        })
    );

    CARRY4 \simple_cpu_inst/alu_inst/acc0_inferred__4/i__carry__2  (
        .CI(\simple_cpu_inst/alu_inst/acc0_inferred__4/i__carry__1_n_0 ),
        .CYINIT(1'b0),
        .DI({
            i__carry__2_i_1__2_n_0,
            i__carry__2_i_2__1_n_0,
            i__carry__2_i_3__1_n_0,
            i__carry__2_i_4__1_n_0
        }),
        .S({
            i__carry__2_i_5_n_0,
            i__carry__2_i_6_n_0,
            i__carry__2_i_7_n_0,
            i__carry__2_i_8_n_0
        }),
        .CO({
            \simple_cpu_inst/alu_inst/data5 ,
            \simple_cpu_inst/alu_inst/acc0_inferred__4/i__carry__2_n_1 ,
            \simple_cpu_inst/alu_inst/acc0_inferred__4/i__carry__2_n_2 ,
            \simple_cpu_inst/alu_inst/acc0_inferred__4/i__carry__2_n_3 
        })
    );

    LUT4 #(
        .INIT(16'h9009)
    ) i__carry__1_i_8 (
        .I0(\simple_cpu_inst/alu_in2(17) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[17] ),
        .I2(\simple_cpu_inst/alu_in2(16) ),
        .I3(\simple_cpu_inst/alu_in1_reg_n_0_[16] ),
        .O(i__carry__1_i_8_n_0)
    );

    LUT4 #(
        .INIT(16'h44D4)
    ) i__carry__1_i_4__1 (
        .I0(\simple_cpu_inst/alu_in1_reg_n_0_[17] ),
        .I1(\simple_cpu_inst/alu_in2(17) ),
        .I2(\simple_cpu_inst/alu_in2(16) ),
        .I3(\simple_cpu_inst/alu_in1_reg_n_0_[16] ),
        .O(i__carry__1_i_4__1_n_0)
    );

    LUT4 #(
        .INIT(16'h9009)
    ) i__carry__2_i_8 (
        .I0(\simple_cpu_inst/alu_in2(25) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[25] ),
        .I2(\simple_cpu_inst/alu_in2(24) ),
        .I3(\simple_cpu_inst/alu_in1_reg_n_0_[24] ),
        .O(i__carry__2_i_8_n_0)
    );

    LUT4 #(
        .INIT(16'h9009)
    ) i__carry_i_8 (
        .I0(\simple_cpu_inst/alu_in1_reg_n_0_[0] ),
        .I1(\simple_cpu_inst/alu_in2(0) ),
        .I2(\simple_cpu_inst/alu_in1_reg_n_0_[1] ),
        .I3(\simple_cpu_inst/alu_in2(1) ),
        .O(i__carry_i_8_n_0)
    );

    LUT4 #(
        .INIT(16'h9009)
    ) i__carry__1_i_5 (
        .I0(\simple_cpu_inst/alu_in2(23) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[23] ),
        .I2(\simple_cpu_inst/alu_in2(22) ),
        .I3(\simple_cpu_inst/alu_in1_reg_n_0_[22] ),
        .O(i__carry__1_i_5_n_0)
    );

    LUT4 #(
        .INIT(16'h9009)
    ) i__carry__1_i_6 (
        .I0(\simple_cpu_inst/alu_in2(21) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[21] ),
        .I2(\simple_cpu_inst/alu_in2(20) ),
        .I3(\simple_cpu_inst/alu_in1_reg_n_0_[20] ),
        .O(i__carry__1_i_6_n_0)
    );

    LUT4 #(
        .INIT(16'h9009)
    ) i__carry_i_6 (
        .I0(\simple_cpu_inst/alu_in2(5) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[5] ),
        .I2(\simple_cpu_inst/alu_in1_reg_n_0_[4] ),
        .I3(\simple_cpu_inst/alu_in2(4) ),
        .O(i__carry_i_6_n_0)
    );

    LUT4 #(
        .INIT(16'h9009)
    ) i__carry__1_i_7 (
        .I0(\simple_cpu_inst/alu_in2(19) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[19] ),
        .I2(\simple_cpu_inst/alu_in2(18) ),
        .I3(\simple_cpu_inst/alu_in1_reg_n_0_[18] ),
        .O(i__carry__1_i_7_n_0)
    );

    LUT4 #(
        .INIT(16'h9009)
    ) i__carry_i_7 (
        .I0(\simple_cpu_inst/alu_in1_reg_n_0_[3] ),
        .I1(\simple_cpu_inst/alu_in2(3) ),
        .I2(\simple_cpu_inst/alu_in1_reg_n_0_[2] ),
        .I3(\simple_cpu_inst/alu_in2(2) ),
        .O(i__carry_i_7_n_0)
    );

    LUT4 #(
        .INIT(16'h22B2)
    ) i__carry_i_4 (
        .I0(\simple_cpu_inst/alu_in2(1) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[1] ),
        .I2(\simple_cpu_inst/alu_in2(0) ),
        .I3(\simple_cpu_inst/alu_in1_reg_n_0_[0] ),
        .O(i__carry_i_4_n_0)
    );

    LUT4 #(
        .INIT(16'h9009)
    ) i__carry_i_5 (
        .I0(\simple_cpu_inst/alu_in2(7) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[7] ),
        .I2(\simple_cpu_inst/alu_in2(6) ),
        .I3(\simple_cpu_inst/alu_in1_reg_n_0_[6] ),
        .O(i__carry_i_5_n_0)
    );

    LUT4 #(
        .INIT(16'h44D4)
    ) i__carry__1_i_3__1 (
        .I0(\simple_cpu_inst/alu_in1_reg_n_0_[19] ),
        .I1(\simple_cpu_inst/alu_in2(19) ),
        .I2(\simple_cpu_inst/alu_in2(18) ),
        .I3(\simple_cpu_inst/alu_in1_reg_n_0_[18] ),
        .O(i__carry__1_i_3__1_n_0)
    );

    LUT4 #(
        .INIT(16'h44D4)
    ) i__carry__0_i_3__1 (
        .I0(\simple_cpu_inst/alu_in1_reg_n_0_[11] ),
        .I1(\simple_cpu_inst/alu_in2(11) ),
        .I2(\simple_cpu_inst/alu_in2(10) ),
        .I3(\simple_cpu_inst/alu_in1_reg_n_0_[10] ),
        .O(i__carry__0_i_3__1_n_0)
    );

    LUT4 #(
        .INIT(16'h9009)
    ) i__carry__2_i_6 (
        .I0(\simple_cpu_inst/alu_in2(29) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[29] ),
        .I2(\simple_cpu_inst/alu_in2(28) ),
        .I3(\simple_cpu_inst/alu_in1_reg_n_0_[28] ),
        .O(i__carry__2_i_6_n_0)
    );

    LUT4 #(
        .INIT(16'h44D4)
    ) i__carry__1_i_2__1 (
        .I0(\simple_cpu_inst/alu_in1_reg_n_0_[21] ),
        .I1(\simple_cpu_inst/alu_in2(21) ),
        .I2(\simple_cpu_inst/alu_in2(20) ),
        .I3(\simple_cpu_inst/alu_in1_reg_n_0_[20] ),
        .O(i__carry__1_i_2__1_n_0)
    );

    LUT4 #(
        .INIT(16'h44D4)
    ) i__carry__0_i_2__1 (
        .I0(\simple_cpu_inst/alu_in1_reg_n_0_[13] ),
        .I1(\simple_cpu_inst/alu_in2(13) ),
        .I2(\simple_cpu_inst/alu_in2(12) ),
        .I3(\simple_cpu_inst/alu_in1_reg_n_0_[12] ),
        .O(i__carry__0_i_2__1_n_0)
    );

    CARRY4 \simple_cpu_inst/alu_inst/acc0_inferred__4/i__carry  (
        .CI(1'b0),
        .CYINIT(1'b0),
        .DI({
            i__carry_i_1__1_n_0,
            i__carry_i_2__1_n_0,
            i__carry_i_3__0_n_0,
            i__carry_i_4_n_0
        }),
        .S({
            i__carry_i_5_n_0,
            i__carry_i_6_n_0,
            i__carry_i_7_n_0,
            i__carry_i_8_n_0
        }),
        .CO({
            \simple_cpu_inst/alu_inst/acc0_inferred__4/i__carry_n_0 ,
            \simple_cpu_inst/alu_inst/acc0_inferred__4/i__carry_n_1 ,
            \simple_cpu_inst/alu_inst/acc0_inferred__4/i__carry_n_2 ,
            \simple_cpu_inst/alu_inst/acc0_inferred__4/i__carry_n_3 
        })
    );

    CARRY4 \simple_cpu_inst/alu_inst/acc0_inferred__4/i__carry__0  (
        .CI(\simple_cpu_inst/alu_inst/acc0_inferred__4/i__carry_n_0 ),
        .CYINIT(1'b0),
        .DI({
            i__carry__0_i_1__1_n_0,
            i__carry__0_i_2__1_n_0,
            i__carry__0_i_3__1_n_0,
            i__carry__0_i_4__1_n_0
        }),
        .S({
            i__carry__0_i_5_n_0,
            i__carry__0_i_6_n_0,
            i__carry__0_i_7_n_0,
            i__carry__0_i_8_n_0
        }),
        .CO({
            \simple_cpu_inst/alu_inst/acc0_inferred__4/i__carry__0_n_0 ,
            \simple_cpu_inst/alu_inst/acc0_inferred__4/i__carry__0_n_1 ,
            \simple_cpu_inst/alu_inst/acc0_inferred__4/i__carry__0_n_2 ,
            \simple_cpu_inst/alu_inst/acc0_inferred__4/i__carry__0_n_3 
        })
    );

    LUT4 #(
        .INIT(16'h44D4)
    ) i__carry__2_i_4__1 (
        .I0(\simple_cpu_inst/alu_in1_reg_n_0_[25] ),
        .I1(\simple_cpu_inst/alu_in2(25) ),
        .I2(\simple_cpu_inst/alu_in2(24) ),
        .I3(\simple_cpu_inst/alu_in1_reg_n_0_[24] ),
        .O(i__carry__2_i_4__1_n_0)
    );

    LUT4 #(
        .INIT(16'h44D4)
    ) i__carry__1_i_1__1 (
        .I0(\simple_cpu_inst/alu_in1_reg_n_0_[23] ),
        .I1(\simple_cpu_inst/alu_in2(23) ),
        .I2(\simple_cpu_inst/alu_in2(22) ),
        .I3(\simple_cpu_inst/alu_in1_reg_n_0_[22] ),
        .O(i__carry__1_i_1__1_n_0)
    );

    LUT4 #(
        .INIT(16'h44D4)
    ) i__carry__0_i_1__1 (
        .I0(\simple_cpu_inst/alu_in1_reg_n_0_[15] ),
        .I1(\simple_cpu_inst/alu_in2(15) ),
        .I2(\simple_cpu_inst/alu_in2(14) ),
        .I3(\simple_cpu_inst/alu_in1_reg_n_0_[14] ),
        .O(i__carry__0_i_1__1_n_0)
    );

    LUT4 #(
        .INIT(16'h9009)
    ) i__carry__2_i_5 (
        .I0(\simple_cpu_inst/alu_in2(31) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[31] ),
        .I2(\simple_cpu_inst/alu_in2(30) ),
        .I3(\simple_cpu_inst/alu_in1_reg_n_0_[30] ),
        .O(i__carry__2_i_5_n_0)
    );

    LUT4 #(
        .INIT(16'h9009)
    ) i__carry__0_i_8 (
        .I0(\simple_cpu_inst/alu_in2(9) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[9] ),
        .I2(\simple_cpu_inst/alu_in2(8) ),
        .I3(\simple_cpu_inst/alu_in1_reg_n_0_[8] ),
        .O(i__carry__0_i_8_n_0)
    );

    LUT4 #(
        .INIT(16'h22B2)
    ) i__carry_i_3__0 (
        .I0(\simple_cpu_inst/alu_in2(3) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[3] ),
        .I2(\simple_cpu_inst/alu_in2(2) ),
        .I3(\simple_cpu_inst/alu_in1_reg_n_0_[2] ),
        .O(i__carry_i_3__0_n_0)
    );

    LUT4 #(
        .INIT(16'h9009)
    ) i__carry__0_i_6 (
        .I0(\simple_cpu_inst/alu_in2(13) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[13] ),
        .I2(\simple_cpu_inst/alu_in2(12) ),
        .I3(\simple_cpu_inst/alu_in1_reg_n_0_[12] ),
        .O(i__carry__0_i_6_n_0)
    );

    LUT4 #(
        .INIT(16'h9009)
    ) i__carry__0_i_7 (
        .I0(\simple_cpu_inst/alu_in2(11) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[11] ),
        .I2(\simple_cpu_inst/alu_in2(10) ),
        .I3(\simple_cpu_inst/alu_in1_reg_n_0_[10] ),
        .O(i__carry__0_i_7_n_0)
    );

    LUT4 #(
        .INIT(16'h44D4)
    ) i__carry_i_2__1 (
        .I0(\simple_cpu_inst/alu_in1_reg_n_0_[5] ),
        .I1(\simple_cpu_inst/alu_in2(5) ),
        .I2(\simple_cpu_inst/alu_in2(4) ),
        .I3(\simple_cpu_inst/alu_in1_reg_n_0_[4] ),
        .O(i__carry_i_2__1_n_0)
    );

    LUT4 #(
        .INIT(16'h44D4)
    ) i__carry__2_i_3__1 (
        .I0(\simple_cpu_inst/alu_in1_reg_n_0_[27] ),
        .I1(\simple_cpu_inst/alu_in2(27) ),
        .I2(\simple_cpu_inst/alu_in2(26) ),
        .I3(\simple_cpu_inst/alu_in1_reg_n_0_[26] ),
        .O(i__carry__2_i_3__1_n_0)
    );

    LUT4 #(
        .INIT(16'h44D4)
    ) i__carry__0_i_4__1 (
        .I0(\simple_cpu_inst/alu_in1_reg_n_0_[9] ),
        .I1(\simple_cpu_inst/alu_in2(9) ),
        .I2(\simple_cpu_inst/alu_in2(8) ),
        .I3(\simple_cpu_inst/alu_in1_reg_n_0_[8] ),
        .O(i__carry__0_i_4__1_n_0)
    );

    LUT4 #(
        .INIT(16'h44D4)
    ) i__carry__2_i_2__1 (
        .I0(\simple_cpu_inst/alu_in1_reg_n_0_[29] ),
        .I1(\simple_cpu_inst/alu_in2(29) ),
        .I2(\simple_cpu_inst/alu_in2(28) ),
        .I3(\simple_cpu_inst/alu_in1_reg_n_0_[28] ),
        .O(i__carry__2_i_2__1_n_0)
    );

    LUT4 #(
        .INIT(16'h44D4)
    ) i__carry_i_1__1 (
        .I0(\simple_cpu_inst/alu_in1_reg_n_0_[7] ),
        .I1(\simple_cpu_inst/alu_in2(7) ),
        .I2(\simple_cpu_inst/alu_in2(6) ),
        .I3(\simple_cpu_inst/alu_in1_reg_n_0_[6] ),
        .O(i__carry_i_1__1_n_0)
    );

    LUT4 #(
        .INIT(16'h9009)
    ) i__carry__0_i_5 (
        .I0(\simple_cpu_inst/alu_in2(15) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[15] ),
        .I2(\simple_cpu_inst/alu_in2(14) ),
        .I3(\simple_cpu_inst/alu_in1_reg_n_0_[14] ),
        .O(i__carry__0_i_5_n_0)
    );

    LUT4 #(
        .INIT(16'h2F02)
    ) i__carry__2_i_1__2 (
        .I0(\simple_cpu_inst/alu_in2(30) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[30] ),
        .I2(\simple_cpu_inst/alu_in1_reg_n_0_[31] ),
        .I3(\simple_cpu_inst/alu_in2(31) ),
        .O(i__carry__2_i_1__2_n_0)
    );

    LUT4 #(
        .INIT(16'h9009)
    ) i__carry__2_i_7 (
        .I0(\simple_cpu_inst/alu_in2(27) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[27] ),
        .I2(\simple_cpu_inst/alu_in2(26) ),
        .I3(\simple_cpu_inst/alu_in1_reg_n_0_[26] ),
        .O(i__carry__2_i_7_n_0)
    );
endmodule

