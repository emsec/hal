`timescale 1 ps/1 ps
module top(\simple_cpu_inst/alu_in2(21) ,\simple_cpu_inst/alu_in1_reg_n_0_[0] ,\simple_cpu_inst/alu_in1_reg_n_0_[3] ,\simple_cpu_inst/alu_in2(2) ,\simple_cpu_inst/alu_in1_reg_n_0_[2] ,\simple_cpu_inst/alu_in1_reg_n_0_[5] ,\simple_cpu_inst/alu_in1_reg_n_0_[25] ,\simple_cpu_inst/alu_in2(16) ,\simple_cpu_inst/alu_in1_reg_n_0_[30] ,\simple_cpu_inst/alu_in1_reg_n_0_[7] ,\simple_cpu_inst/alu_in2(22) ,\simple_cpu_inst/alu_in2(3) ,\simple_cpu_inst/alu_in2(7) ,\simple_cpu_inst/alu_in1_reg_n_0_[9] ,\simple_cpu_inst/alu_in1_reg_n_0_[14] ,\simple_cpu_inst/alu_in1_reg_n_0_[4] ,\simple_cpu_inst/alu_in2(28) ,\simple_cpu_inst/alu_in2(8) ,\simple_cpu_inst/alu_in2(30) ,\simple_cpu_inst/alu_in2(11) ,\simple_cpu_inst/alu_in2(25) ,\simple_cpu_inst/alu_in1_reg_n_0_[23] ,\simple_cpu_inst/alu_in1_reg_n_0_[26] ,\simple_cpu_inst/alu_in2(19) ,\simple_cpu_inst/alu_in2(29) ,\simple_cpu_inst/alu_in1_reg_n_0_[18] ,\simple_cpu_inst/alu_in2(4) ,\simple_cpu_inst/alu_in1_reg_n_0_[22] ,\simple_cpu_inst/alu_in2(27) ,\simple_cpu_inst/alu_in2(5) ,\simple_cpu_inst/alu_in1_reg_n_0_[16] ,\simple_cpu_inst/alu_in1_reg_n_0_[19] ,\simple_cpu_inst/alu_in1_reg_n_0_[6] ,\simple_cpu_inst/alu_in1_reg_n_0_[21] ,\simple_cpu_inst/alu_in2(24) ,\simple_cpu_inst/alu_in1_reg_n_0_[10] ,\simple_cpu_inst/alu_in2(9) ,\simple_cpu_inst/alu_in2(6) ,\simple_cpu_inst/alu_in2(10) ,\simple_cpu_inst/alu_in2(26) ,\simple_cpu_inst/alu_in2(17) ,\simple_cpu_inst/alu_in1_reg_n_0_[28] ,\simple_cpu_inst/alu_in1_reg_n_0_[11] ,\simple_cpu_inst/alu_in1_reg_n_0_[1] ,\simple_cpu_inst/alu_in1_reg_n_0_[20] ,\simple_cpu_inst/alu_in2(23) ,\simple_cpu_inst/alu_in1_reg_n_0_[15] ,\simple_cpu_inst/alu_in2(31) ,\simple_cpu_inst/alu_in2(14) ,\simple_cpu_inst/alu_in2(12) ,\simple_cpu_inst/alu_in2(0) ,\simple_cpu_inst/alu_in1_reg_n_0_[29] ,\simple_cpu_inst/alu_in2(18) ,\simple_cpu_inst/alu_in1_reg_n_0_[8] ,\simple_cpu_inst/alu_in2(20) ,\simple_cpu_inst/alu_in1_reg_n_0_[31] ,\simple_cpu_inst/alu_in2(13) ,\simple_cpu_inst/alu_in1_reg_n_0_[24] ,\simple_cpu_inst/alu_in2(15) ,\simple_cpu_inst/alu_in1_reg_n_0_[13] ,\simple_cpu_inst/alu_in1_reg_n_0_[12] ,\simple_cpu_inst/alu_in1_reg_n_0_[27] ,\simple_cpu_inst/alu_in2(1) ,\simple_cpu_inst/alu_in1_reg_n_0_[17] ,\simple_cpu_inst/alu_inst/data2(5) ,\simple_cpu_inst/alu_inst/data2(16) ,\simple_cpu_inst/alu_inst/data2(12) ,\simple_cpu_inst/alu_inst/data2(17) ,\simple_cpu_inst/alu_inst/data2(13) ,\simple_cpu_inst/alu_inst/data2(15) ,\simple_cpu_inst/alu_inst/data2(31) ,\simple_cpu_inst/alu_inst/data2(25) ,\simple_cpu_inst/alu_inst/data2(24) ,\simple_cpu_inst/alu_inst/data2(19) ,\simple_cpu_inst/alu_inst/data2(29) ,\simple_cpu_inst/alu_inst/data2(7) ,\simple_cpu_inst/alu_inst/data2(6) ,\simple_cpu_inst/alu_inst/data2(2) ,\simple_cpu_inst/alu_inst/data2(18) ,\simple_cpu_inst/alu_inst/data2(23) ,\simple_cpu_inst/alu_inst/data2(1) ,\simple_cpu_inst/alu_inst/data2(11) ,\simple_cpu_inst/alu_inst/data2(9) ,\NLW_write_addr_reg[3]_i_8_O_UNCONNECTED(0) ,\simple_cpu_inst/alu_inst/data2(10) ,\simple_cpu_inst/alu_inst/data2(30) ,\simple_cpu_inst/alu_inst/data2(4) ,\simple_cpu_inst/alu_inst/data2(22) ,\simple_cpu_inst/alu_inst/data2(8) ,\simple_cpu_inst/alu_inst/data2(21) ,\simple_cpu_inst/alu_inst/data2(14) ,\simple_cpu_inst/alu_inst/data2(28) ,\simple_cpu_inst/alu_inst/data2(27) ,\simple_cpu_inst/alu_inst/data2(20) ,\simple_cpu_inst/alu_inst/data2(3) ,\simple_cpu_inst/alu_inst/data2(26) );
    input \simple_cpu_inst/alu_in2(21) ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[0] ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[3] ;
    input \simple_cpu_inst/alu_in2(2) ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[2] ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[5] ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[25] ;
    input \simple_cpu_inst/alu_in2(16) ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[30] ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[7] ;
    input \simple_cpu_inst/alu_in2(22) ;
    input \simple_cpu_inst/alu_in2(3) ;
    input \simple_cpu_inst/alu_in2(7) ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[9] ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[14] ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[4] ;
    input \simple_cpu_inst/alu_in2(28) ;
    input \simple_cpu_inst/alu_in2(8) ;
    input \simple_cpu_inst/alu_in2(30) ;
    input \simple_cpu_inst/alu_in2(11) ;
    input \simple_cpu_inst/alu_in2(25) ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[23] ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[26] ;
    input \simple_cpu_inst/alu_in2(19) ;
    input \simple_cpu_inst/alu_in2(29) ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[18] ;
    input \simple_cpu_inst/alu_in2(4) ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[22] ;
    input \simple_cpu_inst/alu_in2(27) ;
    input \simple_cpu_inst/alu_in2(5) ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[16] ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[19] ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[6] ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[21] ;
    input \simple_cpu_inst/alu_in2(24) ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[10] ;
    input \simple_cpu_inst/alu_in2(9) ;
    input \simple_cpu_inst/alu_in2(6) ;
    input \simple_cpu_inst/alu_in2(10) ;
    input \simple_cpu_inst/alu_in2(26) ;
    input \simple_cpu_inst/alu_in2(17) ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[28] ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[11] ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[1] ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[20] ;
    input \simple_cpu_inst/alu_in2(23) ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[15] ;
    input \simple_cpu_inst/alu_in2(31) ;
    input \simple_cpu_inst/alu_in2(14) ;
    input \simple_cpu_inst/alu_in2(12) ;
    input \simple_cpu_inst/alu_in2(0) ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[29] ;
    input \simple_cpu_inst/alu_in2(18) ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[8] ;
    input \simple_cpu_inst/alu_in2(20) ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[31] ;
    input \simple_cpu_inst/alu_in2(13) ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[24] ;
    input \simple_cpu_inst/alu_in2(15) ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[13] ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[12] ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[27] ;
    input \simple_cpu_inst/alu_in2(1) ;
    input \simple_cpu_inst/alu_in1_reg_n_0_[17] ;
    output \simple_cpu_inst/alu_inst/data2(5) ;
    output \simple_cpu_inst/alu_inst/data2(16) ;
    output \simple_cpu_inst/alu_inst/data2(12) ;
    output \simple_cpu_inst/alu_inst/data2(17) ;
    output \simple_cpu_inst/alu_inst/data2(13) ;
    output \simple_cpu_inst/alu_inst/data2(15) ;
    output \simple_cpu_inst/alu_inst/data2(31) ;
    output \simple_cpu_inst/alu_inst/data2(25) ;
    output \simple_cpu_inst/alu_inst/data2(24) ;
    output \simple_cpu_inst/alu_inst/data2(19) ;
    output \simple_cpu_inst/alu_inst/data2(29) ;
    output \simple_cpu_inst/alu_inst/data2(7) ;
    output \simple_cpu_inst/alu_inst/data2(6) ;
    output \simple_cpu_inst/alu_inst/data2(2) ;
    output \simple_cpu_inst/alu_inst/data2(18) ;
    output \simple_cpu_inst/alu_inst/data2(23) ;
    output \simple_cpu_inst/alu_inst/data2(1) ;
    output \simple_cpu_inst/alu_inst/data2(11) ;
    output \simple_cpu_inst/alu_inst/data2(9) ;
    output \NLW_write_addr_reg[3]_i_8_O_UNCONNECTED(0) ;
    output \simple_cpu_inst/alu_inst/data2(10) ;
    output \simple_cpu_inst/alu_inst/data2(30) ;
    output \simple_cpu_inst/alu_inst/data2(4) ;
    output \simple_cpu_inst/alu_inst/data2(22) ;
    output \simple_cpu_inst/alu_inst/data2(8) ;
    output \simple_cpu_inst/alu_inst/data2(21) ;
    output \simple_cpu_inst/alu_inst/data2(14) ;
    output \simple_cpu_inst/alu_inst/data2(28) ;
    output \simple_cpu_inst/alu_inst/data2(27) ;
    output \simple_cpu_inst/alu_inst/data2(20) ;
    output \simple_cpu_inst/alu_inst/data2(3) ;
    output \simple_cpu_inst/alu_inst/data2(26) ;
    wire \write_addr[7]_i_13_n_0 ;
    wire \write_addr[7]_i_14_n_0 ;
    wire \write_addr[7]_i_15_n_0 ;
    wire \write_addr_reg[3]_i_8_n_0 ;
    wire \write_addr_reg[15]_i_5_n_1 ;
    wire \write_addr_reg[7]_i_8_n_1 ;
    wire \write_addr[11]_i_12_n_0 ;
    wire \write_addr_reg[3]_i_8_n_1 ;
    wire \write_addr_reg[23]_i_9_n_3 ;
    wire \write_addr_reg[7]_i_8_n_3 ;
    wire \write_addr_reg[7]_i_8_n_0 ;
    wire \write_addr_reg[7]_i_8_n_2 ;
    wire \write_addr[15]_i_10_n_0 ;
    wire \write_addr_reg[15]_i_5_n_0 ;
    wire \write_addr_reg[31]_i_8_n_3 ;
    wire \write_addr_reg[15]_i_5_n_2 ;
    wire \write_addr[3]_i_15_n_0 ;
    wire \write_addr[15]_i_11_n_0 ;
    wire \write_addr[27]_i_16_n_0 ;
    wire \write_addr[19]_i_27_n_0 ;
    wire \write_addr[3]_i_18_n_0 ;
    wire \write_addr_reg[15]_i_5_n_3 ;
    wire \write_addr_reg[31]_i_8_n_2 ;
    wire \write_addr_reg[11]_i_5_n_0 ;
    wire \write_addr[15]_i_12_n_0 ;
    wire \write_addr[27]_i_15_n_0 ;
    wire \write_addr[3]_i_16_n_0 ;
    wire \write_addr[15]_i_13_n_0 ;
    wire \write_addr[27]_i_13_n_0 ;
    wire \write_addr[23]_i_16_n_0 ;
    wire \write_addr[19]_i_29_n_0 ;
    wire \write_addr[19]_i_26_n_0 ;
    wire \write_addr[7]_i_12_n_0 ;
    wire \write_addr[31]_i_15_n_0 ;
    wire \write_addr[31]_i_16_n_0 ;
    wire \write_addr_reg[19]_i_13_n_3 ;
    wire \write_addr[27]_i_14_n_0 ;
    wire \write_addr_reg[23]_i_9_n_1 ;
    wire \write_addr_reg[27]_i_6_n_2 ;
    wire \write_addr_reg[19]_i_13_n_2 ;
    wire \write_addr_reg[19]_i_13_n_1 ;
    wire \write_addr[23]_i_19_n_0 ;
    wire \write_addr[23]_i_18_n_0 ;
    wire \write_addr[11]_i_11_n_0 ;
    wire \write_addr[31]_i_13_n_0 ;
    wire \write_addr[3]_i_17_n_0 ;
    wire \write_addr[23]_i_17_n_0 ;
    wire \write_addr_reg[23]_i_9_n_2 ;
    wire \write_addr_reg[3]_i_8_n_3 ;
    wire \write_addr_reg[23]_i_9_n_0 ;
    wire \write_addr[31]_i_14_n_0 ;
    wire \write_addr_reg[11]_i_5_n_2 ;
    wire \write_addr_reg[3]_i_8_n_2 ;
    wire \write_addr_reg[27]_i_6_n_1 ;
    wire \write_addr[11]_i_13_n_0 ;
    wire \write_addr_reg[31]_i_8_n_1 ;
    wire \write_addr_reg[27]_i_6_n_0 ;
    wire \write_addr_reg[19]_i_13_n_0 ;
    wire \write_addr[11]_i_10_n_0 ;
    wire \write_addr[19]_i_28_n_0 ;
    wire \write_addr_reg[27]_i_6_n_3 ;
    wire \write_addr_reg[11]_i_5_n_1 ;
    wire \write_addr_reg[11]_i_5_n_3 ;

    CARRY4 \write_addr_reg[7]_i_8  (
        .CI(\write_addr_reg[3]_i_8_n_0 ),
        .CYINIT(1'b0 ),
        .DI({
            \simple_cpu_inst/alu_in1_reg_n_0_[7] ,
            \simple_cpu_inst/alu_in1_reg_n_0_[6] ,
            \simple_cpu_inst/alu_in1_reg_n_0_[5] ,
            \simple_cpu_inst/alu_in1_reg_n_0_[4] 
        }),
        .S({
            \write_addr[7]_i_12_n_0 ,
            \write_addr[7]_i_13_n_0 ,
            \write_addr[7]_i_14_n_0 ,
            \write_addr[7]_i_15_n_0 
        }),
        .CO({
            \write_addr_reg[7]_i_8_n_0 ,
            \write_addr_reg[7]_i_8_n_1 ,
            \write_addr_reg[7]_i_8_n_2 ,
            \write_addr_reg[7]_i_8_n_3 
        }),
        .O({
            \simple_cpu_inst/alu_inst/data2(7) ,
            \simple_cpu_inst/alu_inst/data2(6) ,
            \simple_cpu_inst/alu_inst/data2(5) ,
            \simple_cpu_inst/alu_inst/data2(4) 
        })
    );

    LUT2 #(
        .INIT(4'h9)
    ) \write_addr[3]_i_16  (
        .I0(\simple_cpu_inst/alu_in1_reg_n_0_[2] ),
        .I1(\simple_cpu_inst/alu_in2(2) ),
        .O(\write_addr[3]_i_16_n_0 )
    );

    LUT2 #(
        .INIT(4'h9)
    ) \write_addr[7]_i_12  (
        .I0(\simple_cpu_inst/alu_in2(7) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[7] ),
        .O(\write_addr[7]_i_12_n_0 )
    );

    LUT2 #(
        .INIT(4'h9)
    ) \write_addr[3]_i_15  (
        .I0(\simple_cpu_inst/alu_in1_reg_n_0_[3] ),
        .I1(\simple_cpu_inst/alu_in2(3) ),
        .O(\write_addr[3]_i_15_n_0 )
    );

    CARRY4 \write_addr_reg[15]_i_5  (
        .CI(\write_addr_reg[11]_i_5_n_0 ),
        .CYINIT(1'b0 ),
        .DI({
            \simple_cpu_inst/alu_in1_reg_n_0_[15] ,
            \simple_cpu_inst/alu_in1_reg_n_0_[14] ,
            \simple_cpu_inst/alu_in1_reg_n_0_[13] ,
            \simple_cpu_inst/alu_in1_reg_n_0_[12] 
        }),
        .S({
            \write_addr[15]_i_10_n_0 ,
            \write_addr[15]_i_11_n_0 ,
            \write_addr[15]_i_12_n_0 ,
            \write_addr[15]_i_13_n_0 
        }),
        .CO({
            \write_addr_reg[15]_i_5_n_0 ,
            \write_addr_reg[15]_i_5_n_1 ,
            \write_addr_reg[15]_i_5_n_2 ,
            \write_addr_reg[15]_i_5_n_3 
        }),
        .O({
            \simple_cpu_inst/alu_inst/data2(15) ,
            \simple_cpu_inst/alu_inst/data2(14) ,
            \simple_cpu_inst/alu_inst/data2(13) ,
            \simple_cpu_inst/alu_inst/data2(12) 
        })
    );

    LUT2 #(
        .INIT(4'h9)
    ) \write_addr[27]_i_15  (
        .I0(\simple_cpu_inst/alu_in2(25) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[25] ),
        .O(\write_addr[27]_i_15_n_0 )
    );

    LUT2 #(
        .INIT(4'h9)
    ) \write_addr[27]_i_14  (
        .I0(\simple_cpu_inst/alu_in2(26) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[26] ),
        .O(\write_addr[27]_i_14_n_0 )
    );

    LUT2 #(
        .INIT(4'h9)
    ) \write_addr[7]_i_15  (
        .I0(\simple_cpu_inst/alu_in1_reg_n_0_[4] ),
        .I1(\simple_cpu_inst/alu_in2(4) ),
        .O(\write_addr[7]_i_15_n_0 )
    );

    LUT2 #(
        .INIT(4'h9)
    ) \write_addr[27]_i_13  (
        .I0(\simple_cpu_inst/alu_in2(27) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[27] ),
        .O(\write_addr[27]_i_13_n_0 )
    );

    LUT2 #(
        .INIT(4'h9)
    ) \write_addr[7]_i_14  (
        .I0(\simple_cpu_inst/alu_in2(5) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[5] ),
        .O(\write_addr[7]_i_14_n_0 )
    );

    LUT2 #(
        .INIT(4'h9)
    ) \write_addr[7]_i_13  (
        .I0(\simple_cpu_inst/alu_in2(6) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[6] ),
        .O(\write_addr[7]_i_13_n_0 )
    );

    CARRY4 \write_addr_reg[19]_i_13  (
        .CI(\write_addr_reg[15]_i_5_n_0 ),
        .CYINIT(1'b0 ),
        .DI({
            \simple_cpu_inst/alu_in1_reg_n_0_[19] ,
            \simple_cpu_inst/alu_in1_reg_n_0_[18] ,
            \simple_cpu_inst/alu_in1_reg_n_0_[17] ,
            \simple_cpu_inst/alu_in1_reg_n_0_[16] 
        }),
        .S({
            \write_addr[19]_i_26_n_0 ,
            \write_addr[19]_i_27_n_0 ,
            \write_addr[19]_i_28_n_0 ,
            \write_addr[19]_i_29_n_0 
        }),
        .CO({
            \write_addr_reg[19]_i_13_n_0 ,
            \write_addr_reg[19]_i_13_n_1 ,
            \write_addr_reg[19]_i_13_n_2 ,
            \write_addr_reg[19]_i_13_n_3 
        }),
        .O({
            \simple_cpu_inst/alu_inst/data2(19) ,
            \simple_cpu_inst/alu_inst/data2(18) ,
            \simple_cpu_inst/alu_inst/data2(17) ,
            \simple_cpu_inst/alu_inst/data2(16) 
        })
    );

    LUT2 #(
        .INIT(4'h9)
    ) \write_addr[15]_i_13  (
        .I0(\simple_cpu_inst/alu_in2(12) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[12] ),
        .O(\write_addr[15]_i_13_n_0 )
    );

    LUT2 #(
        .INIT(4'h9)
    ) \write_addr[15]_i_12  (
        .I0(\simple_cpu_inst/alu_in2(13) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[13] ),
        .O(\write_addr[15]_i_12_n_0 )
    );

    LUT2 #(
        .INIT(4'h9)
    ) \write_addr[11]_i_11  (
        .I0(\simple_cpu_inst/alu_in2(10) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[10] ),
        .O(\write_addr[11]_i_11_n_0 )
    );

    LUT2 #(
        .INIT(4'h9)
    ) \write_addr[11]_i_10  (
        .I0(\simple_cpu_inst/alu_in2(11) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[11] ),
        .O(\write_addr[11]_i_10_n_0 )
    );

    LUT2 #(
        .INIT(4'h9)
    ) \write_addr[19]_i_28  (
        .I0(\simple_cpu_inst/alu_in2(17) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[17] ),
        .O(\write_addr[19]_i_28_n_0 )
    );

    LUT2 #(
        .INIT(4'h9)
    ) \write_addr[23]_i_19  (
        .I0(\simple_cpu_inst/alu_in2(20) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[20] ),
        .O(\write_addr[23]_i_19_n_0 )
    );

    LUT2 #(
        .INIT(4'h9)
    ) \write_addr[19]_i_27  (
        .I0(\simple_cpu_inst/alu_in2(18) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[18] ),
        .O(\write_addr[19]_i_27_n_0 )
    );

    LUT2 #(
        .INIT(4'h9)
    ) \write_addr[23]_i_18  (
        .I0(\simple_cpu_inst/alu_in2(21) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[21] ),
        .O(\write_addr[23]_i_18_n_0 )
    );

    LUT2 #(
        .INIT(4'h9)
    ) \write_addr[19]_i_26  (
        .I0(\simple_cpu_inst/alu_in2(19) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[19] ),
        .O(\write_addr[19]_i_26_n_0 )
    );

    LUT2 #(
        .INIT(4'h9)
    ) \write_addr[23]_i_17  (
        .I0(\simple_cpu_inst/alu_in2(22) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[22] ),
        .O(\write_addr[23]_i_17_n_0 )
    );

    LUT2 #(
        .INIT(4'h9)
    ) \write_addr[15]_i_11  (
        .I0(\simple_cpu_inst/alu_in2(14) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[14] ),
        .O(\write_addr[15]_i_11_n_0 )
    );

    LUT2 #(
        .INIT(4'h9)
    ) \write_addr[3]_i_18  (
        .I0(\simple_cpu_inst/alu_in1_reg_n_0_[0] ),
        .I1(\simple_cpu_inst/alu_in2(0) ),
        .O(\write_addr[3]_i_18_n_0 )
    );

    LUT2 #(
        .INIT(4'h9)
    ) \write_addr[31]_i_16  (
        .I0(\simple_cpu_inst/alu_in2(28) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[28] ),
        .O(\write_addr[31]_i_16_n_0 )
    );

    CARRY4 \write_addr_reg[3]_i_8  (
        .CI(1'b0 ),
        .CYINIT(1'b1 ),
        .DI({
            \simple_cpu_inst/alu_in1_reg_n_0_[3] ,
            \simple_cpu_inst/alu_in1_reg_n_0_[2] ,
            \simple_cpu_inst/alu_in1_reg_n_0_[1] ,
            \simple_cpu_inst/alu_in1_reg_n_0_[0] 
        }),
        .S({
            \write_addr[3]_i_15_n_0 ,
            \write_addr[3]_i_16_n_0 ,
            \write_addr[3]_i_17_n_0 ,
            \write_addr[3]_i_18_n_0 
        }),
        .CO({
            \write_addr_reg[3]_i_8_n_0 ,
            \write_addr_reg[3]_i_8_n_1 ,
            \write_addr_reg[3]_i_8_n_2 ,
            \write_addr_reg[3]_i_8_n_3 
        }),
        .O({
            \simple_cpu_inst/alu_inst/data2(3) ,
            \simple_cpu_inst/alu_inst/data2(2) ,
            \simple_cpu_inst/alu_inst/data2(1) ,
            \NLW_write_addr_reg[3]_i_8_O_UNCONNECTED(0) 
        })
    );

    LUT2 #(
        .INIT(4'h9)
    ) \write_addr[23]_i_16  (
        .I0(\simple_cpu_inst/alu_in2(23) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[23] ),
        .O(\write_addr[23]_i_16_n_0 )
    );

    LUT2 #(
        .INIT(4'h9)
    ) \write_addr[15]_i_10  (
        .I0(\simple_cpu_inst/alu_in2(15) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[15] ),
        .O(\write_addr[15]_i_10_n_0 )
    );

    LUT2 #(
        .INIT(4'h9)
    ) \write_addr[3]_i_17  (
        .I0(\simple_cpu_inst/alu_in1_reg_n_0_[1] ),
        .I1(\simple_cpu_inst/alu_in2(1) ),
        .O(\write_addr[3]_i_17_n_0 )
    );

    LUT2 #(
        .INIT(4'h9)
    ) \write_addr[31]_i_15  (
        .I0(\simple_cpu_inst/alu_in2(29) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[29] ),
        .O(\write_addr[31]_i_15_n_0 )
    );

    LUT2 #(
        .INIT(4'h9)
    ) \write_addr[31]_i_14  (
        .I0(\simple_cpu_inst/alu_in2(30) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[30] ),
        .O(\write_addr[31]_i_14_n_0 )
    );

    CARRY4 \write_addr_reg[31]_i_8  (
        .CI(\write_addr_reg[27]_i_6_n_0 ),
        .CYINIT(1'b0 ),
        .DI({
            1'b0 ,
            \simple_cpu_inst/alu_in1_reg_n_0_[30] ,
            \simple_cpu_inst/alu_in1_reg_n_0_[29] ,
            \simple_cpu_inst/alu_in1_reg_n_0_[28] 
        }),
        .S({
            \write_addr[31]_i_13_n_0 ,
            \write_addr[31]_i_14_n_0 ,
            \write_addr[31]_i_15_n_0 ,
            \write_addr[31]_i_16_n_0 
        }),
        .CO({
            1'bz,
            \write_addr_reg[31]_i_8_n_1 ,
            \write_addr_reg[31]_i_8_n_2 ,
            \write_addr_reg[31]_i_8_n_3 
        }),
        .O({
            \simple_cpu_inst/alu_inst/data2(31) ,
            \simple_cpu_inst/alu_inst/data2(30) ,
            \simple_cpu_inst/alu_inst/data2(29) ,
            \simple_cpu_inst/alu_inst/data2(28) 
        })
    );

    LUT2 #(
        .INIT(4'h9)
    ) \write_addr[31]_i_13  (
        .I0(\simple_cpu_inst/alu_in2(31) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[31] ),
        .O(\write_addr[31]_i_13_n_0 )
    );

    LUT2 #(
        .INIT(4'h9)
    ) \write_addr[19]_i_29  (
        .I0(\simple_cpu_inst/alu_in2(16) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[16] ),
        .O(\write_addr[19]_i_29_n_0 )
    );

    LUT2 #(
        .INIT(4'h9)
    ) \write_addr[27]_i_16  (
        .I0(\simple_cpu_inst/alu_in2(24) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[24] ),
        .O(\write_addr[27]_i_16_n_0 )
    );

    CARRY4 \write_addr_reg[27]_i_6  (
        .CI(\write_addr_reg[23]_i_9_n_0 ),
        .CYINIT(1'b0 ),
        .DI({
            \simple_cpu_inst/alu_in1_reg_n_0_[27] ,
            \simple_cpu_inst/alu_in1_reg_n_0_[26] ,
            \simple_cpu_inst/alu_in1_reg_n_0_[25] ,
            \simple_cpu_inst/alu_in1_reg_n_0_[24] 
        }),
        .S({
            \write_addr[27]_i_13_n_0 ,
            \write_addr[27]_i_14_n_0 ,
            \write_addr[27]_i_15_n_0 ,
            \write_addr[27]_i_16_n_0 
        }),
        .CO({
            \write_addr_reg[27]_i_6_n_0 ,
            \write_addr_reg[27]_i_6_n_1 ,
            \write_addr_reg[27]_i_6_n_2 ,
            \write_addr_reg[27]_i_6_n_3 
        }),
        .O({
            \simple_cpu_inst/alu_inst/data2(27) ,
            \simple_cpu_inst/alu_inst/data2(26) ,
            \simple_cpu_inst/alu_inst/data2(25) ,
            \simple_cpu_inst/alu_inst/data2(24) 
        })
    );

    CARRY4 \write_addr_reg[23]_i_9  (
        .CI(\write_addr_reg[19]_i_13_n_0 ),
        .CYINIT(1'b0 ),
        .DI({
            \simple_cpu_inst/alu_in1_reg_n_0_[23] ,
            \simple_cpu_inst/alu_in1_reg_n_0_[22] ,
            \simple_cpu_inst/alu_in1_reg_n_0_[21] ,
            \simple_cpu_inst/alu_in1_reg_n_0_[20] 
        }),
        .S({
            \write_addr[23]_i_16_n_0 ,
            \write_addr[23]_i_17_n_0 ,
            \write_addr[23]_i_18_n_0 ,
            \write_addr[23]_i_19_n_0 
        }),
        .CO({
            \write_addr_reg[23]_i_9_n_0 ,
            \write_addr_reg[23]_i_9_n_1 ,
            \write_addr_reg[23]_i_9_n_2 ,
            \write_addr_reg[23]_i_9_n_3 
        }),
        .O({
            \simple_cpu_inst/alu_inst/data2(23) ,
            \simple_cpu_inst/alu_inst/data2(22) ,
            \simple_cpu_inst/alu_inst/data2(21) ,
            \simple_cpu_inst/alu_inst/data2(20) 
        })
    );

    LUT2 #(
        .INIT(4'h9)
    ) \write_addr[11]_i_13  (
        .I0(\simple_cpu_inst/alu_in2(8) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[8] ),
        .O(\write_addr[11]_i_13_n_0 )
    );

    LUT2 #(
        .INIT(4'h9)
    ) \write_addr[11]_i_12  (
        .I0(\simple_cpu_inst/alu_in2(9) ),
        .I1(\simple_cpu_inst/alu_in1_reg_n_0_[9] ),
        .O(\write_addr[11]_i_12_n_0 )
    );

    CARRY4 \write_addr_reg[11]_i_5  (
        .CI(\write_addr_reg[7]_i_8_n_0 ),
        .CYINIT(1'b0 ),
        .DI({
            \simple_cpu_inst/alu_in1_reg_n_0_[11] ,
            \simple_cpu_inst/alu_in1_reg_n_0_[10] ,
            \simple_cpu_inst/alu_in1_reg_n_0_[9] ,
            \simple_cpu_inst/alu_in1_reg_n_0_[8] 
        }),
        .S({
            \write_addr[11]_i_10_n_0 ,
            \write_addr[11]_i_11_n_0 ,
            \write_addr[11]_i_12_n_0 ,
            \write_addr[11]_i_13_n_0 
        }),
        .CO({
            \write_addr_reg[11]_i_5_n_0 ,
            \write_addr_reg[11]_i_5_n_1 ,
            \write_addr_reg[11]_i_5_n_2 ,
            \write_addr_reg[11]_i_5_n_3 
        }),
        .O({
            \simple_cpu_inst/alu_inst/data2(11) ,
            \simple_cpu_inst/alu_inst/data2(10) ,
            \simple_cpu_inst/alu_inst/data2(9) ,
            \simple_cpu_inst/alu_inst/data2(8) 
        })
    );
endmodule

