//-----------------------------------------------// 
//----	SB_MAC16 DSP Primitive             ------//
//-----------------------------------------------// 
`timescale 1ps/1ps
module SB_MAC16 (
		A,
		B,
		C,
		D,
		O,
		CLK,
		CE,
		IRSTTOP,
	    IRSTBOT,
		ORSTTOP,
		ORSTBOT,
		AHOLD,
		BHOLD,
		CHOLD,
		DHOLD,
		OHOLDTOP,
		OHOLDBOT,
		OLOADTOP,
		OLOADBOT,
		ADDSUBTOP,
		ADDSUBBOT,
		CO,
		CI,  		//from bottom tile
		ACCUMCI, 	// Carry input from MAC CO below
		ACCUMCO, 	// Carry output to above MAC block.    
		SIGNEXTIN,
		SIGNEXTOUT
);
output 	[31:0] O;	 // Output [31:0]
input	[15:0] A;        // data  to upper mult block / upper accum block.
input	[15:0] B;        // data  to lower mult block / lower accum block.   
input	[15:0] C;        // direct data  to upper accum block. 
input	[15:0] D;        // direct data  to lower accum block.
input	CLK;	         // Clock for MAC16 elements 
input	CE;              // Clock enable . global control 
input	IRSTTOP;         // Active High  reset for  A,C registers,upper half multplier pipeline regs(16). 
input	IRSTBOT;         // Active High reset for  B,D registers, lower half multiplier pipeline regs(16), 32 bit result pipelines regs   
input	ORSTTOP;	 // Active High reset for top accum registers O[31:16]
input	ORSTBOT;         // Active High reset for bottom accum registers O[15:0]   
input   AHOLD;           // Active High hold data signal for A register
input   BHOLD;           // Active High hold data signal for B register   
input   CHOLD;           // Active High hold data signal for C register
input   DHOLD;           // Active High hold data signal for D register 
input   OHOLDTOP;        // Active High hold data signal for top accum registers O[31:16]
input   OHOLDBOT;        // Active High hold data signal for bottom  accum registers O[15:0]     
input 	OLOADTOP;        // Load top accum regiser with  direct input C or Registered data C.  
input 	OLOADBOT;        // Load bottom accum regisers with direct input D or Registered data D
input 	ADDSUBTOP;       // Control for Add/Sub operation for top accum . 0-addition , 1-subtraction.  
input 	ADDSUBBOT;       // Control for Add/Sub operation for bottom accum . 0-addition , 1-subtraction.
output  CO;              // top accumulator carry out to next LUT
input 	CI;              // bottom accumaltor carry in signal from lower LUT block. 
input   ACCUMCI;         // Carry in from  MAC16 below
output  ACCUMCO;         // Carry out to MAC16 above
input   SIGNEXTIN;	 // Single bit Sign extenstion from MAC16 below         
output  SIGNEXTOUT;      // Single bit Sign extenstion to MAC16 above


parameter NEG_TRIGGER = 1'b0;    
parameter C_REG = 1'b0;     			// C0
parameter A_REG = 1'b0;     			// C1
parameter B_REG = 1'b0;     			// C2
parameter D_REG = 1'b0;     			// C3

parameter TOP_8x8_MULT_REG = 1'b0; 		//C4
parameter BOT_8x8_MULT_REG = 1'b0; 		//C5
parameter PIPELINE_16x16_MULT_REG1 = 1'b0; 	//C6
parameter PIPELINE_16x16_MULT_REG2 = 1'b0; 	//C7

parameter TOPOUTPUT_SELECT =  2'b00; 		//COMB, ACCUM_REG, MULT_8x8, MULT_16x16  // {C9,C8} = 00, 01, 10, 11
parameter TOPADDSUB_LOWERINPUT = 2'b00; 	//DATA, MULT_8x8, MULT_16x16, SIGNEXT    // {C11,C10} = 00, 01, 10, 11
parameter TOPADDSUB_UPPERINPUT = 1'b0; 		//ACCUM_REG, DATAC  			 //  C12 = 0, 1
parameter TOPADDSUB_CARRYSELECT = 2'b00; 	//LOGIC0, LOGIC1, LCOCAS, GENERATED_CARRY (LCO) // {C14, C13} = 00, 01, 10, 11

parameter BOTOUTPUT_SELECT =  2'b00; 		//COMB, ACCUM_REG, MULT_8x8, MULT_16x16   // {C16,C15} = 00, 01, 10, 11
parameter BOTADDSUB_LOWERINPUT = 2'b00; 	//DATA, MULT_8x8, MULT_16x16, SIGNEXTIN   // {C18,C17} = 00, 01, 10, 11
parameter BOTADDSUB_UPPERINPUT = 1'b0;  	//ACCUM_REG, DATAD   			  // C19 = 0, 1
parameter BOTADDSUB_CARRYSELECT = 2'b00; 	//LOGIC0, LOGIC1, ACCUMCI, CI  		  // {C21, C20} = 00, 01, 10, 11
parameter MODE_8x8 = 1'b0; 			// C22 

parameter A_SIGNED = 1'b0;  			// C23
parameter B_SIGNED = 1'b0;  			// C24	 

//--------- local params ----------------------------------------------------// 
localparam cbits_inreg   	= {D_REG,B_REG,A_REG,C_REG}; 
localparam cbits_mpyreg   	= {PIPELINE_16x16_MULT_REG2,PIPELINE_16x16_MULT_REG1,BOT_8x8_MULT_REG,TOP_8x8_MULT_REG};
localparam cbits_topmac	 	= {TOPADDSUB_CARRYSELECT,TOPADDSUB_UPPERINPUT,TOPADDSUB_LOWERINPUT,TOPOUTPUT_SELECT};
localparam cbits_botmac	 	= {BOTADDSUB_CARRYSELECT,BOTADDSUB_UPPERINPUT,BOTADDSUB_LOWERINPUT,BOTOUTPUT_SELECT};
localparam cbits_sign	 	= {B_SIGNED,A_SIGNED,MODE_8x8}; 
localparam cbits 	  	= {cbits_sign,cbits_botmac,cbits_topmac,cbits_mpyreg,cbits_inreg}; 

wire CLK_g , intCLK; 
reg NOTIFIER;


//------------------- initial block --------------------------------------// 
	
	initial 
begin 
	
	
	
	if( (TOPOUTPUT_SELECT != 2'b00 )&& (TOPOUTPUT_SELECT != 2'b01 ) && (TOPOUTPUT_SELECT != 2'b10 ) && (TOPOUTPUT_SELECT !=2'b11 ) ) begin 
	$display("Error: TOPOUTPUT_SELECT parameter is set to incorrect value. Exiting Simulation ...."); 
	$finish;	
	end 
	if( (TOPADDSUB_LOWERINPUT != 2'b00) && (TOPADDSUB_LOWERINPUT != 2'b01) && (TOPADDSUB_LOWERINPUT != 2'b10) && (TOPADDSUB_LOWERINPUT != 2'b11) ) begin 
	$display("Error: TOPADDSUB_LOWERINPUT parameter is set to incorrect value. Exiting Simulation ...."); 
	$finish; 
	end 
	if( (TOPADDSUB_UPPERINPUT != 1'b0 ) && (TOPADDSUB_UPPERINPUT != 1'b1) ) begin
	$display("Error: TOPADDSUB_UPPERINPUT parameter is set to incorrect value. Exiting Simulation ....");
        $finish;
        end
	if( (TOPADDSUB_CARRYSELECT != 2'b00 )&&(TOPADDSUB_CARRYSELECT != 2'b01) && (TOPADDSUB_CARRYSELECT != 2'b10) &&(TOPADDSUB_CARRYSELECT != 2'b11)) begin 
	$display("Error: TOPADDSUB_CARRYSELECT parameter is set to incorrect value. Exiting Simulation ....");
        $finish;
        end

	
	if( (BOTOUTPUT_SELECT != 2'b00 )&& (BOTOUTPUT_SELECT != 2'b01 ) && (BOTOUTPUT_SELECT != 2'b10 ) && (BOTOUTPUT_SELECT !=2'b11 ) ) begin 
	$display("Error: BOTOUTPUT_SELECT parameter is set to incorrect value. Exiting Simulation ...."); 
	$finish;	
	end 
	if( (BOTADDSUB_LOWERINPUT != 2'b00) && (BOTADDSUB_LOWERINPUT != 2'b01) && (BOTADDSUB_LOWERINPUT != 2'b10) && (BOTADDSUB_LOWERINPUT != 2'b11) ) begin 
	$display("Error: BOTADDSUB_LOWERINPUT parameter is set to incorrect value. Exiting Simulation ...."); 
	$finish; 
	end 
	if( (BOTADDSUB_UPPERINPUT != 1'b0 ) && (BOTADDSUB_UPPERINPUT != 1'b1) ) begin
	$display("Error:BOTADDSUB_UPPERINPUT parameter is set to incorrect value. Exiting Simulation ....");
        $finish;
        end
	if( (BOTADDSUB_CARRYSELECT != 2'b00 ) && (BOTADDSUB_CARRYSELECT != 2'b01) && (BOTADDSUB_CARRYSELECT != 2'b10) && (BOTADDSUB_CARRYSELECT != 2'b11)) begin 
	$display("Error: BOTADDSUB_CARRYSELECT parameter is set to incorrect value. Exiting Simulation ....");
        $finish;
        end
	
	//Validation for mode8x8.
		if (PIPELINE_16x16_MULT_REG1 == 1'b1 || PIPELINE_16x16_MULT_REG2 ==1'b1 ) begin   		
		$display ("**************  INFO  ***********************************"); 
		$display ("Info : To Reset 16x16 multiplier INTERNAL PIPELINE REGISTER assert both IRSTTOP and IRSTBOT signals") ;  
	        $display ("Info : To Reset 16x16 multiplier OUTPUT  REGISTER   assert IRSTBOT signal");  	
		$display ("**********************************************************"); 	
		end else if ( (PIPELINE_16x16_MULT_REG1 == 1'b1 || PIPELINE_16x16_MULT_REG2 ==1'b1) &&  MODE_8x8 == 1'b1) begin
		  
		$display ("***********  ERROR  ****************************************"); 
		$display ("Error : MODE_8x8 parameter is set to 1. To use 16x16 mulitplier internal and output registers it should be set to 0.Exiting Simulation ...."); 
		
		$display ("***************************************************************"); 	
		$finish; 
		end else if( (PIPELINE_16x16_MULT_REG1 == 1'b0 &&  PIPELINE_16x16_MULT_REG2 ==1'b0)  &&  MODE_8x8 == 1'b0 ) begin
                $display ("************ WARNING  **********************************************");
                $display ("Warning : When 16x16 multiplier PIPELINE REGISTERS are not used, set MODE_8x8 to 1(power save mode) ");
                $display ("*******************************************************************");
		end 


end	// initial  

//-------------------------- Default input signals -------------------------------------// 
assign (weak0,weak1) CE 	= 1'b1; 
assign (weak0,weak1) A  	= 16'b0; 
assign (weak0,weak1) B  	= 16'b0; 
assign (weak0,weak1) C  	= 16'b0; 
assign (weak0,weak1) D  	= 16'b0; 
assign (weak0,weak1) AHOLD 	= 1'b0; 
assign (weak0,weak1) BHOLD 	= 1'b0; 
assign (weak0,weak1) CHOLD 	= 1'b0; 
assign (weak0,weak1) DHOLD    	= 1'b0; 
assign (weak0,weak1) IRSTTOP  	= 1'b0; 
assign (weak0,weak1) IRSTBOT  	= 1'b0; 
assign (weak0,weak1) ORSTTOP  	= 1'b0; 
assign (weak0,weak1) ORSTBOT  	= 1'b0; 
assign (weak0,weak1) OLOADTOP 	= 1'b0; 
assign (weak0,weak1) OLOADBOT 	= 1'b0; 
assign (weak0,weak1) ADDSUBTOP	= 1'b0; 
assign (weak0,weak1) ADDSUBBOT  = 1'b0; 
assign (weak0,weak1) OHOLDTOP   = 1'b0; 
assign (weak0,weak1) OHOLDBOT	= 1'b0;   
assign (weak0,weak1) CI		= 1'b0;   
assign (weak0,weak1) ACCUMCI	= 1'b0;   


//---------------------------Logic section --------------------------------------------// 

assign CLK_g = (CLK & CE);  				// CE=0 disables entire clock  
assign intCLK = (CLK_g ^ NEG_TRIGGER);			// Clock Polarity control 

 mac16_physical  mac16physical_i (
	 .CLK(intCLK) ,
	 .A(A) ,
	 .B(B) ,
	 .C(C) ,
	 .D(D) ,
	 .IHRST(IRSTTOP),
	 .ILRST(IRSTBOT),
	 .OHRST(ORSTTOP),
	 .OLRST(ORSTBOT),
	 .AHLD(AHOLD),
	 .BHLD(BHOLD),
	 .CHLD(CHOLD),
	 .DHLD(DHOLD),
		
	 .OHHLD(OHOLDTOP),
	 .OLHLD(OHOLDBOT),
	 .OHADS(ADDSUBTOP),
	 .OLADS(ADDSUBBOT),
	 .OHLDA(OLOADTOP),
	 .OLLDA(OLOADBOT),
	 .CICAS(ACCUMCI),
	 .CI(CI),
	 .SIGNEXTIN(SIGNEXTIN),
	 .SIGNEXTOUT(SIGNEXTOUT),
	 .COCAS(ACCUMCO),
	 .CO(CO),
	 .O(O), 
	 .CBIT(cbits)
    );
`ifdef TIMINGCHECK		
specify


		 (A[0] *> O[0])=(0.0,0.0); 
        (A[0] *> O[1])=(0.0,0.0); 
        (A[0] *> O[2])=(0.0,0.0); 
        (A[0] *> O[3])=(0.0,0.0); 
        (A[0] *> O[4])=(0.0,0.0); 
        (A[0] *> O[5])=(0.0,0.0); 
        (A[0] *> O[6])=(0.0,0.0); 
        (A[0] *> O[7])=(0.0,0.0); 
        (A[0] *> O[8])=(0.0,0.0); 
        (A[0] *> O[9])=(0.0,0.0); 
        (A[0] *> O[10])=(0.0,0.0); 
        (A[0] *> O[11])=(0.0,0.0); 
        (A[0] *> O[12])=(0.0,0.0); 
        (A[0] *> O[13])=(0.0,0.0); 
        (A[0] *> O[14])=(0.0,0.0); 
        (A[0] *> O[15])=(0.0,0.0); 
        (A[0] *> O[16])=(0.0,0.0); 
        (A[0] *> O[17])=(0.0,0.0); 
        (A[0] *> O[18])=(0.0,0.0); 
        (A[0] *> O[19])=(0.0,0.0); 
        (A[0] *> O[20])=(0.0,0.0); 
        (A[0] *> O[21])=(0.0,0.0); 
        (A[0] *> O[22])=(0.0,0.0); 
        (A[0] *> O[23])=(0.0,0.0); 
        (A[0] *> O[24])=(0.0,0.0); 
        (A[0] *> O[25])=(0.0,0.0); 
        (A[0] *> O[26])=(0.0,0.0); 
        (A[0] *> O[27])=(0.0,0.0); 
        (A[0] *> O[28])=(0.0,0.0); 
        (A[0] *> O[29])=(0.0,0.0); 
        (A[0] *> O[30])=(0.0,0.0); 
        (A[0] *> O[31])=(0.0,0.0); 
        (A[1] *> O[0])=(0.0,0.0); 
        (A[1] *> O[1])=(0.0,0.0); 
        (A[1] *> O[2])=(0.0,0.0); 
        (A[1] *> O[3])=(0.0,0.0); 
        (A[1] *> O[4])=(0.0,0.0); 
        (A[1] *> O[5])=(0.0,0.0); 
        (A[1] *> O[6])=(0.0,0.0); 
        (A[1] *> O[7])=(0.0,0.0); 
        (A[1] *> O[8])=(0.0,0.0); 
        (A[1] *> O[9])=(0.0,0.0); 
        (A[1] *> O[10])=(0.0,0.0); 
        (A[1] *> O[11])=(0.0,0.0); 
        (A[1] *> O[12])=(0.0,0.0); 
        (A[1] *> O[13])=(0.0,0.0); 
        (A[1] *> O[14])=(0.0,0.0); 
        (A[1] *> O[15])=(0.0,0.0); 
        (A[1] *> O[16])=(0.0,0.0); 
        (A[1] *> O[17])=(0.0,0.0); 
        (A[1] *> O[18])=(0.0,0.0); 
        (A[1] *> O[19])=(0.0,0.0); 
        (A[1] *> O[20])=(0.0,0.0); 
        (A[1] *> O[21])=(0.0,0.0); 
        (A[1] *> O[22])=(0.0,0.0); 
        (A[1] *> O[23])=(0.0,0.0); 
        (A[1] *> O[24])=(0.0,0.0); 
        (A[1] *> O[25])=(0.0,0.0); 
        (A[1] *> O[26])=(0.0,0.0); 
        (A[1] *> O[27])=(0.0,0.0); 
        (A[1] *> O[28])=(0.0,0.0); 
        (A[1] *> O[29])=(0.0,0.0); 
        (A[1] *> O[30])=(0.0,0.0); 
        (A[1] *> O[31])=(0.0,0.0); 
        (A[2] *> O[0])=(0.0,0.0); 
        (A[2] *> O[1])=(0.0,0.0); 
        (A[2] *> O[2])=(0.0,0.0); 
        (A[2] *> O[3])=(0.0,0.0); 
        (A[2] *> O[4])=(0.0,0.0); 
        (A[2] *> O[5])=(0.0,0.0); 
        (A[2] *> O[6])=(0.0,0.0); 
        (A[2] *> O[7])=(0.0,0.0); 
        (A[2] *> O[8])=(0.0,0.0); 
        (A[2] *> O[9])=(0.0,0.0); 
        (A[2] *> O[10])=(0.0,0.0); 
        (A[2] *> O[11])=(0.0,0.0); 
        (A[2] *> O[12])=(0.0,0.0); 
        (A[2] *> O[13])=(0.0,0.0); 
        (A[2] *> O[14])=(0.0,0.0); 
        (A[2] *> O[15])=(0.0,0.0); 
        (A[2] *> O[16])=(0.0,0.0); 
        (A[2] *> O[17])=(0.0,0.0); 
        (A[2] *> O[18])=(0.0,0.0); 
        (A[2] *> O[19])=(0.0,0.0); 
        (A[2] *> O[20])=(0.0,0.0); 
        (A[2] *> O[21])=(0.0,0.0); 
        (A[2] *> O[22])=(0.0,0.0); 
        (A[2] *> O[23])=(0.0,0.0); 
        (A[2] *> O[24])=(0.0,0.0); 
        (A[2] *> O[25])=(0.0,0.0); 
        (A[2] *> O[26])=(0.0,0.0); 
        (A[2] *> O[27])=(0.0,0.0); 
        (A[2] *> O[28])=(0.0,0.0); 
        (A[2] *> O[29])=(0.0,0.0); 
        (A[2] *> O[30])=(0.0,0.0); 
        (A[2] *> O[31])=(0.0,0.0); 
        (A[3] *> O[0])=(0.0,0.0); 
        (A[3] *> O[1])=(0.0,0.0); 
        (A[3] *> O[2])=(0.0,0.0); 
        (A[3] *> O[3])=(0.0,0.0); 
        (A[3] *> O[4])=(0.0,0.0); 
        (A[3] *> O[5])=(0.0,0.0); 
        (A[3] *> O[6])=(0.0,0.0); 
        (A[3] *> O[7])=(0.0,0.0); 
        (A[3] *> O[8])=(0.0,0.0); 
        (A[3] *> O[9])=(0.0,0.0); 
        (A[3] *> O[10])=(0.0,0.0); 
        (A[3] *> O[11])=(0.0,0.0); 
        (A[3] *> O[12])=(0.0,0.0); 
        (A[3] *> O[13])=(0.0,0.0); 
        (A[3] *> O[14])=(0.0,0.0); 
        (A[3] *> O[15])=(0.0,0.0); 
        (A[3] *> O[16])=(0.0,0.0); 
        (A[3] *> O[17])=(0.0,0.0); 
        (A[3] *> O[18])=(0.0,0.0); 
        (A[3] *> O[19])=(0.0,0.0); 
        (A[3] *> O[20])=(0.0,0.0); 
        (A[3] *> O[21])=(0.0,0.0); 
        (A[3] *> O[22])=(0.0,0.0); 
        (A[3] *> O[23])=(0.0,0.0); 
        (A[3] *> O[24])=(0.0,0.0); 
        (A[3] *> O[25])=(0.0,0.0); 
        (A[3] *> O[26])=(0.0,0.0); 
        (A[3] *> O[27])=(0.0,0.0); 
        (A[3] *> O[28])=(0.0,0.0); 
        (A[3] *> O[29])=(0.0,0.0); 
        (A[3] *> O[30])=(0.0,0.0); 
        (A[3] *> O[31])=(0.0,0.0); 
        (A[4] *> O[0])=(0.0,0.0); 
        (A[4] *> O[1])=(0.0,0.0); 
        (A[4] *> O[2])=(0.0,0.0); 
        (A[4] *> O[3])=(0.0,0.0); 
        (A[4] *> O[4])=(0.0,0.0); 
        (A[4] *> O[5])=(0.0,0.0); 
        (A[4] *> O[6])=(0.0,0.0); 
        (A[4] *> O[7])=(0.0,0.0); 
        (A[4] *> O[8])=(0.0,0.0); 
        (A[4] *> O[9])=(0.0,0.0); 
        (A[4] *> O[10])=(0.0,0.0); 
        (A[4] *> O[11])=(0.0,0.0); 
        (A[4] *> O[12])=(0.0,0.0); 
        (A[4] *> O[13])=(0.0,0.0); 
        (A[4] *> O[14])=(0.0,0.0); 
        (A[4] *> O[15])=(0.0,0.0); 
        (A[4] *> O[16])=(0.0,0.0); 
        (A[4] *> O[17])=(0.0,0.0); 
        (A[4] *> O[18])=(0.0,0.0); 
        (A[4] *> O[19])=(0.0,0.0); 
        (A[4] *> O[20])=(0.0,0.0); 
        (A[4] *> O[21])=(0.0,0.0); 
        (A[4] *> O[22])=(0.0,0.0); 
        (A[4] *> O[23])=(0.0,0.0); 
        (A[4] *> O[24])=(0.0,0.0); 
        (A[4] *> O[25])=(0.0,0.0); 
        (A[4] *> O[26])=(0.0,0.0); 
        (A[4] *> O[27])=(0.0,0.0); 
        (A[4] *> O[28])=(0.0,0.0); 
        (A[4] *> O[29])=(0.0,0.0); 
        (A[4] *> O[30])=(0.0,0.0); 
        (A[4] *> O[31])=(0.0,0.0); 
        (A[5] *> O[0])=(0.0,0.0); 
        (A[5] *> O[1])=(0.0,0.0); 
        (A[5] *> O[2])=(0.0,0.0); 
        (A[5] *> O[3])=(0.0,0.0); 
        (A[5] *> O[4])=(0.0,0.0); 
        (A[5] *> O[5])=(0.0,0.0); 
        (A[5] *> O[6])=(0.0,0.0); 
        (A[5] *> O[7])=(0.0,0.0); 
        (A[5] *> O[8])=(0.0,0.0); 
        (A[5] *> O[9])=(0.0,0.0); 
        (A[5] *> O[10])=(0.0,0.0); 
        (A[5] *> O[11])=(0.0,0.0); 
        (A[5] *> O[12])=(0.0,0.0); 
        (A[5] *> O[13])=(0.0,0.0); 
        (A[5] *> O[14])=(0.0,0.0); 
        (A[5] *> O[15])=(0.0,0.0); 
        (A[5] *> O[16])=(0.0,0.0); 
        (A[5] *> O[17])=(0.0,0.0); 
        (A[5] *> O[18])=(0.0,0.0); 
        (A[5] *> O[19])=(0.0,0.0); 
        (A[5] *> O[20])=(0.0,0.0); 
        (A[5] *> O[21])=(0.0,0.0); 
        (A[5] *> O[22])=(0.0,0.0); 
        (A[5] *> O[23])=(0.0,0.0); 
        (A[5] *> O[24])=(0.0,0.0); 
        (A[5] *> O[25])=(0.0,0.0); 
        (A[5] *> O[26])=(0.0,0.0); 
        (A[5] *> O[27])=(0.0,0.0); 
        (A[5] *> O[28])=(0.0,0.0); 
        (A[5] *> O[29])=(0.0,0.0); 
        (A[5] *> O[30])=(0.0,0.0); 
        (A[5] *> O[31])=(0.0,0.0); 
        (A[6] *> O[0])=(0.0,0.0); 
        (A[6] *> O[1])=(0.0,0.0); 
        (A[6] *> O[2])=(0.0,0.0); 
        (A[6] *> O[3])=(0.0,0.0); 
        (A[6] *> O[4])=(0.0,0.0); 
        (A[6] *> O[5])=(0.0,0.0); 
        (A[6] *> O[6])=(0.0,0.0); 
        (A[6] *> O[7])=(0.0,0.0); 
        (A[6] *> O[8])=(0.0,0.0); 
        (A[6] *> O[9])=(0.0,0.0); 
        (A[6] *> O[10])=(0.0,0.0); 
        (A[6] *> O[11])=(0.0,0.0); 
        (A[6] *> O[12])=(0.0,0.0); 
        (A[6] *> O[13])=(0.0,0.0); 
        (A[6] *> O[14])=(0.0,0.0); 
        (A[6] *> O[15])=(0.0,0.0); 
        (A[6] *> O[16])=(0.0,0.0); 
        (A[6] *> O[17])=(0.0,0.0); 
        (A[6] *> O[18])=(0.0,0.0); 
        (A[6] *> O[19])=(0.0,0.0); 
        (A[6] *> O[20])=(0.0,0.0); 
        (A[6] *> O[21])=(0.0,0.0); 
        (A[6] *> O[22])=(0.0,0.0); 
        (A[6] *> O[23])=(0.0,0.0); 
        (A[6] *> O[24])=(0.0,0.0); 
        (A[6] *> O[25])=(0.0,0.0); 
        (A[6] *> O[26])=(0.0,0.0); 
        (A[6] *> O[27])=(0.0,0.0); 
        (A[6] *> O[28])=(0.0,0.0); 
        (A[6] *> O[29])=(0.0,0.0); 
        (A[6] *> O[30])=(0.0,0.0); 
        (A[6] *> O[31])=(0.0,0.0); 
        (A[7] *> O[0])=(0.0,0.0); 
        (A[7] *> O[1])=(0.0,0.0); 
        (A[7] *> O[2])=(0.0,0.0); 
        (A[7] *> O[3])=(0.0,0.0); 
        (A[7] *> O[4])=(0.0,0.0); 
        (A[7] *> O[5])=(0.0,0.0); 
        (A[7] *> O[6])=(0.0,0.0); 
        (A[7] *> O[7])=(0.0,0.0); 
        (A[7] *> O[8])=(0.0,0.0); 
        (A[7] *> O[9])=(0.0,0.0); 
        (A[7] *> O[10])=(0.0,0.0); 
        (A[7] *> O[11])=(0.0,0.0); 
        (A[7] *> O[12])=(0.0,0.0); 
        (A[7] *> O[13])=(0.0,0.0); 
        (A[7] *> O[14])=(0.0,0.0); 
        (A[7] *> O[15])=(0.0,0.0); 
        (A[7] *> O[16])=(0.0,0.0); 
        (A[7] *> O[17])=(0.0,0.0); 
        (A[7] *> O[18])=(0.0,0.0); 
        (A[7] *> O[19])=(0.0,0.0); 
        (A[7] *> O[20])=(0.0,0.0); 
        (A[7] *> O[21])=(0.0,0.0); 
        (A[7] *> O[22])=(0.0,0.0); 
        (A[7] *> O[23])=(0.0,0.0); 
        (A[7] *> O[24])=(0.0,0.0); 
        (A[7] *> O[25])=(0.0,0.0); 
        (A[7] *> O[26])=(0.0,0.0); 
        (A[7] *> O[27])=(0.0,0.0); 
        (A[7] *> O[28])=(0.0,0.0); 
        (A[7] *> O[29])=(0.0,0.0); 
        (A[7] *> O[30])=(0.0,0.0); 
        (A[7] *> O[31])=(0.0,0.0); 
        (A[8] *> O[0])=(0.0,0.0); 
        (A[8] *> O[1])=(0.0,0.0); 
        (A[8] *> O[2])=(0.0,0.0); 
        (A[8] *> O[3])=(0.0,0.0); 
        (A[8] *> O[4])=(0.0,0.0); 
        (A[8] *> O[5])=(0.0,0.0); 
        (A[8] *> O[6])=(0.0,0.0); 
        (A[8] *> O[7])=(0.0,0.0); 
        (A[8] *> O[8])=(0.0,0.0); 
        (A[8] *> O[9])=(0.0,0.0); 
        (A[8] *> O[10])=(0.0,0.0); 
        (A[8] *> O[11])=(0.0,0.0); 
        (A[8] *> O[12])=(0.0,0.0); 
        (A[8] *> O[13])=(0.0,0.0); 
        (A[8] *> O[14])=(0.0,0.0); 
        (A[8] *> O[15])=(0.0,0.0); 
        (A[8] *> O[16])=(0.0,0.0); 
        (A[8] *> O[17])=(0.0,0.0); 
        (A[8] *> O[18])=(0.0,0.0); 
        (A[8] *> O[19])=(0.0,0.0); 
        (A[8] *> O[20])=(0.0,0.0); 
        (A[8] *> O[21])=(0.0,0.0); 
        (A[8] *> O[22])=(0.0,0.0); 
        (A[8] *> O[23])=(0.0,0.0); 
        (A[8] *> O[24])=(0.0,0.0); 
        (A[8] *> O[25])=(0.0,0.0); 
        (A[8] *> O[26])=(0.0,0.0); 
        (A[8] *> O[27])=(0.0,0.0); 
        (A[8] *> O[28])=(0.0,0.0); 
        (A[8] *> O[29])=(0.0,0.0); 
        (A[8] *> O[30])=(0.0,0.0); 
        (A[8] *> O[31])=(0.0,0.0); 
        (A[9] *> O[0])=(0.0,0.0); 
        (A[9] *> O[1])=(0.0,0.0); 
        (A[9] *> O[2])=(0.0,0.0); 
        (A[9] *> O[3])=(0.0,0.0); 
        (A[9] *> O[4])=(0.0,0.0); 
        (A[9] *> O[5])=(0.0,0.0); 
        (A[9] *> O[6])=(0.0,0.0); 
        (A[9] *> O[7])=(0.0,0.0); 
        (A[9] *> O[8])=(0.0,0.0); 
        (A[9] *> O[9])=(0.0,0.0); 
        (A[9] *> O[10])=(0.0,0.0); 
        (A[9] *> O[11])=(0.0,0.0); 
        (A[9] *> O[12])=(0.0,0.0); 
        (A[9] *> O[13])=(0.0,0.0); 
        (A[9] *> O[14])=(0.0,0.0); 
        (A[9] *> O[15])=(0.0,0.0); 
        (A[9] *> O[16])=(0.0,0.0); 
        (A[9] *> O[17])=(0.0,0.0); 
        (A[9] *> O[18])=(0.0,0.0); 
        (A[9] *> O[19])=(0.0,0.0); 
        (A[9] *> O[20])=(0.0,0.0); 
        (A[9] *> O[21])=(0.0,0.0); 
        (A[9] *> O[22])=(0.0,0.0); 
        (A[9] *> O[23])=(0.0,0.0); 
        (A[9] *> O[24])=(0.0,0.0); 
        (A[9] *> O[25])=(0.0,0.0); 
        (A[9] *> O[26])=(0.0,0.0); 
        (A[9] *> O[27])=(0.0,0.0); 
        (A[9] *> O[28])=(0.0,0.0); 
        (A[9] *> O[29])=(0.0,0.0); 
        (A[9] *> O[30])=(0.0,0.0); 
        (A[9] *> O[31])=(0.0,0.0); 
        (A[10] *> O[0])=(0.0,0.0); 
        (A[10] *> O[1])=(0.0,0.0); 
        (A[10] *> O[2])=(0.0,0.0); 
        (A[10] *> O[3])=(0.0,0.0); 
        (A[10] *> O[4])=(0.0,0.0); 
        (A[10] *> O[5])=(0.0,0.0); 
        (A[10] *> O[6])=(0.0,0.0); 
        (A[10] *> O[7])=(0.0,0.0); 
        (A[10] *> O[8])=(0.0,0.0); 
        (A[10] *> O[9])=(0.0,0.0); 
        (A[10] *> O[10])=(0.0,0.0); 
        (A[10] *> O[11])=(0.0,0.0); 
        (A[10] *> O[12])=(0.0,0.0); 
        (A[10] *> O[13])=(0.0,0.0); 
        (A[10] *> O[14])=(0.0,0.0); 
        (A[10] *> O[15])=(0.0,0.0); 
        (A[10] *> O[16])=(0.0,0.0); 
        (A[10] *> O[17])=(0.0,0.0); 
        (A[10] *> O[18])=(0.0,0.0); 
        (A[10] *> O[19])=(0.0,0.0); 
        (A[10] *> O[20])=(0.0,0.0); 
        (A[10] *> O[21])=(0.0,0.0); 
        (A[10] *> O[22])=(0.0,0.0); 
        (A[10] *> O[23])=(0.0,0.0); 
        (A[10] *> O[24])=(0.0,0.0); 
        (A[10] *> O[25])=(0.0,0.0); 
        (A[10] *> O[26])=(0.0,0.0); 
        (A[10] *> O[27])=(0.0,0.0); 
        (A[10] *> O[28])=(0.0,0.0); 
        (A[10] *> O[29])=(0.0,0.0); 
        (A[10] *> O[30])=(0.0,0.0); 
        (A[10] *> O[31])=(0.0,0.0); 
        (A[11] *> O[0])=(0.0,0.0); 
        (A[11] *> O[1])=(0.0,0.0); 
        (A[11] *> O[2])=(0.0,0.0); 
        (A[11] *> O[3])=(0.0,0.0); 
        (A[11] *> O[4])=(0.0,0.0); 
        (A[11] *> O[5])=(0.0,0.0); 
        (A[11] *> O[6])=(0.0,0.0); 
        (A[11] *> O[7])=(0.0,0.0); 
        (A[11] *> O[8])=(0.0,0.0); 
        (A[11] *> O[9])=(0.0,0.0); 
        (A[11] *> O[10])=(0.0,0.0); 
        (A[11] *> O[11])=(0.0,0.0); 
        (A[11] *> O[12])=(0.0,0.0); 
        (A[11] *> O[13])=(0.0,0.0); 
        (A[11] *> O[14])=(0.0,0.0); 
        (A[11] *> O[15])=(0.0,0.0); 
        (A[11] *> O[16])=(0.0,0.0); 
        (A[11] *> O[17])=(0.0,0.0); 
        (A[11] *> O[18])=(0.0,0.0); 
        (A[11] *> O[19])=(0.0,0.0); 
        (A[11] *> O[20])=(0.0,0.0); 
        (A[11] *> O[21])=(0.0,0.0); 
        (A[11] *> O[22])=(0.0,0.0); 
        (A[11] *> O[23])=(0.0,0.0); 
        (A[11] *> O[24])=(0.0,0.0); 
        (A[11] *> O[25])=(0.0,0.0); 
        (A[11] *> O[26])=(0.0,0.0); 
        (A[11] *> O[27])=(0.0,0.0); 
        (A[11] *> O[28])=(0.0,0.0); 
        (A[11] *> O[29])=(0.0,0.0); 
        (A[11] *> O[30])=(0.0,0.0); 
        (A[11] *> O[31])=(0.0,0.0); 
        (A[12] *> O[0])=(0.0,0.0); 
        (A[12] *> O[1])=(0.0,0.0); 
        (A[12] *> O[2])=(0.0,0.0); 
        (A[12] *> O[3])=(0.0,0.0); 
        (A[12] *> O[4])=(0.0,0.0); 
        (A[12] *> O[5])=(0.0,0.0); 
        (A[12] *> O[6])=(0.0,0.0); 
        (A[12] *> O[7])=(0.0,0.0); 
        (A[12] *> O[8])=(0.0,0.0); 
        (A[12] *> O[9])=(0.0,0.0); 
        (A[12] *> O[10])=(0.0,0.0); 
        (A[12] *> O[11])=(0.0,0.0); 
        (A[12] *> O[12])=(0.0,0.0); 
        (A[12] *> O[13])=(0.0,0.0); 
        (A[12] *> O[14])=(0.0,0.0); 
        (A[12] *> O[15])=(0.0,0.0); 
        (A[12] *> O[16])=(0.0,0.0); 
        (A[12] *> O[17])=(0.0,0.0); 
        (A[12] *> O[18])=(0.0,0.0); 
        (A[12] *> O[19])=(0.0,0.0); 
        (A[12] *> O[20])=(0.0,0.0); 
        (A[12] *> O[21])=(0.0,0.0); 
        (A[12] *> O[22])=(0.0,0.0); 
        (A[12] *> O[23])=(0.0,0.0); 
        (A[12] *> O[24])=(0.0,0.0); 
        (A[12] *> O[25])=(0.0,0.0); 
        (A[12] *> O[26])=(0.0,0.0); 
        (A[12] *> O[27])=(0.0,0.0); 
        (A[12] *> O[28])=(0.0,0.0); 
        (A[12] *> O[29])=(0.0,0.0); 
        (A[12] *> O[30])=(0.0,0.0); 
        (A[12] *> O[31])=(0.0,0.0); 
        (A[13] *> O[0])=(0.0,0.0); 
        (A[13] *> O[1])=(0.0,0.0); 
        (A[13] *> O[2])=(0.0,0.0); 
        (A[13] *> O[3])=(0.0,0.0); 
        (A[13] *> O[4])=(0.0,0.0); 
        (A[13] *> O[5])=(0.0,0.0); 
        (A[13] *> O[6])=(0.0,0.0); 
        (A[13] *> O[7])=(0.0,0.0); 
        (A[13] *> O[8])=(0.0,0.0); 
        (A[13] *> O[9])=(0.0,0.0); 
        (A[13] *> O[10])=(0.0,0.0); 
        (A[13] *> O[11])=(0.0,0.0); 
        (A[13] *> O[12])=(0.0,0.0); 
        (A[13] *> O[13])=(0.0,0.0); 
        (A[13] *> O[14])=(0.0,0.0); 
        (A[13] *> O[15])=(0.0,0.0); 
        (A[13] *> O[16])=(0.0,0.0); 
        (A[13] *> O[17])=(0.0,0.0); 
        (A[13] *> O[18])=(0.0,0.0); 
        (A[13] *> O[19])=(0.0,0.0); 
        (A[13] *> O[20])=(0.0,0.0); 
        (A[13] *> O[21])=(0.0,0.0); 
        (A[13] *> O[22])=(0.0,0.0); 
        (A[13] *> O[23])=(0.0,0.0); 
        (A[13] *> O[24])=(0.0,0.0); 
        (A[13] *> O[25])=(0.0,0.0); 
        (A[13] *> O[26])=(0.0,0.0); 
        (A[13] *> O[27])=(0.0,0.0); 
        (A[13] *> O[28])=(0.0,0.0); 
        (A[13] *> O[29])=(0.0,0.0); 
        (A[13] *> O[30])=(0.0,0.0); 
        (A[13] *> O[31])=(0.0,0.0); 
        (A[14] *> O[0])=(0.0,0.0); 
        (A[14] *> O[1])=(0.0,0.0); 
        (A[14] *> O[2])=(0.0,0.0); 
        (A[14] *> O[3])=(0.0,0.0); 
        (A[14] *> O[4])=(0.0,0.0); 
        (A[14] *> O[5])=(0.0,0.0); 
        (A[14] *> O[6])=(0.0,0.0); 
        (A[14] *> O[7])=(0.0,0.0); 
        (A[14] *> O[8])=(0.0,0.0); 
        (A[14] *> O[9])=(0.0,0.0); 
        (A[14] *> O[10])=(0.0,0.0); 
        (A[14] *> O[11])=(0.0,0.0); 
        (A[14] *> O[12])=(0.0,0.0); 
        (A[14] *> O[13])=(0.0,0.0); 
        (A[14] *> O[14])=(0.0,0.0); 
        (A[14] *> O[15])=(0.0,0.0); 
        (A[14] *> O[16])=(0.0,0.0); 
        (A[14] *> O[17])=(0.0,0.0); 
        (A[14] *> O[18])=(0.0,0.0); 
        (A[14] *> O[19])=(0.0,0.0); 
        (A[14] *> O[20])=(0.0,0.0); 
        (A[14] *> O[21])=(0.0,0.0); 
        (A[14] *> O[22])=(0.0,0.0); 
        (A[14] *> O[23])=(0.0,0.0); 
        (A[14] *> O[24])=(0.0,0.0); 
        (A[14] *> O[25])=(0.0,0.0); 
        (A[14] *> O[26])=(0.0,0.0); 
        (A[14] *> O[27])=(0.0,0.0); 
        (A[14] *> O[28])=(0.0,0.0); 
        (A[14] *> O[29])=(0.0,0.0); 
        (A[14] *> O[30])=(0.0,0.0); 
        (A[14] *> O[31])=(0.0,0.0); 
        (A[15] *> O[0])=(0.0,0.0); 
        (A[15] *> O[1])=(0.0,0.0); 
        (A[15] *> O[2])=(0.0,0.0); 
        (A[15] *> O[3])=(0.0,0.0); 
        (A[15] *> O[4])=(0.0,0.0); 
        (A[15] *> O[5])=(0.0,0.0); 
        (A[15] *> O[6])=(0.0,0.0); 
        (A[15] *> O[7])=(0.0,0.0); 
        (A[15] *> O[8])=(0.0,0.0); 
        (A[15] *> O[9])=(0.0,0.0); 
        (A[15] *> O[10])=(0.0,0.0); 
        (A[15] *> O[11])=(0.0,0.0); 
        (A[15] *> O[12])=(0.0,0.0); 
        (A[15] *> O[13])=(0.0,0.0); 
        (A[15] *> O[14])=(0.0,0.0); 
        (A[15] *> O[15])=(0.0,0.0); 
        (A[15] *> O[16])=(0.0,0.0); 
        (A[15] *> O[17])=(0.0,0.0); 
        (A[15] *> O[18])=(0.0,0.0); 
        (A[15] *> O[19])=(0.0,0.0); 
        (A[15] *> O[20])=(0.0,0.0); 
        (A[15] *> O[21])=(0.0,0.0); 
        (A[15] *> O[22])=(0.0,0.0); 
        (A[15] *> O[23])=(0.0,0.0); 
        (A[15] *> O[24])=(0.0,0.0); 
        (A[15] *> O[25])=(0.0,0.0); 
        (A[15] *> O[26])=(0.0,0.0); 
        (A[15] *> O[27])=(0.0,0.0); 
        (A[15] *> O[28])=(0.0,0.0); 
        (A[15] *> O[29])=(0.0,0.0); 
        (A[15] *> O[30])=(0.0,0.0); 
        (A[15] *> O[31])=(0.0,0.0); 
        (B[0] *> O[0])=(0.0,0.0); 
        (B[0] *> O[1])=(0.0,0.0); 
        (B[0] *> O[2])=(0.0,0.0); 
        (B[0] *> O[3])=(0.0,0.0); 
        (B[0] *> O[4])=(0.0,0.0); 
        (B[0] *> O[5])=(0.0,0.0); 
        (B[0] *> O[6])=(0.0,0.0); 
        (B[0] *> O[7])=(0.0,0.0); 
        (B[0] *> O[8])=(0.0,0.0); 
        (B[0] *> O[9])=(0.0,0.0); 
        (B[0] *> O[10])=(0.0,0.0); 
        (B[0] *> O[11])=(0.0,0.0); 
        (B[0] *> O[12])=(0.0,0.0); 
        (B[0] *> O[13])=(0.0,0.0); 
        (B[0] *> O[14])=(0.0,0.0); 
        (B[0] *> O[15])=(0.0,0.0); 
        (B[0] *> O[16])=(0.0,0.0); 
        (B[0] *> O[17])=(0.0,0.0); 
        (B[0] *> O[18])=(0.0,0.0); 
        (B[0] *> O[19])=(0.0,0.0); 
        (B[0] *> O[20])=(0.0,0.0); 
        (B[0] *> O[21])=(0.0,0.0); 
        (B[0] *> O[22])=(0.0,0.0); 
        (B[0] *> O[23])=(0.0,0.0); 
        (B[0] *> O[24])=(0.0,0.0); 
        (B[0] *> O[25])=(0.0,0.0); 
        (B[0] *> O[26])=(0.0,0.0); 
        (B[0] *> O[27])=(0.0,0.0); 
        (B[0] *> O[28])=(0.0,0.0); 
        (B[0] *> O[29])=(0.0,0.0); 
        (B[0] *> O[30])=(0.0,0.0); 
        (B[0] *> O[31])=(0.0,0.0); 
        (B[1] *> O[0])=(0.0,0.0); 
        (B[1] *> O[1])=(0.0,0.0); 
        (B[1] *> O[2])=(0.0,0.0); 
        (B[1] *> O[3])=(0.0,0.0); 
        (B[1] *> O[4])=(0.0,0.0); 
        (B[1] *> O[5])=(0.0,0.0); 
        (B[1] *> O[6])=(0.0,0.0); 
        (B[1] *> O[7])=(0.0,0.0); 
        (B[1] *> O[8])=(0.0,0.0); 
        (B[1] *> O[9])=(0.0,0.0); 
        (B[1] *> O[10])=(0.0,0.0); 
        (B[1] *> O[11])=(0.0,0.0); 
        (B[1] *> O[12])=(0.0,0.0); 
        (B[1] *> O[13])=(0.0,0.0); 
        (B[1] *> O[14])=(0.0,0.0); 
        (B[1] *> O[15])=(0.0,0.0); 
        (B[1] *> O[16])=(0.0,0.0); 
        (B[1] *> O[17])=(0.0,0.0); 
        (B[1] *> O[18])=(0.0,0.0); 
        (B[1] *> O[19])=(0.0,0.0); 
        (B[1] *> O[20])=(0.0,0.0); 
        (B[1] *> O[21])=(0.0,0.0); 
        (B[1] *> O[22])=(0.0,0.0); 
        (B[1] *> O[23])=(0.0,0.0); 
        (B[1] *> O[24])=(0.0,0.0); 
        (B[1] *> O[25])=(0.0,0.0); 
        (B[1] *> O[26])=(0.0,0.0); 
        (B[1] *> O[27])=(0.0,0.0); 
        (B[1] *> O[28])=(0.0,0.0); 
        (B[1] *> O[29])=(0.0,0.0); 
        (B[1] *> O[30])=(0.0,0.0); 
        (B[1] *> O[31])=(0.0,0.0); 
        (B[2] *> O[0])=(0.0,0.0); 
        (B[2] *> O[1])=(0.0,0.0); 
        (B[2] *> O[2])=(0.0,0.0); 
        (B[2] *> O[3])=(0.0,0.0); 
        (B[2] *> O[4])=(0.0,0.0); 
        (B[2] *> O[5])=(0.0,0.0); 
        (B[2] *> O[6])=(0.0,0.0); 
        (B[2] *> O[7])=(0.0,0.0); 
        (B[2] *> O[8])=(0.0,0.0); 
        (B[2] *> O[9])=(0.0,0.0); 
        (B[2] *> O[10])=(0.0,0.0); 
        (B[2] *> O[11])=(0.0,0.0); 
        (B[2] *> O[12])=(0.0,0.0); 
        (B[2] *> O[13])=(0.0,0.0); 
        (B[2] *> O[14])=(0.0,0.0); 
        (B[2] *> O[15])=(0.0,0.0); 
        (B[2] *> O[16])=(0.0,0.0); 
        (B[2] *> O[17])=(0.0,0.0); 
        (B[2] *> O[18])=(0.0,0.0); 
        (B[2] *> O[19])=(0.0,0.0); 
        (B[2] *> O[20])=(0.0,0.0); 
        (B[2] *> O[21])=(0.0,0.0); 
        (B[2] *> O[22])=(0.0,0.0); 
        (B[2] *> O[23])=(0.0,0.0); 
        (B[2] *> O[24])=(0.0,0.0); 
        (B[2] *> O[25])=(0.0,0.0); 
        (B[2] *> O[26])=(0.0,0.0); 
        (B[2] *> O[27])=(0.0,0.0); 
        (B[2] *> O[28])=(0.0,0.0); 
        (B[2] *> O[29])=(0.0,0.0); 
        (B[2] *> O[30])=(0.0,0.0); 
        (B[2] *> O[31])=(0.0,0.0); 
        (B[3] *> O[0])=(0.0,0.0); 
        (B[3] *> O[1])=(0.0,0.0); 
        (B[3] *> O[2])=(0.0,0.0); 
        (B[3] *> O[3])=(0.0,0.0); 
        (B[3] *> O[4])=(0.0,0.0); 
        (B[3] *> O[5])=(0.0,0.0); 
        (B[3] *> O[6])=(0.0,0.0); 
        (B[3] *> O[7])=(0.0,0.0); 
        (B[3] *> O[8])=(0.0,0.0); 
        (B[3] *> O[9])=(0.0,0.0); 
        (B[3] *> O[10])=(0.0,0.0); 
        (B[3] *> O[11])=(0.0,0.0); 
        (B[3] *> O[12])=(0.0,0.0); 
        (B[3] *> O[13])=(0.0,0.0); 
        (B[3] *> O[14])=(0.0,0.0); 
        (B[3] *> O[15])=(0.0,0.0); 
        (B[3] *> O[16])=(0.0,0.0); 
        (B[3] *> O[17])=(0.0,0.0); 
        (B[3] *> O[18])=(0.0,0.0); 
        (B[3] *> O[19])=(0.0,0.0); 
        (B[3] *> O[20])=(0.0,0.0); 
        (B[3] *> O[21])=(0.0,0.0); 
        (B[3] *> O[22])=(0.0,0.0); 
        (B[3] *> O[23])=(0.0,0.0); 
        (B[3] *> O[24])=(0.0,0.0); 
        (B[3] *> O[25])=(0.0,0.0); 
        (B[3] *> O[26])=(0.0,0.0); 
        (B[3] *> O[27])=(0.0,0.0); 
        (B[3] *> O[28])=(0.0,0.0); 
        (B[3] *> O[29])=(0.0,0.0); 
        (B[3] *> O[30])=(0.0,0.0); 
        (B[3] *> O[31])=(0.0,0.0); 
        (B[4] *> O[0])=(0.0,0.0); 
        (B[4] *> O[1])=(0.0,0.0); 
        (B[4] *> O[2])=(0.0,0.0); 
        (B[4] *> O[3])=(0.0,0.0); 
        (B[4] *> O[4])=(0.0,0.0); 
        (B[4] *> O[5])=(0.0,0.0); 
        (B[4] *> O[6])=(0.0,0.0); 
        (B[4] *> O[7])=(0.0,0.0); 
        (B[4] *> O[8])=(0.0,0.0); 
        (B[4] *> O[9])=(0.0,0.0); 
        (B[4] *> O[10])=(0.0,0.0); 
        (B[4] *> O[11])=(0.0,0.0); 
        (B[4] *> O[12])=(0.0,0.0); 
        (B[4] *> O[13])=(0.0,0.0); 
        (B[4] *> O[14])=(0.0,0.0); 
        (B[4] *> O[15])=(0.0,0.0); 
        (B[4] *> O[16])=(0.0,0.0); 
        (B[4] *> O[17])=(0.0,0.0); 
        (B[4] *> O[18])=(0.0,0.0); 
        (B[4] *> O[19])=(0.0,0.0); 
        (B[4] *> O[20])=(0.0,0.0); 
        (B[4] *> O[21])=(0.0,0.0); 
        (B[4] *> O[22])=(0.0,0.0); 
        (B[4] *> O[23])=(0.0,0.0); 
        (B[4] *> O[24])=(0.0,0.0); 
        (B[4] *> O[25])=(0.0,0.0); 
        (B[4] *> O[26])=(0.0,0.0); 
        (B[4] *> O[27])=(0.0,0.0); 
        (B[4] *> O[28])=(0.0,0.0); 
        (B[4] *> O[29])=(0.0,0.0); 
        (B[4] *> O[30])=(0.0,0.0); 
        (B[4] *> O[31])=(0.0,0.0); 
        (B[5] *> O[0])=(0.0,0.0); 
        (B[5] *> O[1])=(0.0,0.0); 
        (B[5] *> O[2])=(0.0,0.0); 
        (B[5] *> O[3])=(0.0,0.0); 
        (B[5] *> O[4])=(0.0,0.0); 
        (B[5] *> O[5])=(0.0,0.0); 
        (B[5] *> O[6])=(0.0,0.0); 
        (B[5] *> O[7])=(0.0,0.0); 
        (B[5] *> O[8])=(0.0,0.0); 
        (B[5] *> O[9])=(0.0,0.0); 
        (B[5] *> O[10])=(0.0,0.0); 
        (B[5] *> O[11])=(0.0,0.0); 
        (B[5] *> O[12])=(0.0,0.0); 
        (B[5] *> O[13])=(0.0,0.0); 
        (B[5] *> O[14])=(0.0,0.0); 
        (B[5] *> O[15])=(0.0,0.0); 
        (B[5] *> O[16])=(0.0,0.0); 
        (B[5] *> O[17])=(0.0,0.0); 
        (B[5] *> O[18])=(0.0,0.0); 
        (B[5] *> O[19])=(0.0,0.0); 
        (B[5] *> O[20])=(0.0,0.0); 
        (B[5] *> O[21])=(0.0,0.0); 
        (B[5] *> O[22])=(0.0,0.0); 
        (B[5] *> O[23])=(0.0,0.0); 
        (B[5] *> O[24])=(0.0,0.0); 
        (B[5] *> O[25])=(0.0,0.0); 
        (B[5] *> O[26])=(0.0,0.0); 
        (B[5] *> O[27])=(0.0,0.0); 
        (B[5] *> O[28])=(0.0,0.0); 
        (B[5] *> O[29])=(0.0,0.0); 
        (B[5] *> O[30])=(0.0,0.0); 
        (B[5] *> O[31])=(0.0,0.0); 
        (B[6] *> O[0])=(0.0,0.0); 
        (B[6] *> O[1])=(0.0,0.0); 
        (B[6] *> O[2])=(0.0,0.0); 
        (B[6] *> O[3])=(0.0,0.0); 
        (B[6] *> O[4])=(0.0,0.0); 
        (B[6] *> O[5])=(0.0,0.0); 
        (B[6] *> O[6])=(0.0,0.0); 
        (B[6] *> O[7])=(0.0,0.0); 
        (B[6] *> O[8])=(0.0,0.0); 
        (B[6] *> O[9])=(0.0,0.0); 
        (B[6] *> O[10])=(0.0,0.0); 
        (B[6] *> O[11])=(0.0,0.0); 
        (B[6] *> O[12])=(0.0,0.0); 
        (B[6] *> O[13])=(0.0,0.0); 
        (B[6] *> O[14])=(0.0,0.0); 
        (B[6] *> O[15])=(0.0,0.0); 
        (B[6] *> O[16])=(0.0,0.0); 
        (B[6] *> O[17])=(0.0,0.0); 
        (B[6] *> O[18])=(0.0,0.0); 
        (B[6] *> O[19])=(0.0,0.0); 
        (B[6] *> O[20])=(0.0,0.0); 
        (B[6] *> O[21])=(0.0,0.0); 
        (B[6] *> O[22])=(0.0,0.0); 
        (B[6] *> O[23])=(0.0,0.0); 
        (B[6] *> O[24])=(0.0,0.0); 
        (B[6] *> O[25])=(0.0,0.0); 
        (B[6] *> O[26])=(0.0,0.0); 
        (B[6] *> O[27])=(0.0,0.0); 
        (B[6] *> O[28])=(0.0,0.0); 
        (B[6] *> O[29])=(0.0,0.0); 
        (B[6] *> O[30])=(0.0,0.0); 
        (B[6] *> O[31])=(0.0,0.0); 
        (B[7] *> O[0])=(0.0,0.0); 
        (B[7] *> O[1])=(0.0,0.0); 
        (B[7] *> O[2])=(0.0,0.0); 
        (B[7] *> O[3])=(0.0,0.0); 
        (B[7] *> O[4])=(0.0,0.0); 
        (B[7] *> O[5])=(0.0,0.0); 
        (B[7] *> O[6])=(0.0,0.0); 
        (B[7] *> O[7])=(0.0,0.0); 
        (B[7] *> O[8])=(0.0,0.0); 
        (B[7] *> O[9])=(0.0,0.0); 
        (B[7] *> O[10])=(0.0,0.0); 
        (B[7] *> O[11])=(0.0,0.0); 
        (B[7] *> O[12])=(0.0,0.0); 
        (B[7] *> O[13])=(0.0,0.0); 
        (B[7] *> O[14])=(0.0,0.0); 
        (B[7] *> O[15])=(0.0,0.0); 
        (B[7] *> O[16])=(0.0,0.0); 
        (B[7] *> O[17])=(0.0,0.0); 
        (B[7] *> O[18])=(0.0,0.0); 
        (B[7] *> O[19])=(0.0,0.0); 
        (B[7] *> O[20])=(0.0,0.0); 
        (B[7] *> O[21])=(0.0,0.0); 
        (B[7] *> O[22])=(0.0,0.0); 
        (B[7] *> O[23])=(0.0,0.0); 
        (B[7] *> O[24])=(0.0,0.0); 
        (B[7] *> O[25])=(0.0,0.0); 
        (B[7] *> O[26])=(0.0,0.0); 
        (B[7] *> O[27])=(0.0,0.0); 
        (B[7] *> O[28])=(0.0,0.0); 
        (B[7] *> O[29])=(0.0,0.0); 
        (B[7] *> O[30])=(0.0,0.0); 
        (B[7] *> O[31])=(0.0,0.0); 
        (B[8] *> O[0])=(0.0,0.0); 
        (B[8] *> O[1])=(0.0,0.0); 
        (B[8] *> O[2])=(0.0,0.0); 
        (B[8] *> O[3])=(0.0,0.0); 
        (B[8] *> O[4])=(0.0,0.0); 
        (B[8] *> O[5])=(0.0,0.0); 
        (B[8] *> O[6])=(0.0,0.0); 
        (B[8] *> O[7])=(0.0,0.0); 
        (B[8] *> O[8])=(0.0,0.0); 
        (B[8] *> O[9])=(0.0,0.0); 
        (B[8] *> O[10])=(0.0,0.0); 
        (B[8] *> O[11])=(0.0,0.0); 
        (B[8] *> O[12])=(0.0,0.0); 
        (B[8] *> O[13])=(0.0,0.0); 
        (B[8] *> O[14])=(0.0,0.0); 
        (B[8] *> O[15])=(0.0,0.0); 
        (B[8] *> O[16])=(0.0,0.0); 
        (B[8] *> O[17])=(0.0,0.0); 
        (B[8] *> O[18])=(0.0,0.0); 
        (B[8] *> O[19])=(0.0,0.0); 
        (B[8] *> O[20])=(0.0,0.0); 
        (B[8] *> O[21])=(0.0,0.0); 
        (B[8] *> O[22])=(0.0,0.0); 
        (B[8] *> O[23])=(0.0,0.0); 
        (B[8] *> O[24])=(0.0,0.0); 
        (B[8] *> O[25])=(0.0,0.0); 
        (B[8] *> O[26])=(0.0,0.0); 
        (B[8] *> O[27])=(0.0,0.0); 
        (B[8] *> O[28])=(0.0,0.0); 
        (B[8] *> O[29])=(0.0,0.0); 
        (B[8] *> O[30])=(0.0,0.0); 
        (B[8] *> O[31])=(0.0,0.0); 
        (B[9] *> O[0])=(0.0,0.0); 
        (B[9] *> O[1])=(0.0,0.0); 
        (B[9] *> O[2])=(0.0,0.0); 
        (B[9] *> O[3])=(0.0,0.0); 
        (B[9] *> O[4])=(0.0,0.0); 
        (B[9] *> O[5])=(0.0,0.0); 
        (B[9] *> O[6])=(0.0,0.0); 
        (B[9] *> O[7])=(0.0,0.0); 
        (B[9] *> O[8])=(0.0,0.0); 
        (B[9] *> O[9])=(0.0,0.0); 
        (B[9] *> O[10])=(0.0,0.0); 
        (B[9] *> O[11])=(0.0,0.0); 
        (B[9] *> O[12])=(0.0,0.0); 
        (B[9] *> O[13])=(0.0,0.0); 
        (B[9] *> O[14])=(0.0,0.0); 
        (B[9] *> O[15])=(0.0,0.0); 
        (B[9] *> O[16])=(0.0,0.0); 
        (B[9] *> O[17])=(0.0,0.0); 
        (B[9] *> O[18])=(0.0,0.0); 
        (B[9] *> O[19])=(0.0,0.0); 
        (B[9] *> O[20])=(0.0,0.0); 
        (B[9] *> O[21])=(0.0,0.0); 
        (B[9] *> O[22])=(0.0,0.0); 
        (B[9] *> O[23])=(0.0,0.0); 
        (B[9] *> O[24])=(0.0,0.0); 
        (B[9] *> O[25])=(0.0,0.0); 
        (B[9] *> O[26])=(0.0,0.0); 
        (B[9] *> O[27])=(0.0,0.0); 
        (B[9] *> O[28])=(0.0,0.0); 
        (B[9] *> O[29])=(0.0,0.0); 
        (B[9] *> O[30])=(0.0,0.0); 
        (B[9] *> O[31])=(0.0,0.0); 
        (B[10] *> O[0])=(0.0,0.0); 
        (B[10] *> O[1])=(0.0,0.0); 
        (B[10] *> O[2])=(0.0,0.0); 
        (B[10] *> O[3])=(0.0,0.0); 
        (B[10] *> O[4])=(0.0,0.0); 
        (B[10] *> O[5])=(0.0,0.0); 
        (B[10] *> O[6])=(0.0,0.0); 
        (B[10] *> O[7])=(0.0,0.0); 
        (B[10] *> O[8])=(0.0,0.0); 
        (B[10] *> O[9])=(0.0,0.0); 
        (B[10] *> O[10])=(0.0,0.0); 
        (B[10] *> O[11])=(0.0,0.0); 
        (B[10] *> O[12])=(0.0,0.0); 
        (B[10] *> O[13])=(0.0,0.0); 
        (B[10] *> O[14])=(0.0,0.0); 
        (B[10] *> O[15])=(0.0,0.0); 
        (B[10] *> O[16])=(0.0,0.0); 
        (B[10] *> O[17])=(0.0,0.0); 
        (B[10] *> O[18])=(0.0,0.0); 
        (B[10] *> O[19])=(0.0,0.0); 
        (B[10] *> O[20])=(0.0,0.0); 
        (B[10] *> O[21])=(0.0,0.0); 
        (B[10] *> O[22])=(0.0,0.0); 
        (B[10] *> O[23])=(0.0,0.0); 
        (B[10] *> O[24])=(0.0,0.0); 
        (B[10] *> O[25])=(0.0,0.0); 
        (B[10] *> O[26])=(0.0,0.0); 
        (B[10] *> O[27])=(0.0,0.0); 
        (B[10] *> O[28])=(0.0,0.0); 
        (B[10] *> O[29])=(0.0,0.0); 
        (B[10] *> O[30])=(0.0,0.0); 
        (B[10] *> O[31])=(0.0,0.0); 
        (B[11] *> O[0])=(0.0,0.0); 
        (B[11] *> O[1])=(0.0,0.0); 
        (B[11] *> O[2])=(0.0,0.0); 
        (B[11] *> O[3])=(0.0,0.0); 
        (B[11] *> O[4])=(0.0,0.0); 
        (B[11] *> O[5])=(0.0,0.0); 
        (B[11] *> O[6])=(0.0,0.0); 
        (B[11] *> O[7])=(0.0,0.0); 
        (B[11] *> O[8])=(0.0,0.0); 
        (B[11] *> O[9])=(0.0,0.0); 
        (B[11] *> O[10])=(0.0,0.0); 
        (B[11] *> O[11])=(0.0,0.0); 
        (B[11] *> O[12])=(0.0,0.0); 
        (B[11] *> O[13])=(0.0,0.0); 
        (B[11] *> O[14])=(0.0,0.0); 
        (B[11] *> O[15])=(0.0,0.0); 
        (B[11] *> O[16])=(0.0,0.0); 
        (B[11] *> O[17])=(0.0,0.0); 
        (B[11] *> O[18])=(0.0,0.0); 
        (B[11] *> O[19])=(0.0,0.0); 
        (B[11] *> O[20])=(0.0,0.0); 
        (B[11] *> O[21])=(0.0,0.0); 
        (B[11] *> O[22])=(0.0,0.0); 
        (B[11] *> O[23])=(0.0,0.0); 
        (B[11] *> O[24])=(0.0,0.0); 
        (B[11] *> O[25])=(0.0,0.0); 
        (B[11] *> O[26])=(0.0,0.0); 
        (B[11] *> O[27])=(0.0,0.0); 
        (B[11] *> O[28])=(0.0,0.0); 
        (B[11] *> O[29])=(0.0,0.0); 
        (B[11] *> O[30])=(0.0,0.0); 
        (B[11] *> O[31])=(0.0,0.0); 
        (B[12] *> O[0])=(0.0,0.0); 
        (B[12] *> O[1])=(0.0,0.0); 
        (B[12] *> O[2])=(0.0,0.0); 
        (B[12] *> O[3])=(0.0,0.0); 
        (B[12] *> O[4])=(0.0,0.0); 
        (B[12] *> O[5])=(0.0,0.0); 
        (B[12] *> O[6])=(0.0,0.0); 
        (B[12] *> O[7])=(0.0,0.0); 
        (B[12] *> O[8])=(0.0,0.0); 
        (B[12] *> O[9])=(0.0,0.0); 
        (B[12] *> O[10])=(0.0,0.0); 
        (B[12] *> O[11])=(0.0,0.0); 
        (B[12] *> O[12])=(0.0,0.0); 
        (B[12] *> O[13])=(0.0,0.0); 
        (B[12] *> O[14])=(0.0,0.0); 
        (B[12] *> O[15])=(0.0,0.0); 
        (B[12] *> O[16])=(0.0,0.0); 
        (B[12] *> O[17])=(0.0,0.0); 
        (B[12] *> O[18])=(0.0,0.0); 
        (B[12] *> O[19])=(0.0,0.0); 
        (B[12] *> O[20])=(0.0,0.0); 
        (B[12] *> O[21])=(0.0,0.0); 
        (B[12] *> O[22])=(0.0,0.0); 
        (B[12] *> O[23])=(0.0,0.0); 
        (B[12] *> O[24])=(0.0,0.0); 
        (B[12] *> O[25])=(0.0,0.0); 
        (B[12] *> O[26])=(0.0,0.0); 
        (B[12] *> O[27])=(0.0,0.0); 
        (B[12] *> O[28])=(0.0,0.0); 
        (B[12] *> O[29])=(0.0,0.0); 
        (B[12] *> O[30])=(0.0,0.0); 
        (B[12] *> O[31])=(0.0,0.0); 
        (B[13] *> O[0])=(0.0,0.0); 
        (B[13] *> O[1])=(0.0,0.0); 
        (B[13] *> O[2])=(0.0,0.0); 
        (B[13] *> O[3])=(0.0,0.0); 
        (B[13] *> O[4])=(0.0,0.0); 
        (B[13] *> O[5])=(0.0,0.0); 
        (B[13] *> O[6])=(0.0,0.0); 
        (B[13] *> O[7])=(0.0,0.0); 
        (B[13] *> O[8])=(0.0,0.0); 
        (B[13] *> O[9])=(0.0,0.0); 
        (B[13] *> O[10])=(0.0,0.0); 
        (B[13] *> O[11])=(0.0,0.0); 
        (B[13] *> O[12])=(0.0,0.0); 
        (B[13] *> O[13])=(0.0,0.0); 
        (B[13] *> O[14])=(0.0,0.0); 
        (B[13] *> O[15])=(0.0,0.0); 
        (B[13] *> O[16])=(0.0,0.0); 
        (B[13] *> O[17])=(0.0,0.0); 
        (B[13] *> O[18])=(0.0,0.0); 
        (B[13] *> O[19])=(0.0,0.0); 
        (B[13] *> O[20])=(0.0,0.0); 
        (B[13] *> O[21])=(0.0,0.0); 
        (B[13] *> O[22])=(0.0,0.0); 
        (B[13] *> O[23])=(0.0,0.0); 
        (B[13] *> O[24])=(0.0,0.0); 
        (B[13] *> O[25])=(0.0,0.0); 
        (B[13] *> O[26])=(0.0,0.0); 
        (B[13] *> O[27])=(0.0,0.0); 
        (B[13] *> O[28])=(0.0,0.0); 
        (B[13] *> O[29])=(0.0,0.0); 
        (B[13] *> O[30])=(0.0,0.0); 
        (B[13] *> O[31])=(0.0,0.0); 
        (B[14] *> O[0])=(0.0,0.0); 
        (B[14] *> O[1])=(0.0,0.0); 
        (B[14] *> O[2])=(0.0,0.0); 
        (B[14] *> O[3])=(0.0,0.0); 
        (B[14] *> O[4])=(0.0,0.0); 
        (B[14] *> O[5])=(0.0,0.0); 
        (B[14] *> O[6])=(0.0,0.0); 
        (B[14] *> O[7])=(0.0,0.0); 
        (B[14] *> O[8])=(0.0,0.0); 
        (B[14] *> O[9])=(0.0,0.0); 
        (B[14] *> O[10])=(0.0,0.0); 
        (B[14] *> O[11])=(0.0,0.0); 
        (B[14] *> O[12])=(0.0,0.0); 
        (B[14] *> O[13])=(0.0,0.0); 
        (B[14] *> O[14])=(0.0,0.0); 
        (B[14] *> O[15])=(0.0,0.0); 
        (B[14] *> O[16])=(0.0,0.0); 
        (B[14] *> O[17])=(0.0,0.0); 
        (B[14] *> O[18])=(0.0,0.0); 
        (B[14] *> O[19])=(0.0,0.0); 
        (B[14] *> O[20])=(0.0,0.0); 
        (B[14] *> O[21])=(0.0,0.0); 
        (B[14] *> O[22])=(0.0,0.0); 
        (B[14] *> O[23])=(0.0,0.0); 
        (B[14] *> O[24])=(0.0,0.0); 
        (B[14] *> O[25])=(0.0,0.0); 
        (B[14] *> O[26])=(0.0,0.0); 
        (B[14] *> O[27])=(0.0,0.0); 
        (B[14] *> O[28])=(0.0,0.0); 
        (B[14] *> O[29])=(0.0,0.0); 
        (B[14] *> O[30])=(0.0,0.0); 
        (B[14] *> O[31])=(0.0,0.0); 
        (B[15] *> O[0])=(0.0,0.0); 
        (B[15] *> O[1])=(0.0,0.0); 
        (B[15] *> O[2])=(0.0,0.0); 
        (B[15] *> O[3])=(0.0,0.0); 
        (B[15] *> O[4])=(0.0,0.0); 
        (B[15] *> O[5])=(0.0,0.0); 
        (B[15] *> O[6])=(0.0,0.0); 
        (B[15] *> O[7])=(0.0,0.0); 
        (B[15] *> O[8])=(0.0,0.0); 
        (B[15] *> O[9])=(0.0,0.0); 
        (B[15] *> O[10])=(0.0,0.0); 
        (B[15] *> O[11])=(0.0,0.0); 
        (B[15] *> O[12])=(0.0,0.0); 
        (B[15] *> O[13])=(0.0,0.0); 
        (B[15] *> O[14])=(0.0,0.0); 
        (B[15] *> O[15])=(0.0,0.0); 
        (B[15] *> O[16])=(0.0,0.0); 
        (B[15] *> O[17])=(0.0,0.0); 
        (B[15] *> O[18])=(0.0,0.0); 
        (B[15] *> O[19])=(0.0,0.0); 
        (B[15] *> O[20])=(0.0,0.0); 
        (B[15] *> O[21])=(0.0,0.0); 
        (B[15] *> O[22])=(0.0,0.0); 
        (B[15] *> O[23])=(0.0,0.0); 
        (B[15] *> O[24])=(0.0,0.0); 
        (B[15] *> O[25])=(0.0,0.0); 
        (B[15] *> O[26])=(0.0,0.0); 
        (B[15] *> O[27])=(0.0,0.0); 
        (B[15] *> O[28])=(0.0,0.0); 
        (B[15] *> O[29])=(0.0,0.0); 
        (B[15] *> O[30])=(0.0,0.0); 
        (B[15] *> O[31])=(0.0,0.0); 
        (C[0] *> O[0])=(0.0,0.0); 
        (C[0] *> O[1])=(0.0,0.0); 
        (C[0] *> O[2])=(0.0,0.0); 
        (C[0] *> O[3])=(0.0,0.0); 
        (C[0] *> O[4])=(0.0,0.0); 
        (C[0] *> O[5])=(0.0,0.0); 
        (C[0] *> O[6])=(0.0,0.0); 
        (C[0] *> O[7])=(0.0,0.0); 
        (C[0] *> O[8])=(0.0,0.0); 
        (C[0] *> O[9])=(0.0,0.0); 
        (C[0] *> O[10])=(0.0,0.0); 
        (C[0] *> O[11])=(0.0,0.0); 
        (C[0] *> O[12])=(0.0,0.0); 
        (C[0] *> O[13])=(0.0,0.0); 
        (C[0] *> O[14])=(0.0,0.0); 
        (C[0] *> O[15])=(0.0,0.0); 
        (C[0] *> O[16])=(0.0,0.0); 
        (C[0] *> O[17])=(0.0,0.0); 
        (C[0] *> O[18])=(0.0,0.0); 
        (C[0] *> O[19])=(0.0,0.0); 
        (C[0] *> O[20])=(0.0,0.0); 
        (C[0] *> O[21])=(0.0,0.0); 
        (C[0] *> O[22])=(0.0,0.0); 
        (C[0] *> O[23])=(0.0,0.0); 
        (C[0] *> O[24])=(0.0,0.0); 
        (C[0] *> O[25])=(0.0,0.0); 
        (C[0] *> O[26])=(0.0,0.0); 
        (C[0] *> O[27])=(0.0,0.0); 
        (C[0] *> O[28])=(0.0,0.0); 
        (C[0] *> O[29])=(0.0,0.0); 
        (C[0] *> O[30])=(0.0,0.0); 
        (C[0] *> O[31])=(0.0,0.0); 
        (C[1] *> O[0])=(0.0,0.0); 
        (C[1] *> O[1])=(0.0,0.0); 
        (C[1] *> O[2])=(0.0,0.0); 
        (C[1] *> O[3])=(0.0,0.0); 
        (C[1] *> O[4])=(0.0,0.0); 
        (C[1] *> O[5])=(0.0,0.0); 
        (C[1] *> O[6])=(0.0,0.0); 
        (C[1] *> O[7])=(0.0,0.0); 
        (C[1] *> O[8])=(0.0,0.0); 
        (C[1] *> O[9])=(0.0,0.0); 
        (C[1] *> O[10])=(0.0,0.0); 
        (C[1] *> O[11])=(0.0,0.0); 
        (C[1] *> O[12])=(0.0,0.0); 
        (C[1] *> O[13])=(0.0,0.0); 
        (C[1] *> O[14])=(0.0,0.0); 
        (C[1] *> O[15])=(0.0,0.0); 
        (C[1] *> O[16])=(0.0,0.0); 
        (C[1] *> O[17])=(0.0,0.0); 
        (C[1] *> O[18])=(0.0,0.0); 
        (C[1] *> O[19])=(0.0,0.0); 
        (C[1] *> O[20])=(0.0,0.0); 
        (C[1] *> O[21])=(0.0,0.0); 
        (C[1] *> O[22])=(0.0,0.0); 
        (C[1] *> O[23])=(0.0,0.0); 
        (C[1] *> O[24])=(0.0,0.0); 
        (C[1] *> O[25])=(0.0,0.0); 
        (C[1] *> O[26])=(0.0,0.0); 
        (C[1] *> O[27])=(0.0,0.0); 
        (C[1] *> O[28])=(0.0,0.0); 
        (C[1] *> O[29])=(0.0,0.0); 
        (C[1] *> O[30])=(0.0,0.0); 
        (C[1] *> O[31])=(0.0,0.0); 
        (C[2] *> O[0])=(0.0,0.0); 
        (C[2] *> O[1])=(0.0,0.0); 
        (C[2] *> O[2])=(0.0,0.0); 
        (C[2] *> O[3])=(0.0,0.0); 
        (C[2] *> O[4])=(0.0,0.0); 
        (C[2] *> O[5])=(0.0,0.0); 
        (C[2] *> O[6])=(0.0,0.0); 
        (C[2] *> O[7])=(0.0,0.0); 
        (C[2] *> O[8])=(0.0,0.0); 
        (C[2] *> O[9])=(0.0,0.0); 
        (C[2] *> O[10])=(0.0,0.0); 
        (C[2] *> O[11])=(0.0,0.0); 
        (C[2] *> O[12])=(0.0,0.0); 
        (C[2] *> O[13])=(0.0,0.0); 
        (C[2] *> O[14])=(0.0,0.0); 
        (C[2] *> O[15])=(0.0,0.0); 
        (C[2] *> O[16])=(0.0,0.0); 
        (C[2] *> O[17])=(0.0,0.0); 
        (C[2] *> O[18])=(0.0,0.0); 
        (C[2] *> O[19])=(0.0,0.0); 
        (C[2] *> O[20])=(0.0,0.0); 
        (C[2] *> O[21])=(0.0,0.0); 
        (C[2] *> O[22])=(0.0,0.0); 
        (C[2] *> O[23])=(0.0,0.0); 
        (C[2] *> O[24])=(0.0,0.0); 
        (C[2] *> O[25])=(0.0,0.0); 
        (C[2] *> O[26])=(0.0,0.0); 
        (C[2] *> O[27])=(0.0,0.0); 
        (C[2] *> O[28])=(0.0,0.0); 
        (C[2] *> O[29])=(0.0,0.0); 
        (C[2] *> O[30])=(0.0,0.0); 
        (C[2] *> O[31])=(0.0,0.0); 
        (C[3] *> O[0])=(0.0,0.0); 
        (C[3] *> O[1])=(0.0,0.0); 
        (C[3] *> O[2])=(0.0,0.0); 
        (C[3] *> O[3])=(0.0,0.0); 
        (C[3] *> O[4])=(0.0,0.0); 
        (C[3] *> O[5])=(0.0,0.0); 
        (C[3] *> O[6])=(0.0,0.0); 
        (C[3] *> O[7])=(0.0,0.0); 
        (C[3] *> O[8])=(0.0,0.0); 
        (C[3] *> O[9])=(0.0,0.0); 
        (C[3] *> O[10])=(0.0,0.0); 
        (C[3] *> O[11])=(0.0,0.0); 
        (C[3] *> O[12])=(0.0,0.0); 
        (C[3] *> O[13])=(0.0,0.0); 
        (C[3] *> O[14])=(0.0,0.0); 
        (C[3] *> O[15])=(0.0,0.0); 
        (C[3] *> O[16])=(0.0,0.0); 
        (C[3] *> O[17])=(0.0,0.0); 
        (C[3] *> O[18])=(0.0,0.0); 
        (C[3] *> O[19])=(0.0,0.0); 
        (C[3] *> O[20])=(0.0,0.0); 
        (C[3] *> O[21])=(0.0,0.0); 
        (C[3] *> O[22])=(0.0,0.0); 
        (C[3] *> O[23])=(0.0,0.0); 
        (C[3] *> O[24])=(0.0,0.0); 
        (C[3] *> O[25])=(0.0,0.0); 
        (C[3] *> O[26])=(0.0,0.0); 
        (C[3] *> O[27])=(0.0,0.0); 
        (C[3] *> O[28])=(0.0,0.0); 
        (C[3] *> O[29])=(0.0,0.0); 
        (C[3] *> O[30])=(0.0,0.0); 
        (C[3] *> O[31])=(0.0,0.0); 
        (C[4] *> O[0])=(0.0,0.0); 
        (C[4] *> O[1])=(0.0,0.0); 
        (C[4] *> O[2])=(0.0,0.0); 
        (C[4] *> O[3])=(0.0,0.0); 
        (C[4] *> O[4])=(0.0,0.0); 
        (C[4] *> O[5])=(0.0,0.0); 
        (C[4] *> O[6])=(0.0,0.0); 
        (C[4] *> O[7])=(0.0,0.0); 
        (C[4] *> O[8])=(0.0,0.0); 
        (C[4] *> O[9])=(0.0,0.0); 
        (C[4] *> O[10])=(0.0,0.0); 
        (C[4] *> O[11])=(0.0,0.0); 
        (C[4] *> O[12])=(0.0,0.0); 
        (C[4] *> O[13])=(0.0,0.0); 
        (C[4] *> O[14])=(0.0,0.0); 
        (C[4] *> O[15])=(0.0,0.0); 
        (C[4] *> O[16])=(0.0,0.0); 
        (C[4] *> O[17])=(0.0,0.0); 
        (C[4] *> O[18])=(0.0,0.0); 
        (C[4] *> O[19])=(0.0,0.0); 
        (C[4] *> O[20])=(0.0,0.0); 
        (C[4] *> O[21])=(0.0,0.0); 
        (C[4] *> O[22])=(0.0,0.0); 
        (C[4] *> O[23])=(0.0,0.0); 
        (C[4] *> O[24])=(0.0,0.0); 
        (C[4] *> O[25])=(0.0,0.0); 
        (C[4] *> O[26])=(0.0,0.0); 
        (C[4] *> O[27])=(0.0,0.0); 
        (C[4] *> O[28])=(0.0,0.0); 
        (C[4] *> O[29])=(0.0,0.0); 
        (C[4] *> O[30])=(0.0,0.0); 
        (C[4] *> O[31])=(0.0,0.0); 
        (C[5] *> O[0])=(0.0,0.0); 
        (C[5] *> O[1])=(0.0,0.0); 
        (C[5] *> O[2])=(0.0,0.0); 
        (C[5] *> O[3])=(0.0,0.0); 
        (C[5] *> O[4])=(0.0,0.0); 
        (C[5] *> O[5])=(0.0,0.0); 
        (C[5] *> O[6])=(0.0,0.0); 
        (C[5] *> O[7])=(0.0,0.0); 
        (C[5] *> O[8])=(0.0,0.0); 
        (C[5] *> O[9])=(0.0,0.0); 
        (C[5] *> O[10])=(0.0,0.0); 
        (C[5] *> O[11])=(0.0,0.0); 
        (C[5] *> O[12])=(0.0,0.0); 
        (C[5] *> O[13])=(0.0,0.0); 
        (C[5] *> O[14])=(0.0,0.0); 
        (C[5] *> O[15])=(0.0,0.0); 
        (C[5] *> O[16])=(0.0,0.0); 
        (C[5] *> O[17])=(0.0,0.0); 
        (C[5] *> O[18])=(0.0,0.0); 
        (C[5] *> O[19])=(0.0,0.0); 
        (C[5] *> O[20])=(0.0,0.0); 
        (C[5] *> O[21])=(0.0,0.0); 
        (C[5] *> O[22])=(0.0,0.0); 
        (C[5] *> O[23])=(0.0,0.0); 
        (C[5] *> O[24])=(0.0,0.0); 
        (C[5] *> O[25])=(0.0,0.0); 
        (C[5] *> O[26])=(0.0,0.0); 
        (C[5] *> O[27])=(0.0,0.0); 
        (C[5] *> O[28])=(0.0,0.0); 
        (C[5] *> O[29])=(0.0,0.0); 
        (C[5] *> O[30])=(0.0,0.0); 
        (C[5] *> O[31])=(0.0,0.0); 
        (C[6] *> O[0])=(0.0,0.0); 
        (C[6] *> O[1])=(0.0,0.0); 
        (C[6] *> O[2])=(0.0,0.0); 
        (C[6] *> O[3])=(0.0,0.0); 
        (C[6] *> O[4])=(0.0,0.0); 
        (C[6] *> O[5])=(0.0,0.0); 
        (C[6] *> O[6])=(0.0,0.0); 
        (C[6] *> O[7])=(0.0,0.0); 
        (C[6] *> O[8])=(0.0,0.0); 
        (C[6] *> O[9])=(0.0,0.0); 
        (C[6] *> O[10])=(0.0,0.0); 
        (C[6] *> O[11])=(0.0,0.0); 
        (C[6] *> O[12])=(0.0,0.0); 
        (C[6] *> O[13])=(0.0,0.0); 
        (C[6] *> O[14])=(0.0,0.0); 
        (C[6] *> O[15])=(0.0,0.0); 
        (C[6] *> O[16])=(0.0,0.0); 
        (C[6] *> O[17])=(0.0,0.0); 
        (C[6] *> O[18])=(0.0,0.0); 
        (C[6] *> O[19])=(0.0,0.0); 
        (C[6] *> O[20])=(0.0,0.0); 
        (C[6] *> O[21])=(0.0,0.0); 
        (C[6] *> O[22])=(0.0,0.0); 
        (C[6] *> O[23])=(0.0,0.0); 
        (C[6] *> O[24])=(0.0,0.0); 
        (C[6] *> O[25])=(0.0,0.0); 
        (C[6] *> O[26])=(0.0,0.0); 
        (C[6] *> O[27])=(0.0,0.0); 
        (C[6] *> O[28])=(0.0,0.0); 
        (C[6] *> O[29])=(0.0,0.0); 
        (C[6] *> O[30])=(0.0,0.0); 
        (C[6] *> O[31])=(0.0,0.0); 
        (C[7] *> O[0])=(0.0,0.0); 
        (C[7] *> O[1])=(0.0,0.0); 
        (C[7] *> O[2])=(0.0,0.0); 
        (C[7] *> O[3])=(0.0,0.0); 
        (C[7] *> O[4])=(0.0,0.0); 
        (C[7] *> O[5])=(0.0,0.0); 
        (C[7] *> O[6])=(0.0,0.0); 
        (C[7] *> O[7])=(0.0,0.0); 
        (C[7] *> O[8])=(0.0,0.0); 
        (C[7] *> O[9])=(0.0,0.0); 
        (C[7] *> O[10])=(0.0,0.0); 
        (C[7] *> O[11])=(0.0,0.0); 
        (C[7] *> O[12])=(0.0,0.0); 
        (C[7] *> O[13])=(0.0,0.0); 
        (C[7] *> O[14])=(0.0,0.0); 
        (C[7] *> O[15])=(0.0,0.0); 
        (C[7] *> O[16])=(0.0,0.0); 
        (C[7] *> O[17])=(0.0,0.0); 
        (C[7] *> O[18])=(0.0,0.0); 
        (C[7] *> O[19])=(0.0,0.0); 
        (C[7] *> O[20])=(0.0,0.0); 
        (C[7] *> O[21])=(0.0,0.0); 
        (C[7] *> O[22])=(0.0,0.0); 
        (C[7] *> O[23])=(0.0,0.0); 
        (C[7] *> O[24])=(0.0,0.0); 
        (C[7] *> O[25])=(0.0,0.0); 
        (C[7] *> O[26])=(0.0,0.0); 
        (C[7] *> O[27])=(0.0,0.0); 
        (C[7] *> O[28])=(0.0,0.0); 
        (C[7] *> O[29])=(0.0,0.0); 
        (C[7] *> O[30])=(0.0,0.0); 
        (C[7] *> O[31])=(0.0,0.0); 
        (C[8] *> O[0])=(0.0,0.0); 
        (C[8] *> O[1])=(0.0,0.0); 
        (C[8] *> O[2])=(0.0,0.0); 
        (C[8] *> O[3])=(0.0,0.0); 
        (C[8] *> O[4])=(0.0,0.0); 
        (C[8] *> O[5])=(0.0,0.0); 
        (C[8] *> O[6])=(0.0,0.0); 
        (C[8] *> O[7])=(0.0,0.0); 
        (C[8] *> O[8])=(0.0,0.0); 
        (C[8] *> O[9])=(0.0,0.0); 
        (C[8] *> O[10])=(0.0,0.0); 
        (C[8] *> O[11])=(0.0,0.0); 
        (C[8] *> O[12])=(0.0,0.0); 
        (C[8] *> O[13])=(0.0,0.0); 
        (C[8] *> O[14])=(0.0,0.0); 
        (C[8] *> O[15])=(0.0,0.0); 
        (C[8] *> O[16])=(0.0,0.0); 
        (C[8] *> O[17])=(0.0,0.0); 
        (C[8] *> O[18])=(0.0,0.0); 
        (C[8] *> O[19])=(0.0,0.0); 
        (C[8] *> O[20])=(0.0,0.0); 
        (C[8] *> O[21])=(0.0,0.0); 
        (C[8] *> O[22])=(0.0,0.0); 
        (C[8] *> O[23])=(0.0,0.0); 
        (C[8] *> O[24])=(0.0,0.0); 
        (C[8] *> O[25])=(0.0,0.0); 
        (C[8] *> O[26])=(0.0,0.0); 
        (C[8] *> O[27])=(0.0,0.0); 
        (C[8] *> O[28])=(0.0,0.0); 
        (C[8] *> O[29])=(0.0,0.0); 
        (C[8] *> O[30])=(0.0,0.0); 
        (C[8] *> O[31])=(0.0,0.0); 
        (C[9] *> O[0])=(0.0,0.0); 
        (C[9] *> O[1])=(0.0,0.0); 
        (C[9] *> O[2])=(0.0,0.0); 
        (C[9] *> O[3])=(0.0,0.0); 
        (C[9] *> O[4])=(0.0,0.0); 
        (C[9] *> O[5])=(0.0,0.0); 
        (C[9] *> O[6])=(0.0,0.0); 
        (C[9] *> O[7])=(0.0,0.0); 
        (C[9] *> O[8])=(0.0,0.0); 
        (C[9] *> O[9])=(0.0,0.0); 
        (C[9] *> O[10])=(0.0,0.0); 
        (C[9] *> O[11])=(0.0,0.0); 
        (C[9] *> O[12])=(0.0,0.0); 
        (C[9] *> O[13])=(0.0,0.0); 
        (C[9] *> O[14])=(0.0,0.0); 
        (C[9] *> O[15])=(0.0,0.0); 
        (C[9] *> O[16])=(0.0,0.0); 
        (C[9] *> O[17])=(0.0,0.0); 
        (C[9] *> O[18])=(0.0,0.0); 
        (C[9] *> O[19])=(0.0,0.0); 
        (C[9] *> O[20])=(0.0,0.0); 
        (C[9] *> O[21])=(0.0,0.0); 
        (C[9] *> O[22])=(0.0,0.0); 
        (C[9] *> O[23])=(0.0,0.0); 
        (C[9] *> O[24])=(0.0,0.0); 
        (C[9] *> O[25])=(0.0,0.0); 
        (C[9] *> O[26])=(0.0,0.0); 
        (C[9] *> O[27])=(0.0,0.0); 
        (C[9] *> O[28])=(0.0,0.0); 
        (C[9] *> O[29])=(0.0,0.0); 
        (C[9] *> O[30])=(0.0,0.0); 
        (C[9] *> O[31])=(0.0,0.0); 
        (C[10] *> O[0])=(0.0,0.0); 
        (C[10] *> O[1])=(0.0,0.0); 
        (C[10] *> O[2])=(0.0,0.0); 
        (C[10] *> O[3])=(0.0,0.0); 
        (C[10] *> O[4])=(0.0,0.0); 
        (C[10] *> O[5])=(0.0,0.0); 
        (C[10] *> O[6])=(0.0,0.0); 
        (C[10] *> O[7])=(0.0,0.0); 
        (C[10] *> O[8])=(0.0,0.0); 
        (C[10] *> O[9])=(0.0,0.0); 
        (C[10] *> O[10])=(0.0,0.0); 
        (C[10] *> O[11])=(0.0,0.0); 
        (C[10] *> O[12])=(0.0,0.0); 
        (C[10] *> O[13])=(0.0,0.0); 
        (C[10] *> O[14])=(0.0,0.0); 
        (C[10] *> O[15])=(0.0,0.0); 
        (C[10] *> O[16])=(0.0,0.0); 
        (C[10] *> O[17])=(0.0,0.0); 
        (C[10] *> O[18])=(0.0,0.0); 
        (C[10] *> O[19])=(0.0,0.0); 
        (C[10] *> O[20])=(0.0,0.0); 
        (C[10] *> O[21])=(0.0,0.0); 
        (C[10] *> O[22])=(0.0,0.0); 
        (C[10] *> O[23])=(0.0,0.0); 
        (C[10] *> O[24])=(0.0,0.0); 
        (C[10] *> O[25])=(0.0,0.0); 
        (C[10] *> O[26])=(0.0,0.0); 
        (C[10] *> O[27])=(0.0,0.0); 
        (C[10] *> O[28])=(0.0,0.0); 
        (C[10] *> O[29])=(0.0,0.0); 
        (C[10] *> O[30])=(0.0,0.0); 
        (C[10] *> O[31])=(0.0,0.0); 
        (C[11] *> O[0])=(0.0,0.0); 
        (C[11] *> O[1])=(0.0,0.0); 
        (C[11] *> O[2])=(0.0,0.0); 
        (C[11] *> O[3])=(0.0,0.0); 
        (C[11] *> O[4])=(0.0,0.0); 
        (C[11] *> O[5])=(0.0,0.0); 
        (C[11] *> O[6])=(0.0,0.0); 
        (C[11] *> O[7])=(0.0,0.0); 
        (C[11] *> O[8])=(0.0,0.0); 
        (C[11] *> O[9])=(0.0,0.0); 
        (C[11] *> O[10])=(0.0,0.0); 
        (C[11] *> O[11])=(0.0,0.0); 
        (C[11] *> O[12])=(0.0,0.0); 
        (C[11] *> O[13])=(0.0,0.0); 
        (C[11] *> O[14])=(0.0,0.0); 
        (C[11] *> O[15])=(0.0,0.0); 
        (C[11] *> O[16])=(0.0,0.0); 
        (C[11] *> O[17])=(0.0,0.0); 
        (C[11] *> O[18])=(0.0,0.0); 
        (C[11] *> O[19])=(0.0,0.0); 
        (C[11] *> O[20])=(0.0,0.0); 
        (C[11] *> O[21])=(0.0,0.0); 
        (C[11] *> O[22])=(0.0,0.0); 
        (C[11] *> O[23])=(0.0,0.0); 
        (C[11] *> O[24])=(0.0,0.0); 
        (C[11] *> O[25])=(0.0,0.0); 
        (C[11] *> O[26])=(0.0,0.0); 
        (C[11] *> O[27])=(0.0,0.0); 
        (C[11] *> O[28])=(0.0,0.0); 
        (C[11] *> O[29])=(0.0,0.0); 
        (C[11] *> O[30])=(0.0,0.0); 
        (C[11] *> O[31])=(0.0,0.0); 
        (C[12] *> O[0])=(0.0,0.0); 
        (C[12] *> O[1])=(0.0,0.0); 
        (C[12] *> O[2])=(0.0,0.0); 
        (C[12] *> O[3])=(0.0,0.0); 
        (C[12] *> O[4])=(0.0,0.0); 
        (C[12] *> O[5])=(0.0,0.0); 
        (C[12] *> O[6])=(0.0,0.0); 
        (C[12] *> O[7])=(0.0,0.0); 
        (C[12] *> O[8])=(0.0,0.0); 
        (C[12] *> O[9])=(0.0,0.0); 
        (C[12] *> O[10])=(0.0,0.0); 
        (C[12] *> O[11])=(0.0,0.0); 
        (C[12] *> O[12])=(0.0,0.0); 
        (C[12] *> O[13])=(0.0,0.0); 
        (C[12] *> O[14])=(0.0,0.0); 
        (C[12] *> O[15])=(0.0,0.0); 
        (C[12] *> O[16])=(0.0,0.0); 
        (C[12] *> O[17])=(0.0,0.0); 
        (C[12] *> O[18])=(0.0,0.0); 
        (C[12] *> O[19])=(0.0,0.0); 
        (C[12] *> O[20])=(0.0,0.0); 
        (C[12] *> O[21])=(0.0,0.0); 
        (C[12] *> O[22])=(0.0,0.0); 
        (C[12] *> O[23])=(0.0,0.0); 
        (C[12] *> O[24])=(0.0,0.0); 
        (C[12] *> O[25])=(0.0,0.0); 
        (C[12] *> O[26])=(0.0,0.0); 
        (C[12] *> O[27])=(0.0,0.0); 
        (C[12] *> O[28])=(0.0,0.0); 
        (C[12] *> O[29])=(0.0,0.0); 
        (C[12] *> O[30])=(0.0,0.0); 
        (C[12] *> O[31])=(0.0,0.0); 
        (C[13] *> O[0])=(0.0,0.0); 
        (C[13] *> O[1])=(0.0,0.0); 
        (C[13] *> O[2])=(0.0,0.0); 
        (C[13] *> O[3])=(0.0,0.0); 
        (C[13] *> O[4])=(0.0,0.0); 
        (C[13] *> O[5])=(0.0,0.0); 
        (C[13] *> O[6])=(0.0,0.0); 
        (C[13] *> O[7])=(0.0,0.0); 
        (C[13] *> O[8])=(0.0,0.0); 
        (C[13] *> O[9])=(0.0,0.0); 
        (C[13] *> O[10])=(0.0,0.0); 
        (C[13] *> O[11])=(0.0,0.0); 
        (C[13] *> O[12])=(0.0,0.0); 
        (C[13] *> O[13])=(0.0,0.0); 
        (C[13] *> O[14])=(0.0,0.0); 
        (C[13] *> O[15])=(0.0,0.0); 
        (C[13] *> O[16])=(0.0,0.0); 
        (C[13] *> O[17])=(0.0,0.0); 
        (C[13] *> O[18])=(0.0,0.0); 
        (C[13] *> O[19])=(0.0,0.0); 
        (C[13] *> O[20])=(0.0,0.0); 
        (C[13] *> O[21])=(0.0,0.0); 
        (C[13] *> O[22])=(0.0,0.0); 
        (C[13] *> O[23])=(0.0,0.0); 
        (C[13] *> O[24])=(0.0,0.0); 
        (C[13] *> O[25])=(0.0,0.0); 
        (C[13] *> O[26])=(0.0,0.0); 
        (C[13] *> O[27])=(0.0,0.0); 
        (C[13] *> O[28])=(0.0,0.0); 
        (C[13] *> O[29])=(0.0,0.0); 
        (C[13] *> O[30])=(0.0,0.0); 
        (C[13] *> O[31])=(0.0,0.0); 
        (C[14] *> O[0])=(0.0,0.0); 
        (C[14] *> O[1])=(0.0,0.0); 
        (C[14] *> O[2])=(0.0,0.0); 
        (C[14] *> O[3])=(0.0,0.0); 
        (C[14] *> O[4])=(0.0,0.0); 
        (C[14] *> O[5])=(0.0,0.0); 
        (C[14] *> O[6])=(0.0,0.0); 
        (C[14] *> O[7])=(0.0,0.0); 
        (C[14] *> O[8])=(0.0,0.0); 
        (C[14] *> O[9])=(0.0,0.0); 
        (C[14] *> O[10])=(0.0,0.0); 
        (C[14] *> O[11])=(0.0,0.0); 
        (C[14] *> O[12])=(0.0,0.0); 
        (C[14] *> O[13])=(0.0,0.0); 
        (C[14] *> O[14])=(0.0,0.0); 
        (C[14] *> O[15])=(0.0,0.0); 
        (C[14] *> O[16])=(0.0,0.0); 
        (C[14] *> O[17])=(0.0,0.0); 
        (C[14] *> O[18])=(0.0,0.0); 
        (C[14] *> O[19])=(0.0,0.0); 
        (C[14] *> O[20])=(0.0,0.0); 
        (C[14] *> O[21])=(0.0,0.0); 
        (C[14] *> O[22])=(0.0,0.0); 
        (C[14] *> O[23])=(0.0,0.0); 
        (C[14] *> O[24])=(0.0,0.0); 
        (C[14] *> O[25])=(0.0,0.0); 
        (C[14] *> O[26])=(0.0,0.0); 
        (C[14] *> O[27])=(0.0,0.0); 
        (C[14] *> O[28])=(0.0,0.0); 
        (C[14] *> O[29])=(0.0,0.0); 
        (C[14] *> O[30])=(0.0,0.0); 
        (C[14] *> O[31])=(0.0,0.0); 
        (C[15] *> O[0])=(0.0,0.0); 
        (C[15] *> O[1])=(0.0,0.0); 
        (C[15] *> O[2])=(0.0,0.0); 
        (C[15] *> O[3])=(0.0,0.0); 
        (C[15] *> O[4])=(0.0,0.0); 
        (C[15] *> O[5])=(0.0,0.0); 
        (C[15] *> O[6])=(0.0,0.0); 
        (C[15] *> O[7])=(0.0,0.0); 
        (C[15] *> O[8])=(0.0,0.0); 
        (C[15] *> O[9])=(0.0,0.0); 
        (C[15] *> O[10])=(0.0,0.0); 
        (C[15] *> O[11])=(0.0,0.0); 
        (C[15] *> O[12])=(0.0,0.0); 
        (C[15] *> O[13])=(0.0,0.0); 
        (C[15] *> O[14])=(0.0,0.0); 
        (C[15] *> O[15])=(0.0,0.0); 
        (C[15] *> O[16])=(0.0,0.0); 
        (C[15] *> O[17])=(0.0,0.0); 
        (C[15] *> O[18])=(0.0,0.0); 
        (C[15] *> O[19])=(0.0,0.0); 
        (C[15] *> O[20])=(0.0,0.0); 
        (C[15] *> O[21])=(0.0,0.0); 
        (C[15] *> O[22])=(0.0,0.0); 
        (C[15] *> O[23])=(0.0,0.0); 
        (C[15] *> O[24])=(0.0,0.0); 
        (C[15] *> O[25])=(0.0,0.0); 
        (C[15] *> O[26])=(0.0,0.0); 
        (C[15] *> O[27])=(0.0,0.0); 
        (C[15] *> O[28])=(0.0,0.0); 
        (C[15] *> O[29])=(0.0,0.0); 
        (C[15] *> O[30])=(0.0,0.0); 
        (C[15] *> O[31])=(0.0,0.0); 
        (D[0] *> O[0])=(0.0,0.0); 
        (D[0] *> O[1])=(0.0,0.0); 
        (D[0] *> O[2])=(0.0,0.0); 
        (D[0] *> O[3])=(0.0,0.0); 
        (D[0] *> O[4])=(0.0,0.0); 
        (D[0] *> O[5])=(0.0,0.0); 
        (D[0] *> O[6])=(0.0,0.0); 
        (D[0] *> O[7])=(0.0,0.0); 
        (D[0] *> O[8])=(0.0,0.0); 
        (D[0] *> O[9])=(0.0,0.0); 
        (D[0] *> O[10])=(0.0,0.0); 
        (D[0] *> O[11])=(0.0,0.0); 
        (D[0] *> O[12])=(0.0,0.0); 
        (D[0] *> O[13])=(0.0,0.0); 
        (D[0] *> O[14])=(0.0,0.0); 
        (D[0] *> O[15])=(0.0,0.0); 
        (D[0] *> O[16])=(0.0,0.0); 
        (D[0] *> O[17])=(0.0,0.0); 
        (D[0] *> O[18])=(0.0,0.0); 
        (D[0] *> O[19])=(0.0,0.0); 
        (D[0] *> O[20])=(0.0,0.0); 
        (D[0] *> O[21])=(0.0,0.0); 
        (D[0] *> O[22])=(0.0,0.0); 
        (D[0] *> O[23])=(0.0,0.0); 
        (D[0] *> O[24])=(0.0,0.0); 
        (D[0] *> O[25])=(0.0,0.0); 
        (D[0] *> O[26])=(0.0,0.0); 
        (D[0] *> O[27])=(0.0,0.0); 
        (D[0] *> O[28])=(0.0,0.0); 
        (D[0] *> O[29])=(0.0,0.0); 
        (D[0] *> O[30])=(0.0,0.0); 
        (D[0] *> O[31])=(0.0,0.0); 
        (D[1] *> O[0])=(0.0,0.0); 
        (D[1] *> O[1])=(0.0,0.0); 
        (D[1] *> O[2])=(0.0,0.0); 
        (D[1] *> O[3])=(0.0,0.0); 
        (D[1] *> O[4])=(0.0,0.0); 
        (D[1] *> O[5])=(0.0,0.0); 
        (D[1] *> O[6])=(0.0,0.0); 
        (D[1] *> O[7])=(0.0,0.0); 
        (D[1] *> O[8])=(0.0,0.0); 
        (D[1] *> O[9])=(0.0,0.0); 
        (D[1] *> O[10])=(0.0,0.0); 
        (D[1] *> O[11])=(0.0,0.0); 
        (D[1] *> O[12])=(0.0,0.0); 
        (D[1] *> O[13])=(0.0,0.0); 
        (D[1] *> O[14])=(0.0,0.0); 
        (D[1] *> O[15])=(0.0,0.0); 
        (D[1] *> O[16])=(0.0,0.0); 
        (D[1] *> O[17])=(0.0,0.0); 
        (D[1] *> O[18])=(0.0,0.0); 
        (D[1] *> O[19])=(0.0,0.0); 
        (D[1] *> O[20])=(0.0,0.0); 
        (D[1] *> O[21])=(0.0,0.0); 
        (D[1] *> O[22])=(0.0,0.0); 
        (D[1] *> O[23])=(0.0,0.0); 
        (D[1] *> O[24])=(0.0,0.0); 
        (D[1] *> O[25])=(0.0,0.0); 
        (D[1] *> O[26])=(0.0,0.0); 
        (D[1] *> O[27])=(0.0,0.0); 
        (D[1] *> O[28])=(0.0,0.0); 
        (D[1] *> O[29])=(0.0,0.0); 
        (D[1] *> O[30])=(0.0,0.0); 
        (D[1] *> O[31])=(0.0,0.0); 
        (D[2] *> O[0])=(0.0,0.0); 
        (D[2] *> O[1])=(0.0,0.0); 
        (D[2] *> O[2])=(0.0,0.0); 
        (D[2] *> O[3])=(0.0,0.0); 
        (D[2] *> O[4])=(0.0,0.0); 
        (D[2] *> O[5])=(0.0,0.0); 
        (D[2] *> O[6])=(0.0,0.0); 
        (D[2] *> O[7])=(0.0,0.0); 
        (D[2] *> O[8])=(0.0,0.0); 
        (D[2] *> O[9])=(0.0,0.0); 
        (D[2] *> O[10])=(0.0,0.0); 
        (D[2] *> O[11])=(0.0,0.0); 
        (D[2] *> O[12])=(0.0,0.0); 
        (D[2] *> O[13])=(0.0,0.0); 
        (D[2] *> O[14])=(0.0,0.0); 
        (D[2] *> O[15])=(0.0,0.0); 
        (D[2] *> O[16])=(0.0,0.0); 
        (D[2] *> O[17])=(0.0,0.0); 
        (D[2] *> O[18])=(0.0,0.0); 
        (D[2] *> O[19])=(0.0,0.0); 
        (D[2] *> O[20])=(0.0,0.0); 
        (D[2] *> O[21])=(0.0,0.0); 
        (D[2] *> O[22])=(0.0,0.0); 
        (D[2] *> O[23])=(0.0,0.0); 
        (D[2] *> O[24])=(0.0,0.0); 
        (D[2] *> O[25])=(0.0,0.0); 
        (D[2] *> O[26])=(0.0,0.0); 
        (D[2] *> O[27])=(0.0,0.0); 
        (D[2] *> O[28])=(0.0,0.0); 
        (D[2] *> O[29])=(0.0,0.0); 
        (D[2] *> O[30])=(0.0,0.0); 
        (D[2] *> O[31])=(0.0,0.0); 
        (D[3] *> O[0])=(0.0,0.0); 
        (D[3] *> O[1])=(0.0,0.0); 
        (D[3] *> O[2])=(0.0,0.0); 
        (D[3] *> O[3])=(0.0,0.0); 
        (D[3] *> O[4])=(0.0,0.0); 
        (D[3] *> O[5])=(0.0,0.0); 
        (D[3] *> O[6])=(0.0,0.0); 
        (D[3] *> O[7])=(0.0,0.0); 
        (D[3] *> O[8])=(0.0,0.0); 
        (D[3] *> O[9])=(0.0,0.0); 
        (D[3] *> O[10])=(0.0,0.0); 
        (D[3] *> O[11])=(0.0,0.0); 
        (D[3] *> O[12])=(0.0,0.0); 
        (D[3] *> O[13])=(0.0,0.0); 
        (D[3] *> O[14])=(0.0,0.0); 
        (D[3] *> O[15])=(0.0,0.0); 
        (D[3] *> O[16])=(0.0,0.0); 
        (D[3] *> O[17])=(0.0,0.0); 
        (D[3] *> O[18])=(0.0,0.0); 
        (D[3] *> O[19])=(0.0,0.0); 
        (D[3] *> O[20])=(0.0,0.0); 
        (D[3] *> O[21])=(0.0,0.0); 
        (D[3] *> O[22])=(0.0,0.0); 
        (D[3] *> O[23])=(0.0,0.0); 
        (D[3] *> O[24])=(0.0,0.0); 
        (D[3] *> O[25])=(0.0,0.0); 
        (D[3] *> O[26])=(0.0,0.0); 
        (D[3] *> O[27])=(0.0,0.0); 
        (D[3] *> O[28])=(0.0,0.0); 
        (D[3] *> O[29])=(0.0,0.0); 
        (D[3] *> O[30])=(0.0,0.0); 
        (D[3] *> O[31])=(0.0,0.0); 
        (D[4] *> O[0])=(0.0,0.0); 
        (D[4] *> O[1])=(0.0,0.0); 
        (D[4] *> O[2])=(0.0,0.0); 
        (D[4] *> O[3])=(0.0,0.0); 
        (D[4] *> O[4])=(0.0,0.0); 
        (D[4] *> O[5])=(0.0,0.0); 
        (D[4] *> O[6])=(0.0,0.0); 
        (D[4] *> O[7])=(0.0,0.0); 
        (D[4] *> O[8])=(0.0,0.0); 
        (D[4] *> O[9])=(0.0,0.0); 
        (D[4] *> O[10])=(0.0,0.0); 
        (D[4] *> O[11])=(0.0,0.0); 
        (D[4] *> O[12])=(0.0,0.0); 
        (D[4] *> O[13])=(0.0,0.0); 
        (D[4] *> O[14])=(0.0,0.0); 
        (D[4] *> O[15])=(0.0,0.0); 
        (D[4] *> O[16])=(0.0,0.0); 
        (D[4] *> O[17])=(0.0,0.0); 
        (D[4] *> O[18])=(0.0,0.0); 
        (D[4] *> O[19])=(0.0,0.0); 
        (D[4] *> O[20])=(0.0,0.0); 
        (D[4] *> O[21])=(0.0,0.0); 
        (D[4] *> O[22])=(0.0,0.0); 
        (D[4] *> O[23])=(0.0,0.0); 
        (D[4] *> O[24])=(0.0,0.0); 
        (D[4] *> O[25])=(0.0,0.0); 
        (D[4] *> O[26])=(0.0,0.0); 
        (D[4] *> O[27])=(0.0,0.0); 
        (D[4] *> O[28])=(0.0,0.0); 
        (D[4] *> O[29])=(0.0,0.0); 
        (D[4] *> O[30])=(0.0,0.0); 
        (D[4] *> O[31])=(0.0,0.0); 
        (D[5] *> O[0])=(0.0,0.0); 
        (D[5] *> O[1])=(0.0,0.0); 
        (D[5] *> O[2])=(0.0,0.0); 
        (D[5] *> O[3])=(0.0,0.0); 
        (D[5] *> O[4])=(0.0,0.0); 
        (D[5] *> O[5])=(0.0,0.0); 
        (D[5] *> O[6])=(0.0,0.0); 
        (D[5] *> O[7])=(0.0,0.0); 
        (D[5] *> O[8])=(0.0,0.0); 
        (D[5] *> O[9])=(0.0,0.0); 
        (D[5] *> O[10])=(0.0,0.0); 
        (D[5] *> O[11])=(0.0,0.0); 
        (D[5] *> O[12])=(0.0,0.0); 
        (D[5] *> O[13])=(0.0,0.0); 
        (D[5] *> O[14])=(0.0,0.0); 
        (D[5] *> O[15])=(0.0,0.0); 
        (D[5] *> O[16])=(0.0,0.0); 
        (D[5] *> O[17])=(0.0,0.0); 
        (D[5] *> O[18])=(0.0,0.0); 
        (D[5] *> O[19])=(0.0,0.0); 
        (D[5] *> O[20])=(0.0,0.0); 
        (D[5] *> O[21])=(0.0,0.0); 
        (D[5] *> O[22])=(0.0,0.0); 
        (D[5] *> O[23])=(0.0,0.0); 
        (D[5] *> O[24])=(0.0,0.0); 
        (D[5] *> O[25])=(0.0,0.0); 
        (D[5] *> O[26])=(0.0,0.0); 
        (D[5] *> O[27])=(0.0,0.0); 
        (D[5] *> O[28])=(0.0,0.0); 
        (D[5] *> O[29])=(0.0,0.0); 
        (D[5] *> O[30])=(0.0,0.0); 
        (D[5] *> O[31])=(0.0,0.0); 
        (D[6] *> O[0])=(0.0,0.0); 
        (D[6] *> O[1])=(0.0,0.0); 
        (D[6] *> O[2])=(0.0,0.0); 
        (D[6] *> O[3])=(0.0,0.0); 
        (D[6] *> O[4])=(0.0,0.0); 
        (D[6] *> O[5])=(0.0,0.0); 
        (D[6] *> O[6])=(0.0,0.0); 
        (D[6] *> O[7])=(0.0,0.0); 
        (D[6] *> O[8])=(0.0,0.0); 
        (D[6] *> O[9])=(0.0,0.0); 
        (D[6] *> O[10])=(0.0,0.0); 
        (D[6] *> O[11])=(0.0,0.0); 
        (D[6] *> O[12])=(0.0,0.0); 
        (D[6] *> O[13])=(0.0,0.0); 
        (D[6] *> O[14])=(0.0,0.0); 
        (D[6] *> O[15])=(0.0,0.0); 
        (D[6] *> O[16])=(0.0,0.0); 
        (D[6] *> O[17])=(0.0,0.0); 
        (D[6] *> O[18])=(0.0,0.0); 
        (D[6] *> O[19])=(0.0,0.0); 
        (D[6] *> O[20])=(0.0,0.0); 
        (D[6] *> O[21])=(0.0,0.0); 
        (D[6] *> O[22])=(0.0,0.0); 
        (D[6] *> O[23])=(0.0,0.0); 
        (D[6] *> O[24])=(0.0,0.0); 
        (D[6] *> O[25])=(0.0,0.0); 
        (D[6] *> O[26])=(0.0,0.0); 
        (D[6] *> O[27])=(0.0,0.0); 
        (D[6] *> O[28])=(0.0,0.0); 
        (D[6] *> O[29])=(0.0,0.0); 
        (D[6] *> O[30])=(0.0,0.0); 
        (D[6] *> O[31])=(0.0,0.0); 
        (D[7] *> O[0])=(0.0,0.0); 
        (D[7] *> O[1])=(0.0,0.0); 
        (D[7] *> O[2])=(0.0,0.0); 
        (D[7] *> O[3])=(0.0,0.0); 
        (D[7] *> O[4])=(0.0,0.0); 
        (D[7] *> O[5])=(0.0,0.0); 
        (D[7] *> O[6])=(0.0,0.0); 
        (D[7] *> O[7])=(0.0,0.0); 
        (D[7] *> O[8])=(0.0,0.0); 
        (D[7] *> O[9])=(0.0,0.0); 
        (D[7] *> O[10])=(0.0,0.0); 
        (D[7] *> O[11])=(0.0,0.0); 
        (D[7] *> O[12])=(0.0,0.0); 
        (D[7] *> O[13])=(0.0,0.0); 
        (D[7] *> O[14])=(0.0,0.0); 
        (D[7] *> O[15])=(0.0,0.0); 
        (D[7] *> O[16])=(0.0,0.0); 
        (D[7] *> O[17])=(0.0,0.0); 
        (D[7] *> O[18])=(0.0,0.0); 
        (D[7] *> O[19])=(0.0,0.0); 
        (D[7] *> O[20])=(0.0,0.0); 
        (D[7] *> O[21])=(0.0,0.0); 
        (D[7] *> O[22])=(0.0,0.0); 
        (D[7] *> O[23])=(0.0,0.0); 
        (D[7] *> O[24])=(0.0,0.0); 
        (D[7] *> O[25])=(0.0,0.0); 
        (D[7] *> O[26])=(0.0,0.0); 
        (D[7] *> O[27])=(0.0,0.0); 
        (D[7] *> O[28])=(0.0,0.0); 
        (D[7] *> O[29])=(0.0,0.0); 
        (D[7] *> O[30])=(0.0,0.0); 
        (D[7] *> O[31])=(0.0,0.0); 
        (D[8] *> O[0])=(0.0,0.0); 
        (D[8] *> O[1])=(0.0,0.0); 
        (D[8] *> O[2])=(0.0,0.0); 
        (D[8] *> O[3])=(0.0,0.0); 
        (D[8] *> O[4])=(0.0,0.0); 
        (D[8] *> O[5])=(0.0,0.0); 
        (D[8] *> O[6])=(0.0,0.0); 
        (D[8] *> O[7])=(0.0,0.0); 
        (D[8] *> O[8])=(0.0,0.0); 
        (D[8] *> O[9])=(0.0,0.0); 
        (D[8] *> O[10])=(0.0,0.0); 
        (D[8] *> O[11])=(0.0,0.0); 
        (D[8] *> O[12])=(0.0,0.0); 
        (D[8] *> O[13])=(0.0,0.0); 
        (D[8] *> O[14])=(0.0,0.0); 
        (D[8] *> O[15])=(0.0,0.0); 
        (D[8] *> O[16])=(0.0,0.0); 
        (D[8] *> O[17])=(0.0,0.0); 
        (D[8] *> O[18])=(0.0,0.0); 
        (D[8] *> O[19])=(0.0,0.0); 
        (D[8] *> O[20])=(0.0,0.0); 
        (D[8] *> O[21])=(0.0,0.0); 
        (D[8] *> O[22])=(0.0,0.0); 
        (D[8] *> O[23])=(0.0,0.0); 
        (D[8] *> O[24])=(0.0,0.0); 
        (D[8] *> O[25])=(0.0,0.0); 
        (D[8] *> O[26])=(0.0,0.0); 
        (D[8] *> O[27])=(0.0,0.0); 
        (D[8] *> O[28])=(0.0,0.0); 
        (D[8] *> O[29])=(0.0,0.0); 
        (D[8] *> O[30])=(0.0,0.0); 
        (D[8] *> O[31])=(0.0,0.0); 
        (D[9] *> O[0])=(0.0,0.0); 
        (D[9] *> O[1])=(0.0,0.0); 
        (D[9] *> O[2])=(0.0,0.0); 
        (D[9] *> O[3])=(0.0,0.0); 
        (D[9] *> O[4])=(0.0,0.0); 
        (D[9] *> O[5])=(0.0,0.0); 
        (D[9] *> O[6])=(0.0,0.0); 
        (D[9] *> O[7])=(0.0,0.0); 
        (D[9] *> O[8])=(0.0,0.0); 
        (D[9] *> O[9])=(0.0,0.0); 
        (D[9] *> O[10])=(0.0,0.0); 
        (D[9] *> O[11])=(0.0,0.0); 
        (D[9] *> O[12])=(0.0,0.0); 
        (D[9] *> O[13])=(0.0,0.0); 
        (D[9] *> O[14])=(0.0,0.0); 
        (D[9] *> O[15])=(0.0,0.0); 
        (D[9] *> O[16])=(0.0,0.0); 
        (D[9] *> O[17])=(0.0,0.0); 
        (D[9] *> O[18])=(0.0,0.0); 
        (D[9] *> O[19])=(0.0,0.0); 
        (D[9] *> O[20])=(0.0,0.0); 
        (D[9] *> O[21])=(0.0,0.0); 
        (D[9] *> O[22])=(0.0,0.0); 
        (D[9] *> O[23])=(0.0,0.0); 
        (D[9] *> O[24])=(0.0,0.0); 
        (D[9] *> O[25])=(0.0,0.0); 
        (D[9] *> O[26])=(0.0,0.0); 
        (D[9] *> O[27])=(0.0,0.0); 
        (D[9] *> O[28])=(0.0,0.0); 
        (D[9] *> O[29])=(0.0,0.0); 
        (D[9] *> O[30])=(0.0,0.0); 
        (D[9] *> O[31])=(0.0,0.0); 
        (D[10] *> O[0])=(0.0,0.0); 
        (D[10] *> O[1])=(0.0,0.0); 
        (D[10] *> O[2])=(0.0,0.0); 
        (D[10] *> O[3])=(0.0,0.0); 
        (D[10] *> O[4])=(0.0,0.0); 
        (D[10] *> O[5])=(0.0,0.0); 
        (D[10] *> O[6])=(0.0,0.0); 
        (D[10] *> O[7])=(0.0,0.0); 
        (D[10] *> O[8])=(0.0,0.0); 
        (D[10] *> O[9])=(0.0,0.0); 
        (D[10] *> O[10])=(0.0,0.0); 
        (D[10] *> O[11])=(0.0,0.0); 
        (D[10] *> O[12])=(0.0,0.0); 
        (D[10] *> O[13])=(0.0,0.0); 
        (D[10] *> O[14])=(0.0,0.0); 
        (D[10] *> O[15])=(0.0,0.0); 
        (D[10] *> O[16])=(0.0,0.0); 
        (D[10] *> O[17])=(0.0,0.0); 
        (D[10] *> O[18])=(0.0,0.0); 
        (D[10] *> O[19])=(0.0,0.0); 
        (D[10] *> O[20])=(0.0,0.0); 
        (D[10] *> O[21])=(0.0,0.0); 
        (D[10] *> O[22])=(0.0,0.0); 
        (D[10] *> O[23])=(0.0,0.0); 
        (D[10] *> O[24])=(0.0,0.0); 
        (D[10] *> O[25])=(0.0,0.0); 
        (D[10] *> O[26])=(0.0,0.0); 
        (D[10] *> O[27])=(0.0,0.0); 
        (D[10] *> O[28])=(0.0,0.0); 
        (D[10] *> O[29])=(0.0,0.0); 
        (D[10] *> O[30])=(0.0,0.0); 
        (D[10] *> O[31])=(0.0,0.0); 
        (D[11] *> O[0])=(0.0,0.0); 
        (D[11] *> O[1])=(0.0,0.0); 
        (D[11] *> O[2])=(0.0,0.0); 
        (D[11] *> O[3])=(0.0,0.0); 
        (D[11] *> O[4])=(0.0,0.0); 
        (D[11] *> O[5])=(0.0,0.0); 
        (D[11] *> O[6])=(0.0,0.0); 
        (D[11] *> O[7])=(0.0,0.0); 
        (D[11] *> O[8])=(0.0,0.0); 
        (D[11] *> O[9])=(0.0,0.0); 
        (D[11] *> O[10])=(0.0,0.0); 
        (D[11] *> O[11])=(0.0,0.0); 
        (D[11] *> O[12])=(0.0,0.0); 
        (D[11] *> O[13])=(0.0,0.0); 
        (D[11] *> O[14])=(0.0,0.0); 
        (D[11] *> O[15])=(0.0,0.0); 
        (D[11] *> O[16])=(0.0,0.0); 
        (D[11] *> O[17])=(0.0,0.0); 
        (D[11] *> O[18])=(0.0,0.0); 
        (D[11] *> O[19])=(0.0,0.0); 
        (D[11] *> O[20])=(0.0,0.0); 
        (D[11] *> O[21])=(0.0,0.0); 
        (D[11] *> O[22])=(0.0,0.0); 
        (D[11] *> O[23])=(0.0,0.0); 
        (D[11] *> O[24])=(0.0,0.0); 
        (D[11] *> O[25])=(0.0,0.0); 
        (D[11] *> O[26])=(0.0,0.0); 
        (D[11] *> O[27])=(0.0,0.0); 
        (D[11] *> O[28])=(0.0,0.0); 
        (D[11] *> O[29])=(0.0,0.0); 
        (D[11] *> O[30])=(0.0,0.0); 
        (D[11] *> O[31])=(0.0,0.0); 
        (D[12] *> O[0])=(0.0,0.0); 
        (D[12] *> O[1])=(0.0,0.0); 
        (D[12] *> O[2])=(0.0,0.0); 
        (D[12] *> O[3])=(0.0,0.0); 
        (D[12] *> O[4])=(0.0,0.0); 
        (D[12] *> O[5])=(0.0,0.0); 
        (D[12] *> O[6])=(0.0,0.0); 
        (D[12] *> O[7])=(0.0,0.0); 
        (D[12] *> O[8])=(0.0,0.0); 
        (D[12] *> O[9])=(0.0,0.0); 
        (D[12] *> O[10])=(0.0,0.0); 
        (D[12] *> O[11])=(0.0,0.0); 
        (D[12] *> O[12])=(0.0,0.0); 
        (D[12] *> O[13])=(0.0,0.0); 
        (D[12] *> O[14])=(0.0,0.0); 
        (D[12] *> O[15])=(0.0,0.0); 
        (D[12] *> O[16])=(0.0,0.0); 
        (D[12] *> O[17])=(0.0,0.0); 
        (D[12] *> O[18])=(0.0,0.0); 
        (D[12] *> O[19])=(0.0,0.0); 
        (D[12] *> O[20])=(0.0,0.0); 
        (D[12] *> O[21])=(0.0,0.0); 
        (D[12] *> O[22])=(0.0,0.0); 
        (D[12] *> O[23])=(0.0,0.0); 
        (D[12] *> O[24])=(0.0,0.0); 
        (D[12] *> O[25])=(0.0,0.0); 
        (D[12] *> O[26])=(0.0,0.0); 
        (D[12] *> O[27])=(0.0,0.0); 
        (D[12] *> O[28])=(0.0,0.0); 
        (D[12] *> O[29])=(0.0,0.0); 
        (D[12] *> O[30])=(0.0,0.0); 
        (D[12] *> O[31])=(0.0,0.0); 
        (D[13] *> O[0])=(0.0,0.0); 
        (D[13] *> O[1])=(0.0,0.0); 
        (D[13] *> O[2])=(0.0,0.0); 
        (D[13] *> O[3])=(0.0,0.0); 
        (D[13] *> O[4])=(0.0,0.0); 
        (D[13] *> O[5])=(0.0,0.0); 
        (D[13] *> O[6])=(0.0,0.0); 
        (D[13] *> O[7])=(0.0,0.0); 
        (D[13] *> O[8])=(0.0,0.0); 
        (D[13] *> O[9])=(0.0,0.0); 
        (D[13] *> O[10])=(0.0,0.0); 
        (D[13] *> O[11])=(0.0,0.0); 
        (D[13] *> O[12])=(0.0,0.0); 
        (D[13] *> O[13])=(0.0,0.0); 
        (D[13] *> O[14])=(0.0,0.0); 
        (D[13] *> O[15])=(0.0,0.0); 
        (D[13] *> O[16])=(0.0,0.0); 
        (D[13] *> O[17])=(0.0,0.0); 
        (D[13] *> O[18])=(0.0,0.0); 
        (D[13] *> O[19])=(0.0,0.0); 
        (D[13] *> O[20])=(0.0,0.0); 
        (D[13] *> O[21])=(0.0,0.0); 
        (D[13] *> O[22])=(0.0,0.0); 
        (D[13] *> O[23])=(0.0,0.0); 
        (D[13] *> O[24])=(0.0,0.0); 
        (D[13] *> O[25])=(0.0,0.0); 
        (D[13] *> O[26])=(0.0,0.0); 
        (D[13] *> O[27])=(0.0,0.0); 
        (D[13] *> O[28])=(0.0,0.0); 
        (D[13] *> O[29])=(0.0,0.0); 
        (D[13] *> O[30])=(0.0,0.0); 
        (D[13] *> O[31])=(0.0,0.0); 
        (D[14] *> O[0])=(0.0,0.0); 
        (D[14] *> O[1])=(0.0,0.0); 
        (D[14] *> O[2])=(0.0,0.0); 
        (D[14] *> O[3])=(0.0,0.0); 
        (D[14] *> O[4])=(0.0,0.0); 
        (D[14] *> O[5])=(0.0,0.0); 
        (D[14] *> O[6])=(0.0,0.0); 
        (D[14] *> O[7])=(0.0,0.0); 
        (D[14] *> O[8])=(0.0,0.0); 
        (D[14] *> O[9])=(0.0,0.0); 
        (D[14] *> O[10])=(0.0,0.0); 
        (D[14] *> O[11])=(0.0,0.0); 
        (D[14] *> O[12])=(0.0,0.0); 
        (D[14] *> O[13])=(0.0,0.0); 
        (D[14] *> O[14])=(0.0,0.0); 
        (D[14] *> O[15])=(0.0,0.0); 
        (D[14] *> O[16])=(0.0,0.0); 
        (D[14] *> O[17])=(0.0,0.0); 
        (D[14] *> O[18])=(0.0,0.0); 
        (D[14] *> O[19])=(0.0,0.0); 
        (D[14] *> O[20])=(0.0,0.0); 
        (D[14] *> O[21])=(0.0,0.0); 
        (D[14] *> O[22])=(0.0,0.0); 
        (D[14] *> O[23])=(0.0,0.0); 
        (D[14] *> O[24])=(0.0,0.0); 
        (D[14] *> O[25])=(0.0,0.0); 
        (D[14] *> O[26])=(0.0,0.0); 
        (D[14] *> O[27])=(0.0,0.0); 
        (D[14] *> O[28])=(0.0,0.0); 
        (D[14] *> O[29])=(0.0,0.0); 
        (D[14] *> O[30])=(0.0,0.0); 
        (D[14] *> O[31])=(0.0,0.0); 
        (D[15] *> O[0])=(0.0,0.0); 
        (D[15] *> O[1])=(0.0,0.0); 
        (D[15] *> O[2])=(0.0,0.0); 
        (D[15] *> O[3])=(0.0,0.0); 
        (D[15] *> O[4])=(0.0,0.0); 
        (D[15] *> O[5])=(0.0,0.0); 
        (D[15] *> O[6])=(0.0,0.0); 
        (D[15] *> O[7])=(0.0,0.0); 
        (D[15] *> O[8])=(0.0,0.0); 
        (D[15] *> O[9])=(0.0,0.0); 
        (D[15] *> O[10])=(0.0,0.0); 
        (D[15] *> O[11])=(0.0,0.0); 
        (D[15] *> O[12])=(0.0,0.0); 
        (D[15] *> O[13])=(0.0,0.0); 
        (D[15] *> O[14])=(0.0,0.0); 
        (D[15] *> O[15])=(0.0,0.0); 
        (D[15] *> O[16])=(0.0,0.0); 
        (D[15] *> O[17])=(0.0,0.0); 
        (D[15] *> O[18])=(0.0,0.0); 
        (D[15] *> O[19])=(0.0,0.0); 
        (D[15] *> O[20])=(0.0,0.0); 
        (D[15] *> O[21])=(0.0,0.0); 
        (D[15] *> O[22])=(0.0,0.0); 
        (D[15] *> O[23])=(0.0,0.0); 
        (D[15] *> O[24])=(0.0,0.0); 
        (D[15] *> O[25])=(0.0,0.0); 
        (D[15] *> O[26])=(0.0,0.0); 
        (D[15] *> O[27])=(0.0,0.0); 
        (D[15] *> O[28])=(0.0,0.0); 
        (D[15] *> O[29])=(0.0,0.0); 
        (D[15] *> O[30])=(0.0,0.0); 
        (D[15] *> O[31])=(0.0,0.0); 
        (IRSTBOT *> O[0])=(0.0,0.0); 
        (IRSTBOT *> O[1])=(0.0,0.0); 
        (IRSTBOT *> O[2])=(0.0,0.0); 
        (IRSTBOT *> O[3])=(0.0,0.0); 
        (IRSTBOT *> O[4])=(0.0,0.0); 
        (IRSTBOT *> O[5])=(0.0,0.0); 
        (IRSTBOT *> O[6])=(0.0,0.0); 
        (IRSTBOT *> O[7])=(0.0,0.0); 
        (IRSTBOT *> O[8])=(0.0,0.0); 
        (IRSTBOT *> O[9])=(0.0,0.0); 
        (IRSTBOT *> O[10])=(0.0,0.0); 
        (IRSTBOT *> O[11])=(0.0,0.0); 
        (IRSTBOT *> O[12])=(0.0,0.0); 
        (IRSTBOT *> O[13])=(0.0,0.0); 
        (IRSTBOT *> O[14])=(0.0,0.0); 
        (IRSTBOT *> O[15])=(0.0,0.0); 
        (IRSTBOT *> O[16])=(0.0,0.0); 
        (IRSTBOT *> O[17])=(0.0,0.0); 
        (IRSTBOT *> O[18])=(0.0,0.0); 
        (IRSTBOT *> O[19])=(0.0,0.0); 
        (IRSTBOT *> O[20])=(0.0,0.0); 
        (IRSTBOT *> O[21])=(0.0,0.0); 
        (IRSTBOT *> O[22])=(0.0,0.0); 
        (IRSTBOT *> O[23])=(0.0,0.0); 
        (IRSTBOT *> O[24])=(0.0,0.0); 
        (IRSTBOT *> O[25])=(0.0,0.0); 
        (IRSTBOT *> O[26])=(0.0,0.0); 
        (IRSTBOT *> O[27])=(0.0,0.0); 
        (IRSTBOT *> O[28])=(0.0,0.0); 
        (IRSTBOT *> O[29])=(0.0,0.0); 
        (IRSTBOT *> O[30])=(0.0,0.0); 
        (IRSTBOT *> O[31])=(0.0,0.0); 
        (ORSTBOT *> O[0])=(0.0,0.0); 
        (ORSTBOT *> O[1])=(0.0,0.0); 
        (ORSTBOT *> O[2])=(0.0,0.0); 
        (ORSTBOT *> O[3])=(0.0,0.0); 
        (ORSTBOT *> O[4])=(0.0,0.0); 
        (ORSTBOT *> O[5])=(0.0,0.0); 
        (ORSTBOT *> O[6])=(0.0,0.0); 
        (ORSTBOT *> O[7])=(0.0,0.0); 
        (ORSTBOT *> O[8])=(0.0,0.0); 
        (ORSTBOT *> O[9])=(0.0,0.0); 
        (ORSTBOT *> O[10])=(0.0,0.0); 
        (ORSTBOT *> O[11])=(0.0,0.0); 
        (ORSTBOT *> O[12])=(0.0,0.0); 
        (ORSTBOT *> O[13])=(0.0,0.0); 
        (ORSTBOT *> O[14])=(0.0,0.0); 
        (ORSTBOT *> O[15])=(0.0,0.0); 
        (ORSTBOT *> O[16])=(0.0,0.0); 
        (ORSTBOT *> O[17])=(0.0,0.0); 
        (ORSTBOT *> O[18])=(0.0,0.0); 
        (ORSTBOT *> O[19])=(0.0,0.0); 
        (ORSTBOT *> O[20])=(0.0,0.0); 
        (ORSTBOT *> O[21])=(0.0,0.0); 
        (ORSTBOT *> O[22])=(0.0,0.0); 
        (ORSTBOT *> O[23])=(0.0,0.0); 
        (ORSTBOT *> O[24])=(0.0,0.0); 
        (ORSTBOT *> O[25])=(0.0,0.0); 
        (ORSTBOT *> O[26])=(0.0,0.0); 
        (ORSTBOT *> O[27])=(0.0,0.0); 
        (ORSTBOT *> O[28])=(0.0,0.0); 
        (ORSTBOT *> O[29])=(0.0,0.0); 
        (ORSTBOT *> O[30])=(0.0,0.0); 
        (ORSTBOT *> O[31])=(0.0,0.0); 
        (ORSTTOP *> O[0])=(0.0,0.0); 
        (ORSTTOP *> O[1])=(0.0,0.0); 
        (ORSTTOP *> O[2])=(0.0,0.0); 
        (ORSTTOP *> O[3])=(0.0,0.0); 
        (ORSTTOP *> O[4])=(0.0,0.0); 
        (ORSTTOP *> O[5])=(0.0,0.0); 
        (ORSTTOP *> O[6])=(0.0,0.0); 
        (ORSTTOP *> O[7])=(0.0,0.0); 
        (ORSTTOP *> O[8])=(0.0,0.0); 
        (ORSTTOP *> O[9])=(0.0,0.0); 
        (ORSTTOP *> O[10])=(0.0,0.0); 
        (ORSTTOP *> O[11])=(0.0,0.0); 
        (ORSTTOP *> O[12])=(0.0,0.0); 
        (ORSTTOP *> O[13])=(0.0,0.0); 
        (ORSTTOP *> O[14])=(0.0,0.0); 
        (ORSTTOP *> O[15])=(0.0,0.0); 
        (ORSTTOP *> O[16])=(0.0,0.0); 
        (ORSTTOP *> O[17])=(0.0,0.0); 
        (ORSTTOP *> O[18])=(0.0,0.0); 
        (ORSTTOP *> O[19])=(0.0,0.0); 
        (ORSTTOP *> O[20])=(0.0,0.0); 
        (ORSTTOP *> O[21])=(0.0,0.0); 
        (ORSTTOP *> O[22])=(0.0,0.0); 
        (ORSTTOP *> O[23])=(0.0,0.0); 
        (ORSTTOP *> O[24])=(0.0,0.0); 
        (ORSTTOP *> O[25])=(0.0,0.0); 
        (ORSTTOP *> O[26])=(0.0,0.0); 
        (ORSTTOP *> O[27])=(0.0,0.0); 
        (ORSTTOP *> O[28])=(0.0,0.0); 
        (ORSTTOP *> O[29])=(0.0,0.0); 
        (ORSTTOP *> O[30])=(0.0,0.0); 
        (ORSTTOP *> O[31])=(0.0,0.0); 
        (OLOADTOP *> O[0])=(0.0,0.0); 
        (OLOADTOP *> O[1])=(0.0,0.0); 
        (OLOADTOP *> O[2])=(0.0,0.0); 
        (OLOADTOP *> O[3])=(0.0,0.0); 
        (OLOADTOP *> O[4])=(0.0,0.0); 
        (OLOADTOP *> O[5])=(0.0,0.0); 
        (OLOADTOP *> O[6])=(0.0,0.0); 
        (OLOADTOP *> O[7])=(0.0,0.0); 
        (OLOADTOP *> O[8])=(0.0,0.0); 
        (OLOADTOP *> O[9])=(0.0,0.0); 
        (OLOADTOP *> O[10])=(0.0,0.0); 
        (OLOADTOP *> O[11])=(0.0,0.0); 
        (OLOADTOP *> O[12])=(0.0,0.0); 
        (OLOADTOP *> O[13])=(0.0,0.0); 
        (OLOADTOP *> O[14])=(0.0,0.0); 
        (OLOADTOP *> O[15])=(0.0,0.0); 
        (OLOADTOP *> O[16])=(0.0,0.0); 
        (OLOADTOP *> O[17])=(0.0,0.0); 
        (OLOADTOP *> O[18])=(0.0,0.0); 
        (OLOADTOP *> O[19])=(0.0,0.0); 
        (OLOADTOP *> O[20])=(0.0,0.0); 
        (OLOADTOP *> O[21])=(0.0,0.0); 
        (OLOADTOP *> O[22])=(0.0,0.0); 
        (OLOADTOP *> O[23])=(0.0,0.0); 
        (OLOADTOP *> O[24])=(0.0,0.0); 
        (OLOADTOP *> O[25])=(0.0,0.0); 
        (OLOADTOP *> O[26])=(0.0,0.0); 
        (OLOADTOP *> O[27])=(0.0,0.0); 
        (OLOADTOP *> O[28])=(0.0,0.0); 
        (OLOADTOP *> O[29])=(0.0,0.0); 
        (OLOADTOP *> O[30])=(0.0,0.0); 
        (OLOADTOP *> O[31])=(0.0,0.0); 
        (OLOADBOT *> O[0])=(0.0,0.0); 
        (OLOADBOT *> O[1])=(0.0,0.0); 
        (OLOADBOT *> O[2])=(0.0,0.0); 
        (OLOADBOT *> O[3])=(0.0,0.0); 
        (OLOADBOT *> O[4])=(0.0,0.0); 
        (OLOADBOT *> O[5])=(0.0,0.0); 
        (OLOADBOT *> O[6])=(0.0,0.0); 
        (OLOADBOT *> O[7])=(0.0,0.0); 
        (OLOADBOT *> O[8])=(0.0,0.0); 
        (OLOADBOT *> O[9])=(0.0,0.0); 
        (OLOADBOT *> O[10])=(0.0,0.0); 
        (OLOADBOT *> O[11])=(0.0,0.0); 
        (OLOADBOT *> O[12])=(0.0,0.0); 
        (OLOADBOT *> O[13])=(0.0,0.0); 
        (OLOADBOT *> O[14])=(0.0,0.0); 
        (OLOADBOT *> O[15])=(0.0,0.0); 
        (OLOADBOT *> O[16])=(0.0,0.0); 
        (OLOADBOT *> O[17])=(0.0,0.0); 
        (OLOADBOT *> O[18])=(0.0,0.0); 
        (OLOADBOT *> O[19])=(0.0,0.0); 
        (OLOADBOT *> O[20])=(0.0,0.0); 
        (OLOADBOT *> O[21])=(0.0,0.0); 
        (OLOADBOT *> O[22])=(0.0,0.0); 
        (OLOADBOT *> O[23])=(0.0,0.0); 
        (OLOADBOT *> O[24])=(0.0,0.0); 
        (OLOADBOT *> O[25])=(0.0,0.0); 
        (OLOADBOT *> O[26])=(0.0,0.0); 
        (OLOADBOT *> O[27])=(0.0,0.0); 
        (OLOADBOT *> O[28])=(0.0,0.0); 
        (OLOADBOT *> O[29])=(0.0,0.0); 
        (OLOADBOT *> O[30])=(0.0,0.0); 
        (OLOADBOT *> O[31])=(0.0,0.0); 
      (OLOADTOP *> CO)=(0.0,0.0);
      (OLOADBOT *> CO)=(0.0,0.0);
      (OLOADTOP *> ACCUMCO)=(0.0,0.0);
      (OLOADBOT *> ACCUMCO)=(0.0,0.0);
        (ADDSUBTOP *> O[0])=(0.0,0.0); 
        (ADDSUBTOP *> O[1])=(0.0,0.0); 
        (ADDSUBTOP *> O[2])=(0.0,0.0); 
        (ADDSUBTOP *> O[3])=(0.0,0.0); 
        (ADDSUBTOP *> O[4])=(0.0,0.0); 
        (ADDSUBTOP *> O[5])=(0.0,0.0); 
        (ADDSUBTOP *> O[6])=(0.0,0.0); 
        (ADDSUBTOP *> O[7])=(0.0,0.0); 
        (ADDSUBTOP *> O[8])=(0.0,0.0); 
        (ADDSUBTOP *> O[9])=(0.0,0.0); 
        (ADDSUBTOP *> O[10])=(0.0,0.0); 
        (ADDSUBTOP *> O[11])=(0.0,0.0); 
        (ADDSUBTOP *> O[12])=(0.0,0.0); 
        (ADDSUBTOP *> O[13])=(0.0,0.0); 
        (ADDSUBTOP *> O[14])=(0.0,0.0); 
        (ADDSUBTOP *> O[15])=(0.0,0.0); 
        (ADDSUBTOP *> O[16])=(0.0,0.0); 
        (ADDSUBTOP *> O[17])=(0.0,0.0); 
        (ADDSUBTOP *> O[18])=(0.0,0.0); 
        (ADDSUBTOP *> O[19])=(0.0,0.0); 
        (ADDSUBTOP *> O[20])=(0.0,0.0); 
        (ADDSUBTOP *> O[21])=(0.0,0.0); 
        (ADDSUBTOP *> O[22])=(0.0,0.0); 
        (ADDSUBTOP *> O[23])=(0.0,0.0); 
        (ADDSUBTOP *> O[24])=(0.0,0.0); 
        (ADDSUBTOP *> O[25])=(0.0,0.0); 
        (ADDSUBTOP *> O[26])=(0.0,0.0); 
        (ADDSUBTOP *> O[27])=(0.0,0.0); 
        (ADDSUBTOP *> O[28])=(0.0,0.0); 
        (ADDSUBTOP *> O[29])=(0.0,0.0); 
        (ADDSUBTOP *> O[30])=(0.0,0.0); 
        (ADDSUBTOP *> O[31])=(0.0,0.0); 
        (ADDSUBBOT *> O[0])=(0.0,0.0); 
        (ADDSUBBOT *> O[1])=(0.0,0.0); 
        (ADDSUBBOT *> O[2])=(0.0,0.0); 
        (ADDSUBBOT *> O[3])=(0.0,0.0); 
        (ADDSUBBOT *> O[4])=(0.0,0.0); 
        (ADDSUBBOT *> O[5])=(0.0,0.0); 
        (ADDSUBBOT *> O[6])=(0.0,0.0); 
        (ADDSUBBOT *> O[7])=(0.0,0.0); 
        (ADDSUBBOT *> O[8])=(0.0,0.0); 
        (ADDSUBBOT *> O[9])=(0.0,0.0); 
        (ADDSUBBOT *> O[10])=(0.0,0.0); 
        (ADDSUBBOT *> O[11])=(0.0,0.0); 
        (ADDSUBBOT *> O[12])=(0.0,0.0); 
        (ADDSUBBOT *> O[13])=(0.0,0.0); 
        (ADDSUBBOT *> O[14])=(0.0,0.0); 
        (ADDSUBBOT *> O[15])=(0.0,0.0); 
        (ADDSUBBOT *> O[16])=(0.0,0.0); 
        (ADDSUBBOT *> O[17])=(0.0,0.0); 
        (ADDSUBBOT *> O[18])=(0.0,0.0); 
        (ADDSUBBOT *> O[19])=(0.0,0.0); 
        (ADDSUBBOT *> O[20])=(0.0,0.0); 
        (ADDSUBBOT *> O[21])=(0.0,0.0); 
        (ADDSUBBOT *> O[22])=(0.0,0.0); 
        (ADDSUBBOT *> O[23])=(0.0,0.0); 
        (ADDSUBBOT *> O[24])=(0.0,0.0); 
        (ADDSUBBOT *> O[25])=(0.0,0.0); 
        (ADDSUBBOT *> O[26])=(0.0,0.0); 
        (ADDSUBBOT *> O[27])=(0.0,0.0); 
        (ADDSUBBOT *> O[28])=(0.0,0.0); 
        (ADDSUBBOT *> O[29])=(0.0,0.0); 
        (ADDSUBBOT *> O[30])=(0.0,0.0); 
        (ADDSUBBOT *> O[31])=(0.0,0.0); 
      (ADDSUBTOP *> CO)=(0.0,0.0);
      (ADDSUBBOT *> CO)=(0.0,0.0);
      (ADDSUBTOP *> ACCUMCO)=(0.0,0.0);
      (ADDSUBBOT *> ACCUMCO)=(0.0,0.0);
        (CLK *> O[0])=(0.0,0.0); 
        (CLK *> O[1])=(0.0,0.0); 
        (CLK *> O[2])=(0.0,0.0); 
        (CLK *> O[3])=(0.0,0.0); 
        (CLK *> O[4])=(0.0,0.0); 
        (CLK *> O[5])=(0.0,0.0); 
        (CLK *> O[6])=(0.0,0.0); 
        (CLK *> O[7])=(0.0,0.0); 
        (CLK *> O[8])=(0.0,0.0); 
        (CLK *> O[9])=(0.0,0.0); 
        (CLK *> O[10])=(0.0,0.0); 
        (CLK *> O[11])=(0.0,0.0); 
        (CLK *> O[12])=(0.0,0.0); 
        (CLK *> O[13])=(0.0,0.0); 
        (CLK *> O[14])=(0.0,0.0); 
        (CLK *> O[15])=(0.0,0.0); 
        (CLK *> O[16])=(0.0,0.0); 
        (CLK *> O[17])=(0.0,0.0); 
        (CLK *> O[18])=(0.0,0.0); 
        (CLK *> O[19])=(0.0,0.0); 
        (CLK *> O[20])=(0.0,0.0); 
        (CLK *> O[21])=(0.0,0.0); 
        (CLK *> O[22])=(0.0,0.0); 
        (CLK *> O[23])=(0.0,0.0); 
        (CLK *> O[24])=(0.0,0.0); 
        (CLK *> O[25])=(0.0,0.0); 
        (CLK *> O[26])=(0.0,0.0); 
        (CLK *> O[27])=(0.0,0.0); 
        (CLK *> O[28])=(0.0,0.0); 
        (CLK *> O[29])=(0.0,0.0); 
        (CLK *> O[30])=(0.0,0.0); 
        (CLK *> O[31])=(0.0,0.0); 
      (CLK *> O)=(0.0,0.0);
      (CLK *> ACCUMCO)=(0.0,0.0);
        (ACCUMCI *> O[0])=(0.0,0.0); 
        (ACCUMCI *> O[1])=(0.0,0.0); 
        (ACCUMCI *> O[2])=(0.0,0.0); 
        (ACCUMCI *> O[3])=(0.0,0.0); 
        (ACCUMCI *> O[4])=(0.0,0.0); 
        (ACCUMCI *> O[5])=(0.0,0.0); 
        (ACCUMCI *> O[6])=(0.0,0.0); 
        (ACCUMCI *> O[7])=(0.0,0.0); 
        (ACCUMCI *> O[8])=(0.0,0.0); 
        (ACCUMCI *> O[9])=(0.0,0.0); 
        (ACCUMCI *> O[10])=(0.0,0.0); 
        (ACCUMCI *> O[11])=(0.0,0.0); 
        (ACCUMCI *> O[12])=(0.0,0.0); 
        (ACCUMCI *> O[13])=(0.0,0.0); 
        (ACCUMCI *> O[14])=(0.0,0.0); 
        (ACCUMCI *> O[15])=(0.0,0.0); 
        (ACCUMCI *> O[16])=(0.0,0.0); 
        (ACCUMCI *> O[17])=(0.0,0.0); 
        (ACCUMCI *> O[18])=(0.0,0.0); 
        (ACCUMCI *> O[19])=(0.0,0.0); 
        (ACCUMCI *> O[20])=(0.0,0.0); 
        (ACCUMCI *> O[21])=(0.0,0.0); 
        (ACCUMCI *> O[22])=(0.0,0.0); 
        (ACCUMCI *> O[23])=(0.0,0.0); 
        (ACCUMCI *> O[24])=(0.0,0.0); 
        (ACCUMCI *> O[25])=(0.0,0.0); 
        (ACCUMCI *> O[26])=(0.0,0.0); 
        (ACCUMCI *> O[27])=(0.0,0.0); 
        (ACCUMCI *> O[28])=(0.0,0.0); 
        (ACCUMCI *> O[29])=(0.0,0.0); 
        (ACCUMCI *> O[30])=(0.0,0.0); 
        (ACCUMCI *> O[31])=(0.0,0.0); 
        (ACCUMCI *> O[0])=(0.0,0.0); 
        (ACCUMCI *> O[1])=(0.0,0.0); 
        (ACCUMCI *> O[2])=(0.0,0.0); 
        (ACCUMCI *> O[3])=(0.0,0.0); 
        (ACCUMCI *> O[4])=(0.0,0.0); 
        (ACCUMCI *> O[5])=(0.0,0.0); 
        (ACCUMCI *> O[6])=(0.0,0.0); 
        (ACCUMCI *> O[7])=(0.0,0.0); 
        (ACCUMCI *> O[8])=(0.0,0.0); 
        (ACCUMCI *> O[9])=(0.0,0.0); 
        (ACCUMCI *> O[10])=(0.0,0.0); 
        (ACCUMCI *> O[11])=(0.0,0.0); 
        (ACCUMCI *> O[12])=(0.0,0.0); 
        (ACCUMCI *> O[13])=(0.0,0.0); 
        (ACCUMCI *> O[14])=(0.0,0.0); 
        (ACCUMCI *> O[15])=(0.0,0.0); 
        (ACCUMCI *> O[16])=(0.0,0.0); 
        (ACCUMCI *> O[17])=(0.0,0.0); 
        (ACCUMCI *> O[18])=(0.0,0.0); 
        (ACCUMCI *> O[19])=(0.0,0.0); 
        (ACCUMCI *> O[20])=(0.0,0.0); 
        (ACCUMCI *> O[21])=(0.0,0.0); 
        (ACCUMCI *> O[22])=(0.0,0.0); 
        (ACCUMCI *> O[23])=(0.0,0.0); 
        (ACCUMCI *> O[24])=(0.0,0.0); 
        (ACCUMCI *> O[25])=(0.0,0.0); 
        (ACCUMCI *> O[26])=(0.0,0.0); 
        (ACCUMCI *> O[27])=(0.0,0.0); 
        (ACCUMCI *> O[28])=(0.0,0.0); 
        (ACCUMCI *> O[29])=(0.0,0.0); 
        (ACCUMCI *> O[30])=(0.0,0.0); 
        (ACCUMCI *> O[31])=(0.0,0.0); 
      (ACCUMCI *> CO)=(0.0,0.0);
      (ACCUMCI *> ACCUMCO)=(0.0,0.0);
        (CI *> O[0])=(0.0,0.0); 
        (CI *> O[1])=(0.0,0.0); 
        (CI *> O[2])=(0.0,0.0); 
        (CI *> O[3])=(0.0,0.0); 
        (CI *> O[4])=(0.0,0.0); 
        (CI *> O[5])=(0.0,0.0); 
        (CI *> O[6])=(0.0,0.0); 
        (CI *> O[7])=(0.0,0.0); 
        (CI *> O[8])=(0.0,0.0); 
        (CI *> O[9])=(0.0,0.0); 
        (CI *> O[10])=(0.0,0.0); 
        (CI *> O[11])=(0.0,0.0); 
        (CI *> O[12])=(0.0,0.0); 
        (CI *> O[13])=(0.0,0.0); 
        (CI *> O[14])=(0.0,0.0); 
        (CI *> O[15])=(0.0,0.0); 
        (CI *> O[16])=(0.0,0.0); 
        (CI *> O[17])=(0.0,0.0); 
        (CI *> O[18])=(0.0,0.0); 
        (CI *> O[19])=(0.0,0.0); 
        (CI *> O[20])=(0.0,0.0); 
        (CI *> O[21])=(0.0,0.0); 
        (CI *> O[22])=(0.0,0.0); 
        (CI *> O[23])=(0.0,0.0); 
        (CI *> O[24])=(0.0,0.0); 
        (CI *> O[25])=(0.0,0.0); 
        (CI *> O[26])=(0.0,0.0); 
        (CI *> O[27])=(0.0,0.0); 
        (CI *> O[28])=(0.0,0.0); 
        (CI *> O[29])=(0.0,0.0); 
        (CI *> O[30])=(0.0,0.0); 
        (CI *> O[31])=(0.0,0.0); 
      (CI *> CO)=(0.0,0.0);
      (CI *> ACCUMCO)=(0.0,0.0);
      (CLK *> SIGNEXTOUT)=(0.0,0.0);
        (A[0] *> CO)=(0.0,0.0); 
        (A[1] *> CO)=(0.0,0.0); 
        (A[2] *> CO)=(0.0,0.0); 
        (A[3] *> CO)=(0.0,0.0); 
        (A[4] *> CO)=(0.0,0.0); 
        (A[5] *> CO)=(0.0,0.0); 
        (A[6] *> CO)=(0.0,0.0); 
        (A[7] *> CO)=(0.0,0.0); 
        (A[8] *> CO)=(0.0,0.0); 
        (A[9] *> CO)=(0.0,0.0); 
        (A[10] *> CO)=(0.0,0.0); 
        (A[11] *> CO)=(0.0,0.0); 
        (A[12] *> CO)=(0.0,0.0); 
        (A[13] *> CO)=(0.0,0.0); 
        (A[14] *> CO)=(0.0,0.0); 
        (A[15] *> CO)=(0.0,0.0); 
        (A[0] *> ACCUMCO)=(0.0,0.0); 
        (A[1] *> ACCUMCO)=(0.0,0.0); 
        (A[2] *> ACCUMCO)=(0.0,0.0); 
        (A[3] *> ACCUMCO)=(0.0,0.0); 
        (A[4] *> ACCUMCO)=(0.0,0.0); 
        (A[5] *> ACCUMCO)=(0.0,0.0); 
        (A[6] *> ACCUMCO)=(0.0,0.0); 
        (A[7] *> ACCUMCO)=(0.0,0.0); 
        (A[8] *> ACCUMCO)=(0.0,0.0); 
        (A[9] *> ACCUMCO)=(0.0,0.0); 
        (A[10] *> ACCUMCO)=(0.0,0.0); 
        (A[11] *> ACCUMCO)=(0.0,0.0); 
        (A[12] *> ACCUMCO)=(0.0,0.0); 
        (A[13] *> ACCUMCO)=(0.0,0.0); 
        (A[14] *> ACCUMCO)=(0.0,0.0); 
        (A[15] *> ACCUMCO)=(0.0,0.0); 
        (A[0] *> SIGNEXTOUT)=(0.0,0.0); 
        (A[1] *> SIGNEXTOUT)=(0.0,0.0); 
        (A[2] *> SIGNEXTOUT)=(0.0,0.0); 
        (A[3] *> SIGNEXTOUT)=(0.0,0.0); 
        (A[4] *> SIGNEXTOUT)=(0.0,0.0); 
        (A[5] *> SIGNEXTOUT)=(0.0,0.0); 
        (A[6] *> SIGNEXTOUT)=(0.0,0.0); 
        (A[7] *> SIGNEXTOUT)=(0.0,0.0); 
        (A[8] *> SIGNEXTOUT)=(0.0,0.0); 
        (A[9] *> SIGNEXTOUT)=(0.0,0.0); 
        (A[10] *> SIGNEXTOUT)=(0.0,0.0); 
        (A[11] *> SIGNEXTOUT)=(0.0,0.0); 
        (A[12] *> SIGNEXTOUT)=(0.0,0.0); 
        (A[13] *> SIGNEXTOUT)=(0.0,0.0); 
        (A[14] *> SIGNEXTOUT)=(0.0,0.0); 
        (A[15] *> SIGNEXTOUT)=(0.0,0.0); 
        (D[0] *> CO)=(0.0,0.0); 
        (D[1] *> CO)=(0.0,0.0); 
        (D[2] *> CO)=(0.0,0.0); 
        (D[3] *> CO)=(0.0,0.0); 
        (D[4] *> CO)=(0.0,0.0); 
        (D[5] *> CO)=(0.0,0.0); 
        (D[6] *> CO)=(0.0,0.0); 
        (D[7] *> CO)=(0.0,0.0); 
        (D[8] *> CO)=(0.0,0.0); 
        (D[9] *> CO)=(0.0,0.0); 
        (D[10] *> CO)=(0.0,0.0); 
        (D[11] *> CO)=(0.0,0.0); 
        (D[12] *> CO)=(0.0,0.0); 
        (D[13] *> CO)=(0.0,0.0); 
        (D[14] *> CO)=(0.0,0.0); 
        (D[15] *> CO)=(0.0,0.0); 
        (D[0] *> ACCUMCO)=(0.0,0.0); 
        (D[1] *> ACCUMCO)=(0.0,0.0); 
        (D[2] *> ACCUMCO)=(0.0,0.0); 
        (D[3] *> ACCUMCO)=(0.0,0.0); 
        (D[4] *> ACCUMCO)=(0.0,0.0); 
        (D[5] *> ACCUMCO)=(0.0,0.0); 
        (D[6] *> ACCUMCO)=(0.0,0.0); 
        (D[7] *> ACCUMCO)=(0.0,0.0); 
        (D[8] *> ACCUMCO)=(0.0,0.0); 
        (D[9] *> ACCUMCO)=(0.0,0.0); 
        (D[10] *> ACCUMCO)=(0.0,0.0); 
        (D[11] *> ACCUMCO)=(0.0,0.0); 
        (D[12] *> ACCUMCO)=(0.0,0.0); 
        (D[13] *> ACCUMCO)=(0.0,0.0); 
        (D[14] *> ACCUMCO)=(0.0,0.0); 
        (D[15] *> ACCUMCO)=(0.0,0.0); 
        (D[0] *> SIGNEXTOUT)=(0.0,0.0); 
        (D[1] *> SIGNEXTOUT)=(0.0,0.0); 
        (D[2] *> SIGNEXTOUT)=(0.0,0.0); 
        (D[3] *> SIGNEXTOUT)=(0.0,0.0); 
        (D[4] *> SIGNEXTOUT)=(0.0,0.0); 
        (D[5] *> SIGNEXTOUT)=(0.0,0.0); 
        (D[6] *> SIGNEXTOUT)=(0.0,0.0); 
        (D[7] *> SIGNEXTOUT)=(0.0,0.0); 
        (D[8] *> SIGNEXTOUT)=(0.0,0.0); 
        (D[9] *> SIGNEXTOUT)=(0.0,0.0); 
        (D[10] *> SIGNEXTOUT)=(0.0,0.0); 
        (D[11] *> SIGNEXTOUT)=(0.0,0.0); 
        (D[12] *> SIGNEXTOUT)=(0.0,0.0); 
        (D[13] *> SIGNEXTOUT)=(0.0,0.0); 
        (D[14] *> SIGNEXTOUT)=(0.0,0.0); 
        (D[15] *> SIGNEXTOUT)=(0.0,0.0); 
        (C[0] *> CO)=(0.0,0.0); 
        (C[1] *> CO)=(0.0,0.0); 
        (C[2] *> CO)=(0.0,0.0); 
        (C[3] *> CO)=(0.0,0.0); 
        (C[4] *> CO)=(0.0,0.0); 
        (C[5] *> CO)=(0.0,0.0); 
        (C[6] *> CO)=(0.0,0.0); 
        (C[7] *> CO)=(0.0,0.0); 
        (C[8] *> CO)=(0.0,0.0); 
        (C[9] *> CO)=(0.0,0.0); 
        (C[10] *> CO)=(0.0,0.0); 
        (C[11] *> CO)=(0.0,0.0); 
        (C[12] *> CO)=(0.0,0.0); 
        (C[13] *> CO)=(0.0,0.0); 
        (C[14] *> CO)=(0.0,0.0); 
        (C[15] *> CO)=(0.0,0.0); 
        (C[0] *> ACCUMCO)=(0.0,0.0); 
        (C[1] *> ACCUMCO)=(0.0,0.0); 
        (C[2] *> ACCUMCO)=(0.0,0.0); 
        (C[3] *> ACCUMCO)=(0.0,0.0); 
        (C[4] *> ACCUMCO)=(0.0,0.0); 
        (C[5] *> ACCUMCO)=(0.0,0.0); 
        (C[6] *> ACCUMCO)=(0.0,0.0); 
        (C[7] *> ACCUMCO)=(0.0,0.0); 
        (C[8] *> ACCUMCO)=(0.0,0.0); 
        (C[9] *> ACCUMCO)=(0.0,0.0); 
        (C[10] *> ACCUMCO)=(0.0,0.0); 
        (C[11] *> ACCUMCO)=(0.0,0.0); 
        (C[12] *> ACCUMCO)=(0.0,0.0); 
        (C[13] *> ACCUMCO)=(0.0,0.0); 
        (C[14] *> ACCUMCO)=(0.0,0.0); 
        (C[15] *> ACCUMCO)=(0.0,0.0); 
        (C[0] *> SIGNEXTOUT)=(0.0,0.0); 
        (C[1] *> SIGNEXTOUT)=(0.0,0.0); 
        (C[2] *> SIGNEXTOUT)=(0.0,0.0); 
        (C[3] *> SIGNEXTOUT)=(0.0,0.0); 
        (C[4] *> SIGNEXTOUT)=(0.0,0.0); 
        (C[5] *> SIGNEXTOUT)=(0.0,0.0); 
        (C[6] *> SIGNEXTOUT)=(0.0,0.0); 
        (C[7] *> SIGNEXTOUT)=(0.0,0.0); 
        (C[8] *> SIGNEXTOUT)=(0.0,0.0); 
        (C[9] *> SIGNEXTOUT)=(0.0,0.0); 
        (C[10] *> SIGNEXTOUT)=(0.0,0.0); 
        (C[11] *> SIGNEXTOUT)=(0.0,0.0); 
        (C[12] *> SIGNEXTOUT)=(0.0,0.0); 
        (C[13] *> SIGNEXTOUT)=(0.0,0.0); 
        (C[14] *> SIGNEXTOUT)=(0.0,0.0); 
        (C[15] *> SIGNEXTOUT)=(0.0,0.0); 
        (B[0] *> CO)=(0.0,0.0); 
        (B[1] *> CO)=(0.0,0.0); 
        (B[2] *> CO)=(0.0,0.0); 
        (B[3] *> CO)=(0.0,0.0); 
        (B[4] *> CO)=(0.0,0.0); 
        (B[5] *> CO)=(0.0,0.0); 
        (B[6] *> CO)=(0.0,0.0); 
        (B[7] *> CO)=(0.0,0.0); 
        (B[8] *> CO)=(0.0,0.0); 
        (B[9] *> CO)=(0.0,0.0); 
        (B[10] *> CO)=(0.0,0.0); 
        (B[11] *> CO)=(0.0,0.0); 
        (B[12] *> CO)=(0.0,0.0); 
        (B[13] *> CO)=(0.0,0.0); 
        (B[14] *> CO)=(0.0,0.0); 
        (B[15] *> CO)=(0.0,0.0); 
        (B[0] *> ACCUMCO)=(0.0,0.0); 
        (B[1] *> ACCUMCO)=(0.0,0.0); 
        (B[2] *> ACCUMCO)=(0.0,0.0); 
        (B[3] *> ACCUMCO)=(0.0,0.0); 
        (B[4] *> ACCUMCO)=(0.0,0.0); 
        (B[5] *> ACCUMCO)=(0.0,0.0); 
        (B[6] *> ACCUMCO)=(0.0,0.0); 
        (B[7] *> ACCUMCO)=(0.0,0.0); 
        (B[8] *> ACCUMCO)=(0.0,0.0); 
        (B[9] *> ACCUMCO)=(0.0,0.0); 
        (B[10] *> ACCUMCO)=(0.0,0.0); 
        (B[11] *> ACCUMCO)=(0.0,0.0); 
        (B[12] *> ACCUMCO)=(0.0,0.0); 
        (B[13] *> ACCUMCO)=(0.0,0.0); 
        (B[14] *> ACCUMCO)=(0.0,0.0); 
        (B[15] *> ACCUMCO)=(0.0,0.0); 
        (B[0] *> SIGNEXTOUT)=(0.0,0.0); 
        (B[1] *> SIGNEXTOUT)=(0.0,0.0); 
        (B[2] *> SIGNEXTOUT)=(0.0,0.0); 
        (B[3] *> SIGNEXTOUT)=(0.0,0.0); 
        (B[4] *> SIGNEXTOUT)=(0.0,0.0); 
        (B[5] *> SIGNEXTOUT)=(0.0,0.0); 
        (B[6] *> SIGNEXTOUT)=(0.0,0.0); 
        (B[7] *> SIGNEXTOUT)=(0.0,0.0); 
        (B[8] *> SIGNEXTOUT)=(0.0,0.0); 
        (B[9] *> SIGNEXTOUT)=(0.0,0.0); 
        (B[10] *> SIGNEXTOUT)=(0.0,0.0); 
        (B[11] *> SIGNEXTOUT)=(0.0,0.0); 
        (B[12] *> SIGNEXTOUT)=(0.0,0.0); 
        (B[13] *> SIGNEXTOUT)=(0.0,0.0); 
        (B[14] *> SIGNEXTOUT)=(0.0,0.0); 
        (B[15] *> SIGNEXTOUT)=(0.0,0.0); 
		(CLK *> CO)=(0.0,0.0); 
	 
		  $recovery( posedge IRSTTOP,posedge CLK , 1.0);
		  $recovery( negedge IRSTTOP, posedge CLK ,1.0);   
		  $removal( posedge IRSTTOP, posedge CLK ,1.0);
		  $removal( negedge IRSTTOP, posedge CLK ,1.0);
		  $recovery(posedge IRSTBOT , posedge CLK ,1.0);
		  $recovery(negedge IRSTBOT , posedge CLK ,1.0);	 
		  $removal(posedge IRSTBOT , posedge CLK ,1.0);
		  $removal(negedge IRSTBOT , posedge CLK ,1.0);
		  $recovery( posedge ORSTTOP, posedge CLK ,1.0);
		  $recovery( negedge ORSTTOP, posedge CLK ,1.0);
		  $removal( posedge ORSTTOP, posedge CLK ,1.0);
		  $removal( negedge ORSTTOP, posedge CLK ,1.0);
		  $recovery(posedge ORSTBOT , posedge CLK ,1.0);
		  $recovery(negedge ORSTBOT , posedge CLK ,1.0);	   
		  $removal(posedge ORSTBOT , posedge CLK ,1.0);
		  $removal(negedge ORSTBOT , posedge CLK ,1.0);
		  $width (posedge CLK, 1.0 ); 
		  $period (posedge CLK, 1.0 ); 

		  $setuphold( posedge CLK,posedge A[0],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge A[0],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge A[1],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge A[1],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge A[2],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge A[2],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge A[3],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge A[3],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge A[4],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge A[4],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge A[5],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge A[5],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge A[6],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge A[6],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge A[7],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge A[7],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge A[8],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge A[8],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge A[9],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge A[9],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge A[10],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge A[10],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge A[11],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge A[11],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge A[12],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge A[12],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge A[13],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge A[13],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge A[14],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge A[14],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge A[15],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge A[15],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge B[0],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge B[0],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge B[1],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge B[1],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge B[2],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge B[2],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge B[3],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge B[3],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge B[4],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge B[4],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge B[5],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge B[5],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge B[6],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge B[6],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge B[7],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge B[7],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge B[8],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge B[8],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge B[9],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge B[9],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge B[10],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge B[10],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge B[11],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge B[11],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge B[12],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge B[12],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge B[13],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge B[13],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge B[14],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge B[14],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge B[15],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge B[15],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge C[0],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge C[0],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge C[1],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge C[1],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge C[2],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge C[2],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge C[3],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge C[3],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge C[4],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge C[4],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge C[5],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge C[5],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge C[6],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge C[6],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge C[7],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge C[7],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge C[8],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge C[8],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge C[9],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge C[9],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge C[10],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge C[10],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge C[11],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge C[11],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge C[12],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge C[12],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge C[13],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge C[13],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge C[14],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge C[14],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge C[15],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge C[15],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge D[0],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge D[0],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge D[1],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge D[1],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge D[2],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge D[2],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge D[3],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge D[3],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge D[4],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge D[4],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge D[5],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge D[5],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge D[6],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge D[6],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge D[7],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge D[7],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge D[8],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge D[8],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge D[9],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge D[9],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge D[10],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge D[10],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge D[11],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge D[11],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge D[12],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge D[12],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge D[13],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge D[13],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge D[14],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge D[14],1.0, 1.0, NOTIFIER);
       $setuphold( posedge CLK,posedge D[15],1.0,1.0, NOTIFIER);
       $setuphold(posedge CLK,negedge D[15],1.0, 1.0, NOTIFIER);
		  
		  
		  
		
		   $setuphold(posedge CLK, posedge AHOLD, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, posedge BHOLD, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, posedge CHOLD, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, posedge DHOLD, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, posedge ADDSUBTOP, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, posedge OHOLDTOP, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, posedge ADDSUBBOT, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, posedge OHOLDBOT, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, posedge OLOADTOP, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, posedge OLOADBOT, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, posedge CI, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, posedge ACCUMCI, 1.0, 1.0, NOTIFIER);	 
		   
		  
		   $setuphold(posedge CLK, negedge AHOLD, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, negedge BHOLD, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, negedge CHOLD, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, negedge DHOLD, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, negedge ADDSUBTOP, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, negedge OHOLDTOP, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, negedge ADDSUBBOT, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, negedge OHOLDBOT, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, negedge OLOADTOP, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, negedge OLOADBOT, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, negedge CI, 1.0, 1.0, NOTIFIER);
		   $setuphold(posedge CLK, negedge ACCUMCI, 1.0, 1.0, NOTIFIER);
 
		 
		 
		 
		 endspecify
`endif		   
		

endmodule

//////////////////////////////////////////////////////////////////////////////////
// mac16_physical
//////////////////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps

module mac16_physical  (
	 CLK ,
	 IHRST,
	 ILRST,
	 OHRST,
	 OLRST,
	 
	 A ,
	 B ,
	 C ,
	 D ,
	 
	 CBIT,
	 
	 AHLD,
	 BHLD,
	 CHLD,
	 DHLD,
	 OHHLD,
	 OLHLD,

 
	 OHADS,
	 OLADS,
	 OHLDA,
	 OLLDA,
	 
	 CICAS,
	 CI,
	 SIGNEXTIN,
	 SIGNEXTOUT,

	 COCAS,
	 CO,
	 O
    );

	 input CLK ;
	 input IHRST;
	 input ILRST;
	 input OHRST;
	 input OLRST;
	 
	 input [15:0] A ;
	 input [15:0] B ;
	 input [15:0] C ;
	 input [15:0] D ;
	 
	 input [24:0] CBIT;
	 
	 input AHLD;
	 input BHLD;
	 input CHLD;
	 input DHLD;
	 input OHHLD;
	 input OLHLD;

 
	 input OHADS;
	 input OLADS;
	 input OHLDA;
	 input OLLDA;
	 
	 input CICAS;
	 input CI;
	 input SIGNEXTIN;
	 output SIGNEXTOUT;
	 
	 output COCAS;
	 output CO;
	 output [31:0] O;
	
	
wire AENA, BENA, CENA, DENA, OHENA, OLENA;
assign AENA = ~AHLD;
assign BENA = ~BHLD;
assign CENA = ~CHLD;
assign DENA = ~DHLD;

assign OHENA = ~OHHLD;
assign OLENA = ~OLHLD;


wire ASEL, BSEL, CSEL, DSEL, FSEL, JKSEL, GSEL, HSEL;
wire OHADDA_SEL, OLADDA_SEL, MPY_8X8_MODE, ASGND, BSGND;
wire [1:0] OHOMUX_SEL, OLOMUX_SEL, OHADDB_SEL, OLADDB_SEL, OHCARRYMUX_SEL, OLCARRYMUX_SEL;

assign ASEL = CBIT[1];
assign BSEL = CBIT[2];
assign CSEL = CBIT[0];
assign DSEL = CBIT[3];

assign FSEL = CBIT[4];
assign JKSEL = CBIT[6];
assign GSEL = CBIT[5];
assign HSEL = CBIT[7];

assign OHOMUX_SEL[1:0] = CBIT[9:8];	
assign OLOMUX_SEL[1:0] = CBIT[16:15];	
assign OHADDA_SEL = CBIT[12];
assign OLADDA_SEL = CBIT[19];
assign OHADDB_SEL[1:0] = CBIT[11:10];	
assign OLADDB_SEL[1:0] = CBIT[18:17];	
assign OHCARRYMUX_SEL[1:0] = CBIT[14:13];
assign OLCARRYMUX_SEL[1:0] = CBIT[21:20];
assign MPY_8X8_MODE = CBIT[22];
assign ASGND = CBIT[23];
assign BSGND = CBIT[24];

wire [15:0] REG_A ;
wire [15:0] REG_B ;
wire [15:0] REG_C ;
wire [15:0] REG_D ;

wire [15:0] OH_8X8;
wire [15:0] OL_8X8;
wire [31:0] O_16X16;

wire MAC16_SIGNOUT_L, MAC16_SIGNOUT_H;

assign SIGNEXTOUT = MAC16_SIGNOUT_H;

REG_BYPASS_MUX  A_REG (
	.D(A) ,
	.Q(REG_A) ,
	.ENA(AENA) ,
	.CLK(CLK) ,
	.RST(IHRST) ,
	.SELM(ASEL) 
); 

REG_BYPASS_MUX  B_REG (
	.D(B) ,
	.Q(REG_B) ,
	.ENA(BENA) ,
	.CLK(CLK) ,
	.RST(ILRST) ,
	.SELM(BSEL) 
); 

REG_BYPASS_MUX  C_REG (
	.D(C) ,
	.Q(REG_C) ,
	.ENA(CENA) ,
	.CLK(CLK) ,
	.RST(IHRST) ,
	.SELM(CSEL) 
); 

REG_BYPASS_MUX  D_REG (
	.D(D) ,
	.Q(REG_D) ,
	.ENA(DENA) ,
	.CLK(CLK) ,
	.RST(ILRST) ,
	.SELM(DSEL) 
); 

MULT_ACCUM HI_MAC (
	.DIRECT_INPUT(REG_C),
	.MULT_INPUT(REG_A),
	.MULT_8x8(OH_8X8[15:0]),
	.MULT_16x16(O_16X16[31:16]),
	.ADDSUB(OHADS),
	.CLK(CLK),
	.CICAS(COCAS_L),
	.CI(CO_L),
	.SIGNEXTIN(MAC16_SIGNOUT_L) ,
	.SIGNEXTOUT(MAC16_SIGNOUT_H) ,
	.LDA(OHLDA),
	.RST(OHRST),
	.ENA(OHENA),
	.COCAS(COCAS),
	.CO(CO),
	.O(O[31:16]),
	.OUTMUX_SEL(OHOMUX_SEL[1:0]),
	.ADDER_A_IN_SEL(OHADDA_SEL),
	.ADDER_B_IN_SEL(OHADDB_SEL[1:0]),
	.CARRYMUX_SEL(OHCARRYMUX_SEL[1:0])
    );

MULT_ACCUM LO_MAC (
	.DIRECT_INPUT(REG_D),
	.MULT_INPUT(REG_B),
	.MULT_8x8(OL_8X8[15:0]),
	.MULT_16x16(O_16X16[15:0]),
	.ADDSUB(OLADS),
	.CLK(CLK),
	.CICAS(CICAS),
	.CI(CI),
	.SIGNEXTIN(SIGNEXTIN) ,
	.SIGNEXTOUT(MAC16_SIGNOUT_L) ,
	.LDA(OLLDA),
	.RST(OLRST),
	.ENA(OLENA),
	.COCAS(COCAS_L),
	.CO(CO_L),
	.O(O[15:0]),
	.OUTMUX_SEL(OLOMUX_SEL[1:0]),
	.ADDER_A_IN_SEL(OLADDA_SEL),
	.ADDER_B_IN_SEL(OLADDB_SEL[1:0]),
	.CARRYMUX_SEL(OLCARRYMUX_SEL[1:0])
    );
	 
MPY16X16 MULTIPLER (
	.clk(CLK),
	.IHRST(IHRST),
	.ILRST(ILRST),
	.FSEL(FSEL),
	.GSEL(GSEL),
	.HSEL(HSEL),
	.JKSEL(JKSEL),
	.MPY_8X8_MODE(MPY_8X8_MODE),
	.ASGND(ASGND),
	.BSGND(BSGND),
	.A(REG_A[15:0]),
	.B(REG_B[15:0]),
	.OH_8X8(OH_8X8[15:0]),
	.OL_8X8(OL_8X8[15:0]),
	.O_16X16(O_16X16[31:0])
);

endmodule



//////////////////////////////////////////////////////////////////////////////////
// Module Name:    MPY16X16
//////////////////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps

//////////////////////////////////////////////////// 
`define  SIGNED_DATA		1'b1
`define  UNSIGNED_DATA		1'b0
////////////////////////////////////////////////////

module booth_encoder(booth_single, booth_double, booth_negtive, multiplier, signed_mpy);
input	[7:0]multiplier;
output	[4:0]booth_single;
output	[4:0]booth_double;
output	[4:0]booth_negtive;
input	signed_mpy;

wire	[10:0]booth_in;
wire	[1:0]sign_ext;
assign sign_ext=(signed_mpy==1'b1)?{2{multiplier[7]}} : 2'b00;

assign booth_in={sign_ext ,multiplier[7:0],1'b0};


assign  booth_negtive[0]=booth_in[2];
assign  booth_negtive[1]=booth_in[4];
assign  booth_negtive[2]=booth_in[6];
assign  booth_negtive[3]=booth_in[8];
assign  booth_negtive[4]=booth_in[10];

assign  booth_single[0]=booth_in[0]^booth_in[1];
assign  booth_single[1]=booth_in[2]^booth_in[3];
assign  booth_single[2]=booth_in[4]^booth_in[5];
assign  booth_single[3]=booth_in[6]^booth_in[7];
assign  booth_single[4]=booth_in[8]^booth_in[9];


assign  booth_double[0]=~(~(booth_in[0] & booth_in[1] & ~booth_in[2]) & ~(~booth_in[0] & ~booth_in[1] & booth_in[2]));
assign  booth_double[1]=~(~(booth_in[2] & booth_in[3] & ~booth_in[4]) & ~(~booth_in[2] & ~booth_in[3] & booth_in[4]));
assign  booth_double[2]=~(~(booth_in[4] & booth_in[5] & ~booth_in[6]) & ~(~booth_in[4] & ~booth_in[5] & booth_in[6]));
assign  booth_double[3]=~(~(booth_in[6] & booth_in[7] & ~booth_in[8]) & ~(~booth_in[6] & ~booth_in[7] & booth_in[8]));
assign  booth_double[4]=~(~(booth_in[8] & booth_in[9] & ~booth_in[10]) & ~(~booth_in[8] & ~booth_in[9] & booth_in[10]));

endmodule // booth_encoder

///////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps 

module booth_selector(pp_out,booth_single, booth_double, booth_negtive,multiplicand, signed_mpy);
input	[7:0]multiplicand;
input	[4:0]booth_single;
input	[4:0]booth_double;
input	[4:0]booth_negtive;
output	[44:0] pp_out;
integer	j;

reg		[8:0] pp0,pp1,pp2,pp3,pp4;

input	signed_mpy;
wire	sign_ext;
assign sign_ext=(signed_mpy==1'b1)?{multiplicand[7]} : 1'b0;


assign pp_out ={pp4, pp3, pp2, pp1, pp0};

wire	[9:0]bs_in;

assign  bs_in={sign_ext ,multiplicand[7:0],1'b0};


always @(booth_negtive or booth_single or bs_in or booth_double)

begin
	for (j=0; j<=8; j=j+1)
	begin
		pp0[j] = (booth_negtive[0]^ ~(~(booth_single[0] & bs_in[j+1]) & ~(booth_double[0] & bs_in[j])));
		pp1[j] = (booth_negtive[1]^ ~(~(booth_single[1] & bs_in[j+1]) & ~(booth_double[1] & bs_in[j])));
		pp2[j] = (booth_negtive[2]^ ~(~(booth_single[2] & bs_in[j+1]) & ~(booth_double[2] & bs_in[j])));
		pp3[j] = (booth_negtive[3]^ ~(~(booth_single[3] & bs_in[j+1]) & ~(booth_double[3] & bs_in[j])));
		pp4[j] = (booth_negtive[4]^ ~(~(booth_single[4] & bs_in[j+1]) & ~(booth_double[4] & bs_in[j])));
	end

end 

endmodule // booth_selector

///////////////////////////////////////////////////////////////////////
`timescale 1ns / 1ps

module MPY8x8(csa_a,csa_b,multiplicand,multiplier,signed_MPD,signed_MPR);
input	[7:0]multiplicand;
input	[7:0]multiplier;
input	signed_MPD, signed_MPR;

output [15:0] csa_a;
output [15:0] csa_b;

wire	[4:0]booth_single;
wire	[4:0]booth_double;
wire	[4:0]booth_negtive;
wire	[4:0]pp_sign;

wire	[44:0]pp_out;
wire	[8:0] PP0,PP1,PP2,PP3,PP4;

assign {PP4, PP3, PP2, PP1, PP0} = pp_out;

booth_encoder booth_encoder
(
.booth_single(booth_single), 
.booth_double(booth_double), 
.booth_negtive(booth_negtive), 
.multiplier(multiplier),
.signed_mpy(signed_MPR)
);


booth_selector booth_selector
(
.pp_out(pp_out),
.booth_single(booth_single), 
.booth_double(booth_double), 
.booth_negtive(booth_negtive),
.multiplicand(multiplicand),
.signed_mpy(signed_MPD)
);

wire	current_MPD_sign;
assign current_MPD_sign = multiplicand[7] & signed_MPD;
//assign pp_sign[0] = (booth_negtive[0] ^ current_MPD_sign) & (booth_single[0] | booth_double[0] | booth_negtive[0]) | (~booth_single[0] & ~booth_double[0] & booth_negtive[0]);
//assign pp_sign[1] = (booth_negtive[1] ^ current_MPD_sign) & (booth_single[1] | booth_double[1] | booth_negtive[1]) | (~booth_single[1] & ~booth_double[1] & booth_negtive[1]);
//assign pp_sign[2] = (booth_negtive[2] ^ current_MPD_sign) & (booth_single[2] | booth_double[2] | booth_negtive[2]) | (~booth_single[2] & ~booth_double[2] & booth_negtive[2]);
//assign pp_sign[3] = (booth_negtive[3] ^ current_MPD_sign) & (booth_single[3] | booth_double[3] | booth_negtive[3]) | (~booth_single[3] & ~booth_double[3] & booth_negtive[3]);
//assign pp_sign[4] = (booth_negtive[4] ^ current_MPD_sign) & (booth_single[4] | booth_double[4] | booth_negtive[4]) | (~booth_single[4] & ~booth_double[4] & booth_negtive[4]);

integer j;
reg [4:0] booth_single_b, booth_double_b, booth_negtive_b;

always @(booth_single or booth_double or booth_negtive)
begin
	for (j=0; j<=4; j=j+1)
	begin
		booth_single_b[j] = ~booth_single[j];
		booth_double_b[j] = ~booth_double[j];
		booth_negtive_b[j] = ~booth_negtive[j];
	end
end 

assign pp_sign[0] = (booth_negtive[0] ^ current_MPD_sign) & ~(booth_single_b[0] & booth_double_b[0] & booth_negtive_b[0]) | (booth_single_b[0] & booth_double_b[0] & booth_negtive[0]);
assign pp_sign[1] = (booth_negtive[1] ^ current_MPD_sign) & ~(booth_single_b[1] & booth_double_b[1] & booth_negtive_b[1]) | (booth_single_b[1] & booth_double_b[1] & booth_negtive[1]);
assign pp_sign[2] = (booth_negtive[2] ^ current_MPD_sign) & ~(booth_single_b[2] & booth_double_b[2] & booth_negtive_b[2]) | (booth_single_b[2] & booth_double_b[2] & booth_negtive[2]);
assign pp_sign[3] = (booth_negtive[3] ^ current_MPD_sign) & ~(booth_single_b[3] & booth_double_b[3] & booth_negtive_b[3]) | (booth_single_b[3] & booth_double_b[3] & booth_negtive[3]);
assign pp_sign[4] = (booth_negtive[4] ^ current_MPD_sign) & ~(booth_single_b[4] & booth_double_b[4] & booth_negtive_b[4]) | (booth_single_b[4] & booth_double_b[4] & booth_negtive[4]);
// Wallace CSA step#1

wire	FA1_R00C14_C, FA1_R00C14_S;
wire	FA1_R00C13_C, FA1_R00C13_S;
wire	FA1_R00C12_C, FA1_R00C12_S;

wire	FA1_R00C11_C, FA1_R00C11_S;
wire	HA1_R03C11_C, HA1_R03C11_S;

wire	FA1_R00C10_C, FA1_R00C10_S;
wire	HA1_R03C10_C, HA1_R03C10_S;

wire	FA1_R00C09_C, FA1_R00C09_S;
wire	HA1_R03C09_C, HA1_R03C09_S;

wire	FA1_R00C08_C, FA1_R00C08_S;
wire	FA1_R03C08_C, FA1_R03C08_S;

wire	FA1_R00C07_C, FA1_R00C07_S;
wire	FA1_R00C06_C, FA1_R00C06_S;
wire	HA1_R03C06_C, HA1_R03C06_S;

wire	FA1_R00C05_C, FA1_R00C05_S;
wire	FA1_R00C04_C, FA1_R00C04_S;

wire	FA1_R00C02_C, FA1_R00C02_S;


fa FA1_R00C14(.Cout(FA1_R00C14_C), .Sum(FA1_R00C14_S), .A(1'b1), .B(PP3[8]), .C(PP4[6]));

fa FA1_R00C13(.Cout(FA1_R00C13_C), .Sum(FA1_R00C13_S), .A(~pp_sign[2]), .B(PP3[7]), .C(PP4[5]));

fa FA1_R00C12(.Cout(FA1_R00C12_C), .Sum(FA1_R00C12_S), .A(1'b1), .B(PP2[8]), .C(PP3[6]));

fa FA1_R00C11(.Cout(FA1_R00C11_C), .Sum(FA1_R00C11_S), .A(~pp_sign[0]), .B(~pp_sign[1]), .C(PP2[7]));
ha HA1_R03C11(.Cout(HA1_R03C11_C), .Sum(HA1_R03C11_S), .A(PP3[5]), .B(PP4[3]));

fa FA1_R00C10(.Cout(FA1_R00C10_C), .Sum(FA1_R00C10_S), .A(pp_sign[0]), .B(PP1[8]), .C(PP2[6]));
ha HA1_R03C10(.Cout(HA1_R03C10_C), .Sum(HA1_R03C10_S), .A(PP3[4]), .B(PP4[2]));

fa FA1_R00C09(.Cout(FA1_R00C09_C), .Sum(FA1_R00C09_S), .A(pp_sign[0]), .B(PP1[7]), .C(PP2[5]));
ha HA1_R03C09(.Cout(HA1_R03C09_C), .Sum(HA1_R03C09_S), .A(PP3[3]), .B(PP4[1]));

fa FA1_R00C08(.Cout(FA1_R00C08_C), .Sum(FA1_R00C08_S), .A(PP0[8]), .B(PP1[6]), .C(PP2[4]));
fa FA1_R03C08(.Cout(FA1_R03C08_C), .Sum(FA1_R03C08_S), .A(PP3[2]), .B(PP4[0]), .C(booth_negtive[4]));

fa FA1_R00C07(.Cout(FA1_R00C07_C), .Sum(FA1_R00C07_S), .A(PP0[7]), .B(PP1[5]), .C(PP2[3]));
fa FA1_R00C06(.Cout(FA1_R00C06_C), .Sum(FA1_R00C06_S), .A(PP0[6]), .B(PP1[4]), .C(PP2[2]));
ha HA1_R03C06(.Cout(HA1_R03C06_C), .Sum(HA1_R03C06_S), .A(PP3[0]), .B(booth_negtive[3]));

fa FA1_R00C05(.Cout(FA1_R00C05_C), .Sum(FA1_R00C05_S), .A(PP0[5]), .B(PP1[3]), .C(PP2[1]));
fa FA1_R00C04(.Cout(FA1_R00C04_C), .Sum(FA1_R00C04_S), .A(PP0[4]), .B(PP1[2]), .C(PP2[0]));

fa FA1_R00C02(.Cout(FA1_R00C02_C), .Sum(FA1_R00C02_S), .A(PP0[2]), .B(PP1[0]), .C(booth_negtive[1]));

// Wallace CSA step#2

wire	FA2_R00C15_C, FA2_R00C15_S;
wire	HA2_R00C14_C, HA2_R00C14_S;
wire	HA2_R00C13_C, HA2_R00C13_S;

wire	FA2_R00C12_C, FA2_R00C12_S;
wire	FA2_R00C11_C, FA2_R00C11_S;
wire	FA2_R00C10_C, FA2_R00C10_S;
wire	FA2_R00C09_C, FA2_R00C09_S;
wire	FA2_R00C08_C, FA2_R00C08_S;
wire	FA2_R00C07_C, FA2_R00C07_S;
wire	FA2_R00C06_C, FA2_R00C06_S;

wire	FA2_R00C03_C, FA2_R00C03_S;


fa FA2_R00C15(.Cout(FA2_R00C15_C), .Sum(FA2_R00C15_S), .A(~pp_sign[3]), .B(PP4[7]), .C(FA1_R00C14_C));

ha HA2_R00C14(.Cout(HA2_R00C14_C), .Sum(HA2_R00C14_S), .A(FA1_R00C14_S), .B(FA1_R00C13_C));
ha HA2_R00C13(.Cout(HA2_R00C13_C), .Sum(HA2_R00C13_S), .A(FA1_R00C13_S), .B(FA1_R00C12_C));

fa FA2_R00C12(.Cout(FA2_R00C12_C), .Sum(FA2_R00C12_S), .A(FA1_R00C12_S), .B(FA1_R00C11_C), .C(HA1_R03C11_C));
fa FA2_R00C11(.Cout(FA2_R00C11_C), .Sum(FA2_R00C11_S), .A(FA1_R00C11_S), .B(FA1_R00C10_C), .C(HA1_R03C11_S));
fa FA2_R00C10(.Cout(FA2_R00C10_C), .Sum(FA2_R00C10_S), .A(FA1_R00C10_S), .B(FA1_R00C09_C), .C(HA1_R03C10_S));
fa FA2_R00C09(.Cout(FA2_R00C09_C), .Sum(FA2_R00C09_S), .A(FA1_R00C09_S), .B(FA1_R00C08_C), .C(HA1_R03C09_S));
fa FA2_R00C08(.Cout(FA2_R00C08_C), .Sum(FA2_R00C08_S), .A(FA1_R00C08_S), .B(FA1_R00C07_C), .C(FA1_R03C08_S));
fa FA2_R00C07(.Cout(FA2_R00C07_C), .Sum(FA2_R00C07_S), .A(FA1_R00C07_S), .B(FA1_R00C06_C), .C(HA1_R03C06_C));
fa FA2_R00C06(.Cout(FA2_R00C06_C), .Sum(FA2_R00C06_S), .A(FA1_R00C06_S), .B(FA1_R00C05_C), .C(HA1_R03C06_S));

fa FA2_R00C03(.Cout(FA2_R00C03_C), .Sum(FA2_R00C03_S), .A(PP0[3]), .B(PP1[1]), .C(FA1_R00C02_C));

// Wallace CSA step#3
wire	HA3_R00C15_C, HA3_R00C15_S;
wire	HA3_R00C14_C, HA3_R00C14_S;
wire	HA3_R00C13_C, HA3_R00C13_S;
wire	FA3_R00C12_C, FA3_R00C12_S;
wire	FA3_R00C11_C, FA3_R00C11_S;
wire	FA3_R00C10_C, FA3_R00C10_S;
wire	FA3_R00C09_C, FA3_R00C09_S;

wire	HA3_R00C08_C, HA3_R00C08_S;
wire	FA3_R00C07_C, FA3_R00C07_S;

wire	HA3_R00C05_C, HA3_R00C05_S;
wire	FA3_R00C04_C, FA3_R00C04_S;


ha HA3_R00C15(.Cout(HA3_R00C15_C), .Sum(HA3_R00C15_S), .A(FA2_R00C15_S), .B(HA2_R00C14_C));
ha HA3_R00C14(.Cout(HA3_R00C14_C), .Sum(HA3_R00C14_S), .A(HA2_R00C14_S), .B(HA2_R00C13_C));
ha HA3_R00C13(.Cout(HA3_R00C13_C), .Sum(HA3_R00C13_S), .A(HA2_R00C13_S), .B(FA2_R00C12_C));
fa FA3_R00C12(.Cout(FA3_R00C12_C), .Sum(FA3_R00C12_S), .A(FA2_R00C12_S), .B(FA2_R00C11_C), .C(PP4[4]));
fa FA3_R00C11(.Cout(FA3_R00C11_C), .Sum(FA3_R00C11_S), .A(FA2_R00C11_S), .B(FA2_R00C10_C), .C(HA1_R03C10_C));
fa FA3_R00C10(.Cout(FA3_R00C10_C), .Sum(FA3_R00C10_S), .A(FA2_R00C10_S), .B(FA2_R00C09_C), .C(HA1_R03C09_C));
fa FA3_R00C09(.Cout(FA3_R00C09_C), .Sum(FA3_R00C09_S), .A(FA2_R00C09_S), .B(FA2_R00C08_C), .C(FA1_R03C08_C));

ha HA3_R00C08(.Cout(HA3_R00C08_C), .Sum(HA3_R00C08_S), .A(FA2_R00C08_S), .B(FA2_R00C07_C));
fa FA3_R00C07(.Cout(FA3_R00C07_C), .Sum(FA3_R00C07_S), .A(FA2_R00C07_S), .B(FA2_R00C06_C), .C(PP3[1]));

ha HA3_R00C05(.Cout(HA3_R00C05_C), .Sum(HA3_R00C05_S), .A(FA1_R00C05_S), .B(FA1_R00C04_C));
fa FA3_R00C04(.Cout(FA3_R00C04_C), .Sum(FA3_R00C04_S), .A(FA1_R00C04_S), .B(booth_negtive[2]), .C(FA2_R00C03_C));


assign csa_a[0] = PP0[0];
assign csa_b[0] = booth_negtive[0];
assign csa_a[1] = PP0[1];
assign csa_b[1] = 1'b0;
assign csa_a[2] = FA1_R00C02_S;
assign csa_b[2] = 1'b0;
assign csa_a[3] = FA2_R00C03_S;
assign csa_b[3] = 1'b0;

assign csa_a[4] = FA3_R00C04_S;
assign csa_b[4] = 1'b0;

assign csa_a[5] = HA3_R00C05_S;
assign csa_b[5] = FA3_R00C04_C;
assign csa_a[6] = FA2_R00C06_S;
assign csa_b[6] = HA3_R00C05_C;
assign csa_a[7] = FA3_R00C07_S;
assign csa_b[7] = 1'b0;
assign csa_a[8] = HA3_R00C08_S;
assign csa_b[8] = FA3_R00C07_C;
assign csa_a[9] = FA3_R00C09_S;
assign csa_b[9] = HA3_R00C08_C;
assign csa_a[10] = FA3_R00C10_S;
assign csa_b[10] = FA3_R00C09_C;
assign csa_a[11] = FA3_R00C11_S;
assign csa_b[11] = FA3_R00C10_C;
assign csa_a[12] = FA3_R00C12_S;
assign csa_b[12] = FA3_R00C11_C;
assign csa_a[13] = HA3_R00C13_S;
assign csa_b[13] = FA3_R00C12_C;
assign csa_a[14] = HA3_R00C14_S;
assign csa_b[14] = HA3_R00C13_C;
assign csa_a[15] = HA3_R00C15_S;
assign csa_b[15] = HA3_R00C14_C;

endmodule // MPY8x8

///////////////////////////////////////////////////////////////////////
`timescale 1ns / 1ps
module MPY16X16(
clk,

IHRST,
ILRST,

FSEL,
GSEL,
HSEL,
JKSEL,
MPY_8X8_MODE,

ASGND,
BSGND,

A,
B,

OH_8X8,
OL_8X8,
O_16X16
);

input clk;

input IHRST;
input ILRST;

input FSEL;
input GSEL;
input HSEL;
input JKSEL;
input MPY_8X8_MODE;

input ASGND;
input BSGND;

input	[15:0]A;
input	[15:0]B;

output [15:0] OH_8X8;
output [15:0] OL_8X8;
output [31:0] O_16X16;


reg 	[31:0]csa_rega, csa_regb;
wire	[152:0]pp_out;

wire	[7:0] MPYG_mpd, MPYG_mpr;
wire	[7:0] MPYJ_mpd, MPYJ_mpr;
wire	[7:0] MPYF_mpd, MPYF_mpr;
wire	[7:0] MPYK_mpd, MPYK_mpr;

wire	MPYG_MPD_sign, MPYG_MPR_sign;
wire	MPYJ_MPD_sign, MPYJ_MPR_sign;
wire	MPYF_MPD_sign, MPYF_MPR_sign;
wire	MPYK_MPD_sign, MPYK_MPR_sign;

assign MPYG_mpd = A[7:0];
assign MPYG_mpr = B[7:0];
assign MPYG_MPD_sign = MPY_8X8_MODE ? ASGND : `UNSIGNED_DATA;
assign MPYG_MPR_sign = MPY_8X8_MODE ? BSGND : `UNSIGNED_DATA;

assign MPYJ_mpd = A[7:0];
assign MPYJ_mpr = B[15:8];
assign MPYJ_MPD_sign = `UNSIGNED_DATA;
assign MPYJ_MPR_sign = BSGND;

assign MPYF_mpd = A[15:8];
assign MPYF_mpr = B[15:8];
assign MPYF_MPD_sign = ASGND;
assign MPYF_MPR_sign = BSGND;

assign MPYK_mpd = A[15:8];
assign MPYK_mpr = B[7:0];
assign MPYK_MPD_sign = ASGND;
assign MPYK_MPR_sign = `UNSIGNED_DATA;

wire	[15:0] MPYG_csa_a, MPYG_csa_b;
wire	[15:0] MPYJ_csa_a, MPYJ_csa_b;
wire	[15:0] MPYF_csa_a, MPYF_csa_b;
wire	[15:0] MPYK_csa_a, MPYK_csa_b;

wire	[15:0] MPYG_o, MPYG_out;
wire	[15:0] MPYJ_o, MPYJ_out;
wire	[15:0] MPYF_o, MPYF_out;
wire	[15:0] MPYK_o, MPYK_out;
reg		[15:0] MPYG_oreg, MPYJ_oreg;
reg		[15:0] MPYF_oreg, MPYK_oreg;

wire	MPYJ_out_sign, MPYK_out_sign;
wire	MPYJK_g, MPYJK_p;

assign MPYJ_out_sign = BSGND ? MPYJ_out[15] : `UNSIGNED_DATA;
assign MPYK_out_sign = ASGND ? MPYK_out[15] : `UNSIGNED_DATA;

assign MPYJK_g = MPYJ_out_sign & MPYK_out_sign;
assign MPYJK_p = MPYJ_out_sign ^ MPYK_out_sign;


MPY8x8 MPY_G(.csa_a(MPYG_csa_a),.csa_b(MPYG_csa_b),.multiplicand(MPYG_mpd),.multiplier(MPYG_mpr),.signed_MPD(MPYG_MPD_sign),.signed_MPR(MPYG_MPR_sign));
MPY8x8 MPY_J(.csa_a(MPYJ_csa_a),.csa_b(MPYJ_csa_b),.multiplicand(MPYJ_mpd),.multiplier(MPYJ_mpr),.signed_MPD(MPYJ_MPD_sign),.signed_MPR(MPYJ_MPR_sign));
MPY8x8 MPY_F(.csa_a(MPYF_csa_a),.csa_b(MPYF_csa_b),.multiplicand(MPYF_mpd),.multiplier(MPYF_mpr),.signed_MPD(MPYF_MPD_sign),.signed_MPR(MPYF_MPR_sign));
MPY8x8 MPY_K(.csa_a(MPYK_csa_a),.csa_b(MPYK_csa_b),.multiplicand(MPYK_mpd),.multiplier(MPYK_mpr),.signed_MPD(MPYK_MPD_sign),.signed_MPR(MPYK_MPR_sign));



wire	[15:0] MPYG_cla_ina, MPYG_cla_inb;

assign MPYG_cla_ina = MPYG_csa_a;
assign MPYG_cla_inb = MPYG_csa_b;

wire	CLA16_G_g, CLA16_G_p, MPYG_ci;
assign MPYG_ci = 1'b0;

wire dangle_g_nodeJ, dangle_p_nodeJ; 
wire dangle_g_nodeF, dangle_p_nodeF; 
wire dangle_g_nodeK, dangle_p_nodeK; 



fcla16 CLA16_G(
.Sum(MPYG_o[15:0]),
.A(MPYG_cla_ina[15:0]),
.B(MPYG_cla_inb[15:0]), 
.G(CLA16_G_g),
.P(CLA16_G_p),
.Cin(MPYG_ci)
);



fcla16 CLA16_J(
.Sum(MPYJ_o[15:0]),
.A(MPYJ_csa_a[15:0]),
.B(MPYJ_csa_b[15:0]), 
.Cin(1'b0),
.G(dangle_g_nodeJ),
.P(dangle_p_nodeJ)
);



fcla16 CLA16_F(
.Sum(MPYF_o[15:0]),
.A(MPYF_csa_a[15:0]),
.B(MPYF_csa_b[15:0]), 
.Cin(1'b0),
.G(dangle_g_nodeF),
.P(dangle_p_nodeF)
);


fcla16 CLA16_K(
.Sum(MPYK_o[15:0]),
.A(MPYK_csa_a[15:0]),
.B(MPYK_csa_b[15:0]), 
.Cin(1'b0),
.G(dangle_g_nodeK), 
.P(dangle_p_nodeK)
);



always @(posedge clk or posedge IHRST)
begin
  if (IHRST)
    MPYF_oreg <= 0;		//#1 0;
  else
    MPYF_oreg <= MPYF_o; 	//#1 MPYF_o;
end

always @(posedge clk or posedge IHRST)
begin
  if (IHRST)
    MPYJ_oreg <=0; 		//#1 0;
  else if (MPY_8X8_MODE)
    MPYJ_oreg <=MPYJ_oreg;	//#1 MPYJ_oreg;
  else
    MPYJ_oreg <=MPYJ_o;  	//#1 MPYJ_o;
end

always @(posedge clk or posedge ILRST)
begin
  if (ILRST)
    MPYK_oreg <=0; 		//#1 0;
  else if (MPY_8X8_MODE)
    MPYK_oreg <=MPYK_oreg; 	//#1 MPYK_oreg;
  else
    MPYK_oreg <=MPYK_o; 	//#1 MPYK_o;
end

always @(posedge clk or posedge ILRST)
begin
  if (ILRST)
    MPYG_oreg <= 0; 		//#1 0;
  else
    MPYG_oreg <= MPYG_o; 	//#1 MPYG_o;
end

 assign MPYG_out = GSEL ? MPYG_oreg : MPYG_o;
 assign MPYJ_out = JKSEL ? MPYJ_oreg : MPYJ_o;

 assign MPYF_out = JKSEL ? MPYF_oreg : MPYF_o;
 assign MPYK_out = FSEL ? MPYK_oreg : MPYK_o;

wire [23:0] csa_oc;
wire [23:0] csa_os;
wire MPYJK_g_b;
assign MPYJK_g_b = ~MPYJK_g;

assign csa_os[23] = MPYJK_p ^ MPYF_out[15];
assign csa_oc[23] = ~(MPYJK_g_b & ~(MPYJK_p & MPYF_out[15]));
assign csa_os[22] = MPYJK_p ^ MPYF_out[14];
assign csa_oc[22] = ~(MPYJK_g_b & ~(MPYJK_p & MPYF_out[14]));
assign csa_os[21] = MPYJK_p ^ MPYF_out[13];
assign csa_oc[21] = ~(MPYJK_g_b & ~(MPYJK_p & MPYF_out[13]));
assign csa_os[20] = MPYJK_p ^ MPYF_out[12];
assign csa_oc[20] = ~(MPYJK_g_b & ~(MPYJK_p & MPYF_out[12]));
assign csa_os[19] = MPYJK_p ^ MPYF_out[11];
assign csa_oc[19] = ~(MPYJK_g_b & ~(MPYJK_p & MPYF_out[11]));
assign csa_os[18] = MPYJK_p ^ MPYF_out[10];
assign csa_oc[18] = ~(MPYJK_g_b & ~(MPYJK_p & MPYF_out[10]));
assign csa_os[17] = MPYJK_p ^ MPYF_out[9];
assign csa_oc[17] = ~(MPYJK_g_b & ~(MPYJK_p & MPYF_out[9]));
assign csa_os[16] = MPYJK_p ^ MPYF_out[8];
assign csa_oc[16] = ~(MPYJK_g_b & ~(MPYJK_p & MPYF_out[8]));

fa FA1_R00C15(.Cout(csa_oc[15]), .Sum(csa_os[15]), .A(MPYJ_out[15]), .B(MPYK_out[15]), .C(MPYF_out[7]));
fa FA1_R00C14(.Cout(csa_oc[14]), .Sum(csa_os[14]), .A(MPYJ_out[14]), .B(MPYK_out[14]), .C(MPYF_out[6]));
fa FA1_R00C13(.Cout(csa_oc[13]), .Sum(csa_os[13]), .A(MPYJ_out[13]), .B(MPYK_out[13]), .C(MPYF_out[5]));
fa FA1_R00C12(.Cout(csa_oc[12]), .Sum(csa_os[12]), .A(MPYJ_out[12]), .B(MPYK_out[12]), .C(MPYF_out[4]));
fa FA1_R00C11(.Cout(csa_oc[11]), .Sum(csa_os[11]), .A(MPYJ_out[11]), .B(MPYK_out[11]), .C(MPYF_out[3]));
fa FA1_R00C10(.Cout(csa_oc[10]), .Sum(csa_os[10]), .A(MPYJ_out[10]), .B(MPYK_out[10]), .C(MPYF_out[2]));
fa FA1_R00C09(.Cout(csa_oc[9]),  .Sum(csa_os[9]),  .A(MPYJ_out[9]),  .B(MPYK_out[9]),  .C(MPYF_out[1]));
fa FA1_R00C08(.Cout(csa_oc[8]),  .Sum(csa_os[8]),  .A(MPYJ_out[8]),  .B(MPYK_out[8]),  .C(MPYF_out[0]));

fa FA1_R00C07(.Cout(csa_oc[7]), .Sum(csa_os[7]), .A(MPYG_out[15]), .B(MPYJ_out[7]), .C(MPYK_out[7]));
fa FA1_R00C06(.Cout(csa_oc[6]), .Sum(csa_os[6]), .A(MPYG_out[14]), .B(MPYJ_out[6]), .C(MPYK_out[6]));
fa FA1_R00C05(.Cout(csa_oc[5]), .Sum(csa_os[5]), .A(MPYG_out[13]), .B(MPYJ_out[5]), .C(MPYK_out[5]));
fa FA1_R00C04(.Cout(csa_oc[4]), .Sum(csa_os[4]), .A(MPYG_out[12]), .B(MPYJ_out[4]), .C(MPYK_out[4]));
fa FA1_R00C03(.Cout(csa_oc[3]), .Sum(csa_os[3]), .A(MPYG_out[11]), .B(MPYJ_out[3]), .C(MPYK_out[3]));
fa FA1_R00C02(.Cout(csa_oc[2]), .Sum(csa_os[2]), .A(MPYG_out[10]), .B(MPYJ_out[2]), .C(MPYK_out[2]));
fa FA1_R00C01(.Cout(csa_oc[1]), .Sum(csa_os[1]), .A(MPYG_out[9]),  .B(MPYJ_out[1]), .C(MPYK_out[1]));
fa FA1_R00C00(.Cout(csa_oc[0]), .Sum(csa_os[0]), .A(MPYG_out[8]),  .B(MPYJ_out[0]), .C(MPYK_out[0]));


wire 	[23:0] cla_ina;
wire 	[23:0] cla_inb;

wire 	[23:0] cla_o;
wire	cla24_g0, cla24_p0;
wire	cla24_g1, cla24_p1;

wire	cla24_cin, cla24_16_cout;

assign cla_ina = csa_os;
assign cla_inb = {csa_oc[22:0],1'b0};
assign cla24_cin = 1'b0 ;


fcla16 CLA24_16(
.Sum(cla_o[15:0]),
.G(cla24_g0),
.P(cla24_p0), 
.A(cla_ina[15:0]),
.B(cla_inb[15:0]), 
.Cin(cla24_cin)
);
assign cla24_16_cout = ~(~cla24_g0 & ~(cla24_p0 & cla24_cin));



fcla8 CLA24_8(
.Sum(cla_o[23:16]),
.G(cla24_g1),
.P(cla24_p1), 
.A(cla_ina[23:16]),
.B(cla_inb[23:16]), 
.Cin(cla24_16_cout)
);

reg 	[31:0]mpy16_reg;

always @(posedge clk or posedge ILRST)
begin
  if (ILRST)
    mpy16_reg <= 0; 		//#1 0;
  else if (MPY_8X8_MODE)
    mpy16_reg <=  mpy16_reg; 	//#1 mpy16_reg;
  else
    mpy16_reg <={cla_o,MPYG_out[7:0]}; 	//#1 {cla_o,MPYG_out[7:0]};
end

assign O_16X16[31:0] = HSEL ? mpy16_reg : {cla_o,MPYG_out[7:0]};

assign OH_8X8 = MPYF_out[15:0];
assign OL_8X8 = MPYG_out[15:0];

endmodule // MPY16x16


//////////////////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps

module MULT_ACCUM(
    DIRECT_INPUT,
    MULT_INPUT,
    MULT_8x8,
    MULT_16x16,
	ADDSUB,
	CLK,
    CICAS,
    CI,
	SIGNEXTIN,
	SIGNEXTOUT,
    LDA,
    RST,
    ENA,
    COCAS,
    CO,
    O,
	OUTMUX_SEL,
	CARRYMUX_SEL,
	ADDER_A_IN_SEL,
	ADDER_B_IN_SEL
    );
	
    input [15:0] DIRECT_INPUT;
    input [15:0] MULT_INPUT;
    input [15:0] MULT_8x8;
    input [15:0] MULT_16x16;
    input ADDSUB;
    input CLK;
    input CICAS;
    input CI;
    input SIGNEXTIN;
    output SIGNEXTOUT;
    input LDA;
    input RST;
    input ENA;
    output COCAS;
    output CO;
    output [15:0] O;
	input [1:0] OUTMUX_SEL;
	input [1:0] CARRYMUX_SEL;
	input ADDER_A_IN_SEL;
	input [1:0] ADDER_B_IN_SEL;

	
	 wire [15:0] ADDER_LOAD_MUX ;
	 wire [15:0] ACCUMULATOR_REG ;
	 wire [15:0] ADDER_SUM ;
	 wire [15:0] ADDER_A_INPUT_MUX ;
	 wire [15:0] ADDER_B_INPUT_MUX ;
	 wire ADDER_CI ;
	 
	 assign SIGNEXTOUT = ADDER_B_INPUT_MUX[15];
	 

OUT_MUX_4 OUTPUT_MULTIPLEXER_TOP (
    .ADDER_COMBINATORIAL (ADDER_LOAD_MUX),
	 .ACCUM_REGISTER(ACCUMULATOR_REG) ,
	 .MULT_8x8(MULT_8x8) ,
	 .MULT_16x16(MULT_16x16),
	 .SELM(OUTMUX_SEL[1:0]) ,
	 .OUT(O)  
	 ) ;
	 
ACCUM_REG ACCUM_REG_TOP (
	.D(ADDER_LOAD_MUX) ,
	.Q(ACCUMULATOR_REG) ,
	.ENA(ENA) ,
	.CLK(CLK) ,
	.RST(RST)
	);
	
ACCUM_ADDER ACCUM_ADDER_TOP(
   .A(ADDER_A_INPUT_MUX) ,
   .B(ADDER_B_INPUT_MUX) ,
	.ADDSUB(ADDSUB) ,
	.CI(ADDER_CI) ,
	.SUM(ADDER_SUM) ,
	.COCAS(COCAS) ,
	.CO(CO)
	);	

LOAD_ADD_MUX LOAD_ADD_TOP (
   .ADDER(ADDER_SUM) ,
	.LOAD_DATA(DIRECT_INPUT) ,
	.LOAD(LDA),
	.OUT(ADDER_LOAD_MUX)
   );
	
ADDER_A_IN_MUX ADDER_A_IN_MUX_TOP (
   .ACCUMULATOR_REG(ACCUMULATOR_REG),
	.DIRECT_INPUT(DIRECT_INPUT) ,
	.SELM(ADDER_A_IN_SEL) ,
	.ADDER_A_MUX(ADDER_A_INPUT_MUX)
   );

ADDER_B_IN_MUX ADDER_B_IN_MUX_TOP (
   .MULT_INPUT(MULT_INPUT) ,
	.MULT_8x8(MULT_8x8) ,
	.MULT_16x16(MULT_16x16) ,
	.SIGNEXTIN(SIGNEXTIN) ,
	.SELM(ADDER_B_IN_SEL[1:0]) ,
	.ADDER_B_MUX(ADDER_B_INPUT_MUX)
	);	

CARRY_IN_MUX CARRY_IN_MUX_TOP (
	.CICAS(CICAS),
	.CI(CI),
	.CARRYMUX_SEL(CARRYMUX_SEL[1:0]),
	.ADDER_CI(ADDER_CI)
	);
	
endmodule

///////////////////////////////////////////////////////////////////////////////////
`timescale 1ns / 1ps

module OUT_MUX_4 (
    ADDER_COMBINATORIAL ,
	ACCUM_REGISTER ,
	MULT_8x8 ,
	MULT_16x16 ,
	SELM ,
	OUT  
	 ) ;

    input [15:0] ADDER_COMBINATORIAL ;
	input [15:0] ACCUM_REGISTER ;
	input [15:0] MULT_8x8 ;
	input [15:0] MULT_16x16 ;
	input [1:0] SELM ;
	output [15:0] OUT;  
	reg [15:0] OUT;  
	 
 
always @(SELM or ADDER_COMBINATORIAL or ACCUM_REGISTER or MULT_8x8 or MULT_16x16)
      case (SELM[1:0])
         2'b00: OUT = ADDER_COMBINATORIAL ; // Combinatorial output
         2'b01: OUT = ACCUM_REGISTER ; // Accumulator register output
         2'b10: OUT = MULT_8x8;  // MULT_8x8
         2'b11: OUT = MULT_16x16;  // MULT_16x16
      endcase	 

endmodule


///////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps

module ACCUM_REG (
	D ,
	Q ,
	ENA ,
	CLK ,
	RST
	);

	input [15:0] D ;
	output [15:0] Q;
	reg [15:0] Q;
	input ENA ;
	input CLK ;
	input RST;
	
	always @(posedge CLK or posedge RST)
      if (RST) // Syncronous reset overrides all other controls
				Q <= 16'h0 ;
		else
			if(ENA) // Update Q whenever LOAD or ENAble asserted
			    Q <=  D ; 	 //#1 D ;
			else
			    Q <= Q ;     //#1 Q ;
		
endmodule 


///////////////////////////////////////////////////////////////////////
`timescale 1ns / 1ps

module LOAD_ADD_MUX (
    ADDER ,
	LOAD_DATA ,
	LOAD,
	OUT
   );

	input [15:0] ADDER ;
	input [15:0] LOAD_DATA ;
	input LOAD;
	output [15:0] OUT;
   
	assign OUT = ( (LOAD) ? LOAD_DATA : ADDER ) ;
	
endmodule


///////////////////////////////////////////////////////////////////////
`timescale 1ns / 1ps

module ADDER_A_IN_MUX (
    ACCUMULATOR_REG ,
	DIRECT_INPUT ,
	SELM ,
	ADDER_A_MUX
   );
	
    input [15:0] ACCUMULATOR_REG ;
	input [15:0] DIRECT_INPUT ;
	input SELM ;
	output [15:0] ADDER_A_MUX;

	assign ADDER_A_MUX = ( (SELM) ? DIRECT_INPUT : ACCUMULATOR_REG ) ;

endmodule


///////////////////////////////////////////////////////////////////////
`timescale 1ns / 1ps

module ADDER_B_IN_MUX (
    MULT_INPUT ,
	MULT_8x8 ,
	MULT_16x16 ,
	SIGNEXTIN ,
	SELM ,
	ADDER_B_MUX
	);

    input [15:0] MULT_INPUT ;
	input [15:0] MULT_8x8 ;
	input [15:0] MULT_16x16 ;
	input SIGNEXTIN ;
	input [1:0] SELM ;
	output [15:0] ADDER_B_MUX;
	
//	wire [15:0] DIRECT_8x8_SELECT ;
//	assign DIRECT_8x8_SELECT = ( (SELM[0]) ? MULT_8x8   : MULT_INPUT) ;
//	assign ADDER_B_MUX       = ( (SELM[1:0]=2'b10) ? MULT_16x16 : DIRECT_8x8_SELECT) ;

	reg [15:0] ADDER_B_MUX;
	
always @(SELM or MULT_INPUT or MULT_8x8 or MULT_16x16 or SIGNEXTIN)
      case (SELM[1:0])
         2'b00: ADDER_B_MUX = MULT_INPUT ; 
         2'b01: ADDER_B_MUX = MULT_8x8 ; 
         2'b10: ADDER_B_MUX = MULT_16x16; 
         2'b11: ADDER_B_MUX = {16{SIGNEXTIN}}; 
      endcase	 
	
endmodule


///////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps
module CARRY_IN_MUX (
	CICAS,
	CI,
	CARRYMUX_SEL,
	ADDER_CI
	);
	
	input CICAS;
	input CI;
	input [1:0] CARRYMUX_SEL;
	output ADDER_CI;
	reg ADDER_CI;
	
always @(CARRYMUX_SEL or CICAS or CI)
      case (CARRYMUX_SEL[1:0])
         2'b00: ADDER_CI = 0 ; 
         2'b01: ADDER_CI = 1 ; 
         2'b10: ADDER_CI = CICAS; 
         2'b11: ADDER_CI = CI; 
      endcase	 

endmodule
	
//////////////////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps

module ACCUM_ADDER (
	A ,
	B ,
	ADDSUB ,
	CI ,
	SUM ,
	COCAS ,
	CO
	);
//parameter A_width =16;
input [15:0] A ;
input [15:0] B ;
input ADDSUB ;
input CI ;
output [15:0] SUM ;
output COCAS, CO;

wire	CLA16_g, CLA16_p;
reg		CO;

wire [15:0] CLA16_SUM;
reg	[15:0] CLA16_A, SUM;
integer j;

always@(ADDSUB or COCAS or A or CLA16_SUM)
begin
	if (ADDSUB)
		begin
		   CO = ~COCAS;
           for (j=0; j<=15; j=j+1)
			begin
			 CLA16_A[j] = ~A[j];
			 SUM[j] = ~CLA16_SUM[j];
			end 
		end   
		else
		begin
		   CO = COCAS;
		   CLA16_A[15:0] = A[15:0];
		   SUM[15:0] = CLA16_SUM[15:0];
		end
end

fcla16 CLA16_ADDER(
.Sum(CLA16_SUM[15:0]),
.A(CLA16_A[15:0]),
.B(B[15:0]), 
.G(CLA16_g),
.P(CLA16_p),
.Cin(CI)
);
assign COCAS= ~(~CLA16_g & ~(CLA16_p & CI));


endmodule


///////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps

module ha (Cout, Sum, A, B);
input A, B;
output Cout, Sum;

assign Cout = A & B;
assign Sum  = A ^ B;

endmodule // ha

///////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps
module fa (Cout, Sum, A, B, C);
input A, B, C;
output Cout, Sum;

//assign Cout = ((A&B) | (B&C) |(A&C));

assign Cout = ~(~(A&B) & ~(B&C) & ~(A&C));
assign Sum  = A^B^C;

endmodule // fa

///////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps

module mpfa (g_b, p,Sum, A, B, Cin);
input A, B, Cin;
output g_b, p, Sum;


assign g_b = ~(A & B);
assign p = A ^ B;

assign Sum  = p ^ Cin;

endmodule // mpfa

///////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps

module mclg4 (cout, g_o, p_o, g_b, p, cin);
input [3:0] g_b, p;
input cin;
output [3:0] cout;
output g_o, p_o;

wire	s1, s2, s3, s4, s5, s6,s7,s8,s9;

wire  [2:0] g;
assign g[0] =~g_b[0];
assign g[1] =~g_b[1];
assign g[2] =~g_b[2];

assign s1 = ~(p[0] & cin);
assign cout[1] =~(g_b[0] & s1);

assign s2 = ~(p[1] & g[0]);
assign s3 = ~(p[1] & p[0] & cin);
assign cout[2] =~(g_b[1] & s2 & s3);

assign s4 = ~(p[2] & g[1]);
assign s5 = ~(p[2] & p[1] & g[0]);
assign s6 = ~(p[2] & p[1] & p[0] & cin);
assign cout[3] =~(g_b[2] & s4 & s5 & s6);

assign s7 =~(p[3] & g[2]);
assign s8 =~(p[3] & p[2] & g[1]);
assign s9 =~(p[3] & p[2] & p[1] & g[0]);
assign g_o =~(g_b[3] & s7 & s8 & s9);

assign p_o =(p[3] & p[2] & p[1] & p[0]);

endmodule // mclg4

///////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps

module mclg16 (cout, g_o, p_o, g, p, cin);
input [3:0] g, p;
input cin;
output [3:0] cout;
output g_o, p_o;

wire	s1, s2, s3, s4, s5, s6, s7,s8,s9;

assign s1 = ~(p[0] & cin);
assign cout[1] =~(~g[0] & s1);

assign s2 = ~(p[1] & g[0]);
assign s3 = ~(p[1] & p[0] & cin);
assign cout[2] =~(~g[1] & s2 & s3);

assign s4 = ~(p[2] & g[1]);
assign s5 = ~(p[2] & p[1] & g[0]);
assign s6 = ~(p[2] & p[1] & p[0] & cin);
assign cout[3] =~(~g[2] & s4 & s5 & s6);

assign s7 =~(p[3] & g[2]);
assign s8 =~(p[3] & p[2] & g[1]);
assign s9 =~(p[3] & p[2] & p[1] & g[0]);
assign g_o =~(~g[3] & s7 & s8 & s9);

assign p_o =(p[3] & p[2] & p[1] & p[0]);

endmodule // mclg16
///////////////////////////////////////////////////////////////////////


`timescale 1ns / 1ps
module fcla16 (Sum, G, P, A, B, Cin);
input [15:0] A, B;
input Cin;
output [15:0] Sum;
output G, P;
wire	[15:0] gtemp1_b;
wire	[15:0] ptemp1;
wire	[15:0] ctemp1;
wire	[3:0] ctemp2;

wire	[3:0] gouta, pouta;
mpfa r01 (.g_b(gtemp1_b[0]), .p(ptemp1[0]), .Sum(Sum[0]), .A(A[0]), .B(B[0]), .Cin(Cin));
mpfa r02 (.g_b(gtemp1_b[1]), .p(ptemp1[1]), .Sum(Sum[1]), .A(A[1]), .B(B[1]), .Cin(ctemp1[1]));
mpfa r03 (.g_b(gtemp1_b[2]), .p(ptemp1[2]), .Sum(Sum[2]), .A(A[2]), .B(B[2]), .Cin(ctemp1[2]));
mpfa r04 (.g_b(gtemp1_b[3]), .p(ptemp1[3]), .Sum(Sum[3]), .A(A[3]), .B(B[3]), .Cin(ctemp1[3]));
mclg4 b1 (.cout(ctemp1[3:0]), .g_o(gouta[0]), .p_o(pouta[0]), .g_b(gtemp1_b[3:0]), .p(ptemp1[3:0]), .cin(Cin));

mpfa r05 (.g_b(gtemp1_b[4]), .p(ptemp1[4]), .Sum(Sum[4]), .A(A[4]), .B(B[4]), .Cin(ctemp2[1]));
mpfa r06 (.g_b(gtemp1_b[5]), .p(ptemp1[5]), .Sum(Sum[5]), .A(A[5]), .B(B[5]), .Cin(ctemp1[5]));
mpfa r07 (.g_b(gtemp1_b[6]), .p(ptemp1[6]), .Sum(Sum[6]), .A(A[6]), .B(B[6]), .Cin(ctemp1[6]));
mpfa r08 (.g_b(gtemp1_b[7]), .p(ptemp1[7]), .Sum(Sum[7]), .A(A[7]), .B(B[7]), .Cin(ctemp1[7]));
mclg4 b2 (.cout(ctemp1[7:4]), .g_o(gouta[1]), .p_o(pouta[1]), .g_b(gtemp1_b[7:4]), .p(ptemp1[7:4]), .cin(ctemp2[1]));

mpfa r09 (.g_b(gtemp1_b[8]), .p(ptemp1[8]), .Sum(Sum[8]), .A(A[8]), .B(B[8]), .Cin(ctemp2[2]));
mpfa r10 (.g_b(gtemp1_b[9]), .p(ptemp1[9]), .Sum(Sum[9]), .A(A[9]), .B(B[9]), .Cin(ctemp1[9]));
mpfa r11 (.g_b(gtemp1_b[10]), .p(ptemp1[10]), .Sum(Sum[10]), .A(A[10]), .B(B[10]), .Cin(ctemp1[10]));
mpfa r12 (.g_b(gtemp1_b[11]), .p(ptemp1[11]), .Sum(Sum[11]), .A(A[11]), .B(B[11]), .Cin(ctemp1[11]));
mclg4 b3 (.cout(ctemp1[11:8]), .g_o(gouta[2]), .p_o(pouta[2]), .g_b(gtemp1_b[11:8]), .p(ptemp1[11:8]), .cin(ctemp2[2]));

mpfa r13 (.g_b(gtemp1_b[12]), .p(ptemp1[12]), .Sum(Sum[12]), .A(A[12]), .B(B[12]), .Cin(ctemp2[3]));
mpfa r14 (.g_b(gtemp1_b[13]), .p(ptemp1[13]), .Sum(Sum[13]), .A(A[13]), .B(B[13]), .Cin(ctemp1[13]));
mpfa r15 (.g_b(gtemp1_b[14]), .p(ptemp1[14]), .Sum(Sum[14]), .A(A[14]), .B(B[14]), .Cin(ctemp1[14]));
mpfa r16 (.g_b(gtemp1_b[15]), .p(ptemp1[15]), .Sum(Sum[15]), .A(A[15]), .B(B[15]), .Cin(ctemp1[15]));
mclg4 b4 (.cout(ctemp1[15:12]), .g_o(gouta[3]), .p_o(pouta[3]), .g_b(gtemp1_b[15:12]), .p(ptemp1[15:12]), .cin(ctemp2[3]));

mclg16 b5 (.cout(ctemp2), .g_o(G), .p_o(P), .g(gouta), .p(pouta), .cin(Cin));
endmodule // fcla16


///////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps

module fcla8 (Sum, G, P, A, B, Cin);
input [7:0] A, B;
input Cin;
output [7:0] Sum;
output G, P;
wire	[7:0] gtemp1;
wire	[7:0] ptemp1;
wire	[7:0] ctemp1;
wire	 ctemp2;

wire	[1:0] gouta, pouta;

mpfa r01 (.g_b(gtemp1[0]), .p(ptemp1[0]), .Sum(Sum[0]), .A(A[0]), .B(B[0]), .Cin(Cin));
mpfa r02 (.g_b(gtemp1[1]), .p(ptemp1[1]), .Sum(Sum[1]), .A(A[1]), .B(B[1]), .Cin(ctemp1[1]));
mpfa r03 (.g_b(gtemp1[2]), .p(ptemp1[2]), .Sum(Sum[2]), .A(A[2]), .B(B[2]), .Cin(ctemp1[2]));
mpfa r04 (.g_b(gtemp1[3]), .p(ptemp1[3]), .Sum(Sum[3]), .A(A[3]), .B(B[3]), .Cin(ctemp1[3]));
mclg4 b1 (.cout(ctemp1[3:0]), .g_o(gouta[0]), .p_o(pouta[0]), .g_b(gtemp1[3:0]), .p(ptemp1[3:0]), .cin(Cin));

mpfa r05 (.g_b(gtemp1[4]), .p(ptemp1[4]), .Sum(Sum[4]), .A(A[4]), .B(B[4]), .Cin(ctemp2));
mpfa r06 (.g_b(gtemp1[5]), .p(ptemp1[5]), .Sum(Sum[5]), .A(A[5]), .B(B[5]), .Cin(ctemp1[5]));
mpfa r07 (.g_b(gtemp1[6]), .p(ptemp1[6]), .Sum(Sum[6]), .A(A[6]), .B(B[6]), .Cin(ctemp1[6]));
mpfa r08 (.g_b(gtemp1[7]), .p(ptemp1[7]), .Sum(Sum[7]), .A(A[7]), .B(B[7]), .Cin(ctemp1[7]));
mclg4 b2 (.cout(ctemp1[7:4]), .g_o(gouta[1]), .p_o(pouta[1]), .g_b(gtemp1[7:4]), .p(ptemp1[7:4]), .cin(ctemp2));

assign ctemp2=~(~gouta[0] & ~(pouta[0] & Cin));

assign G = ~(~gouta[1] & ~(pouta[1] & gouta[0]));
assign P = pouta[1] & pouta[0];

endmodule // fcla8


//////////////////////////////////////////////////////////////////////////////// 

`timescale 1ns / 1ps

module REG_BYPASS_MUX(D, Q, ENA, CLK, RST, SELM);

parameter DATA_WIDTH = 16 ;

input  [DATA_WIDTH - 1 : 0] D ;
output [DATA_WIDTH - 1 : 0] Q ;
input  ENA ;
input  CLK ;
input  RST ;
input  SELM ;

reg    [DATA_WIDTH - 1 : 0] REG_INTERNAL ;

assign Q = ( (SELM) ? REG_INTERNAL : D ) ;

always @ (posedge CLK or posedge RST)
begin
	if (RST)
		REG_INTERNAL <= #1 0 ;
	else if (ENA)
	    REG_INTERNAL <= #1 D ;
	else 
	    REG_INTERNAL <= #1 REG_INTERNAL ;
end

endmodule

