`timescale 1 ps/1 ps
module ibex_top(\u_ibex_core/ex_block_i/adder_in_a(24) ,new_n16__8507_RESYNTH,\u_ibex_core/ex_block_i/adder_in_a(22) ,\u_ibex_core/ex_block_i/adder_in_a(16) ,\u_ibex_core/ex_block_i/adder_in_a(31) ,\u_ibex_core/ex_block_i/adder_in_a(26) ,new_n16__8619_RESYNTH,\u_ibex_core/ex_block_i/adder_in_a(8) ,new_n16__8357_RESYNTH,new_n16__8249_RESYNTH,new_n16__8299_RESYNTH,\u_ibex_core/ex_block_i/adder_in_a(30) ,adder_result_ext_o_carry_i_8_n_0,\u_ibex_core/ex_block_i/adder_in_a(6) ,\u_ibex_core/ex_block_i/adder_in_a(9) ,\u_ibex_core/ex_block_i/adder_in_a(29) ,\u_ibex_core/ex_block_i/adder_in_a(27) ,adder_result_ext_o_carry__7_i_1_n_0,\u_ibex_core/ex_block_i/adder_in_a(19) ,\u_ibex_core/ex_block_i/adder_in_a(14) ,new_n16__8497_RESYNTH,new_n16__8441_RESYNTH,\u_ibex_core/ex_block_i/adder_in_a(28) ,\u_ibex_core/ex_block_i/adder_in_a(25) ,new_n16__8377_RESYNTH,new_n16__8411_RESYNTH,new_n16__8517_RESYNTH,\u_ibex_core/ex_block_i/adder_in_a(5) ,\u_ibex_core/ex_block_i/adder_in_a(4) ,\u_ibex_core/ex_block_i/adder_in_a(17) ,\u_ibex_core/ex_block_i/adder_in_a(12) ,new_n16__8347_RESYNTH,\u_ibex_core/ex_block_i/adder_in_a(15) ,new_n16__8557_RESYNTH,\u_ibex_core/ex_block_i/adder_in_a(23) ,\u_ibex_core/ex_block_i/adder_in_a(20) ,\u_ibex_core/ex_block_i/adder_in_a(21) ,new_n16__8527_RESYNTH,new_n16__8259_RESYNTH,\u_ibex_core/ex_block_i/adder_in_a(11) ,new_n16__8367_RESYNTH,new_n16__8467_RESYNTH,\u_ibex_core/ex_block_i/adder_in_a(1) ,\u_ibex_core/ex_block_i/adder_in_a(13) ,new_n16__8421_RESYNTH,\u_ibex_core/ex_block_i/adder_in_a(10) ,\u_ibex_core/ex_block_i/adder_in_a(18) ,new_n16__8537_RESYNTH,\u_ibex_core/ex_block_i/adder_in_a(2) ,new_n16__8477_RESYNTH,\u_ibex_core/ex_block_i/adder_in_b(0) ,new_n16__8487_RESYNTH,new_n16__8431_RESYNTH,\u_ibex_core/ex_block_i/adder_in_a(7) ,new_n16__8457_RESYNTH,new_n16__8309_RESYNTH,new_n16__8651_RESYNTH,\u_ibex_core/ex_block_i/adder_in_a(3) ,new_n16__8547_RESYNTH,new_n16__8567_RESYNTH,new_n16__8661_RESYNTH,new_n16__8319_RESYNTH,new_n16__8289_RESYNTH,new_n16__8279_RESYNTH,new_n16__8269_RESYNTH,\data_addr_o(10) ,\u_ibex_core/alu_adder_result_ex(0) ,\data_addr_o(20) ,\data_addr_o(27) ,\data_addr_o(28) ,\data_addr_o(23) ,\data_addr_o(6) ,\data_addr_o(30) ,\data_addr_o(4) ,\data_addr_o(31) ,\data_addr_o(25) ,\data_addr_o(11) ,\data_addr_o(21) ,\data_addr_o(7) ,\data_addr_o(13) ,\data_addr_o(2) ,\data_addr_o(8) ,\data_addr_o(17) ,\data_addr_o(9) ,\data_addr_o(29) ,\data_addr_o(26) ,\data_addr_o(19) ,\data_addr_o(12) ,\data_addr_o(24) ,\data_addr_o(5) ,\data_addr_o(15) ,\data_addr_o(18) ,\data_addr_o(14) ,\data_addr_o(16) ,\u_ibex_core/alu_adder_result_ex(1) ,\data_addr_o(22) ,\data_addr_o(3) );
    input \u_ibex_core/ex_block_i/adder_in_a(24) ;
    input new_n16__8507_RESYNTH;
    input \u_ibex_core/ex_block_i/adder_in_a(22) ;
    input \u_ibex_core/ex_block_i/adder_in_a(16) ;
    input \u_ibex_core/ex_block_i/adder_in_a(31) ;
    input \u_ibex_core/ex_block_i/adder_in_a(26) ;
    input new_n16__8619_RESYNTH;
    input \u_ibex_core/ex_block_i/adder_in_a(8) ;
    input new_n16__8357_RESYNTH;
    input new_n16__8249_RESYNTH;
    input new_n16__8299_RESYNTH;
    input \u_ibex_core/ex_block_i/adder_in_a(30) ;
    input adder_result_ext_o_carry_i_8_n_0;
    input \u_ibex_core/ex_block_i/adder_in_a(6) ;
    input \u_ibex_core/ex_block_i/adder_in_a(9) ;
    input \u_ibex_core/ex_block_i/adder_in_a(29) ;
    input \u_ibex_core/ex_block_i/adder_in_a(27) ;
    input adder_result_ext_o_carry__7_i_1_n_0;
    input \u_ibex_core/ex_block_i/adder_in_a(19) ;
    input \u_ibex_core/ex_block_i/adder_in_a(14) ;
    input new_n16__8497_RESYNTH;
    input new_n16__8441_RESYNTH;
    input \u_ibex_core/ex_block_i/adder_in_a(28) ;
    input \u_ibex_core/ex_block_i/adder_in_a(25) ;
    input new_n16__8377_RESYNTH;
    input new_n16__8411_RESYNTH;
    input new_n16__8517_RESYNTH;
    input \u_ibex_core/ex_block_i/adder_in_a(5) ;
    input \u_ibex_core/ex_block_i/adder_in_a(4) ;
    input \u_ibex_core/ex_block_i/adder_in_a(17) ;
    input \u_ibex_core/ex_block_i/adder_in_a(12) ;
    input new_n16__8347_RESYNTH;
    input \u_ibex_core/ex_block_i/adder_in_a(15) ;
    input new_n16__8557_RESYNTH;
    input \u_ibex_core/ex_block_i/adder_in_a(23) ;
    input \u_ibex_core/ex_block_i/adder_in_a(20) ;
    input \u_ibex_core/ex_block_i/adder_in_a(21) ;
    input new_n16__8527_RESYNTH;
    input new_n16__8259_RESYNTH;
    input \u_ibex_core/ex_block_i/adder_in_a(11) ;
    input new_n16__8367_RESYNTH;
    input new_n16__8467_RESYNTH;
    input \u_ibex_core/ex_block_i/adder_in_a(1) ;
    input \u_ibex_core/ex_block_i/adder_in_a(13) ;
    input new_n16__8421_RESYNTH;
    input \u_ibex_core/ex_block_i/adder_in_a(10) ;
    input \u_ibex_core/ex_block_i/adder_in_a(18) ;
    input new_n16__8537_RESYNTH;
    input \u_ibex_core/ex_block_i/adder_in_a(2) ;
    input new_n16__8477_RESYNTH;
    input \u_ibex_core/ex_block_i/adder_in_b(0) ;
    input new_n16__8487_RESYNTH;
    input new_n16__8431_RESYNTH;
    input \u_ibex_core/ex_block_i/adder_in_a(7) ;
    input new_n16__8457_RESYNTH;
    input new_n16__8309_RESYNTH;
    input new_n16__8651_RESYNTH;
    input \u_ibex_core/ex_block_i/adder_in_a(3) ;
    input new_n16__8547_RESYNTH;
    input new_n16__8567_RESYNTH;
    input new_n16__8661_RESYNTH;
    input new_n16__8319_RESYNTH;
    input new_n16__8289_RESYNTH;
    input new_n16__8279_RESYNTH;
    input new_n16__8269_RESYNTH;
    output \data_addr_o(10) ;
    output \u_ibex_core/alu_adder_result_ex(0) ;
    output \data_addr_o(20) ;
    output \data_addr_o(27) ;
    output \data_addr_o(28) ;
    output \data_addr_o(23) ;
    output \data_addr_o(6) ;
    output \data_addr_o(30) ;
    output \data_addr_o(4) ;
    output \data_addr_o(31) ;
    output \data_addr_o(25) ;
    output \data_addr_o(11) ;
    output \data_addr_o(21) ;
    output \data_addr_o(7) ;
    output \data_addr_o(13) ;
    output \data_addr_o(2) ;
    output \data_addr_o(8) ;
    output \data_addr_o(17) ;
    output \data_addr_o(9) ;
    output \data_addr_o(29) ;
    output \data_addr_o(26) ;
    output \data_addr_o(19) ;
    output \data_addr_o(12) ;
    output \data_addr_o(24) ;
    output \data_addr_o(5) ;
    output \data_addr_o(15) ;
    output \data_addr_o(18) ;
    output \data_addr_o(14) ;
    output \data_addr_o(16) ;
    output \u_ibex_core/alu_adder_result_ex(1) ;
    output \data_addr_o(22) ;
    output \data_addr_o(3) ;
    wire adder_result_ext_o_carry__3_i_8_n_0;
    wire \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__0_n_3 ;
    wire adder_result_ext_o_carry__5_i_6_n_0;
    wire \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry_n_0 ;
    wire new_n7__8291_RESYNTH;
    wire adder_result_ext_o_carry__4_i_5_n_0;
    wire \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__5_n_0 ;
    wire new_n7__8459_RESYNTH;
    wire adder_result_ext_o_carry__2_i_6_n_0;
    wire new_n7__8301_RESYNTH;
    wire adder_result_ext_o_carry__5_i_7_n_0;
    wire adder_result_ext_o_carry__4_i_7_n_0;
    wire \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__3_n_1 ;
    wire adder_result_ext_o_carry__5_i_8_n_0;
    wire adder_result_ext_o_carry__1_i_5_n_0;
    wire new_n7__8653_RESYNTH;
    wire \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__0_n_0 ;
    wire \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__2_n_3 ;
    wire \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__4_n_0 ;
    wire adder_result_ext_o_carry__2_i_7_n_0;
    wire \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__5_n_1 ;
    wire adder_result_ext_o_carry_i_7_n_0;
    wire new_n7__8349_RESYNTH;
    wire \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__5_n_2 ;
    wire adder_result_ext_o_carry__3_i_5_n_0;
    wire \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__2_n_0 ;
    wire \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__5_n_3 ;
    wire new_n7__8559_RESYNTH;
    wire \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__0_n_2 ;
    wire \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__6_n_2 ;
    wire adder_result_ext_o_carry__1_i_6_n_0;
    wire adder_result_ext_o_carry__5_i_5_n_0;
    wire \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__6_n_3 ;
    wire new_n7__8519_RESYNTH;
    wire adder_result_ext_o_carry__6_i_6_n_0;
    wire new_n7__8509_RESYNTH;
    wire new_n7__8469_RESYNTH;
    wire \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__2_n_2 ;
    wire new_n7__8369_RESYNTH;
    wire new_n7__8281_RESYNTH;
    wire new_n7__8489_RESYNTH;
    wire \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__6_n_1 ;
    wire new_n7__8311_RESYNTH;
    wire new_n7__8479_RESYNTH;
    wire new_n7__8321_RESYNTH;
    wire adder_result_ext_o_carry_i_5_n_0;
    wire new_n7__8443_RESYNTH;
    wire adder_result_ext_o_carry__4_i_6_n_0;
    wire adder_result_ext_o_carry__0_i_5_n_0;
    wire adder_result_ext_o_carry__6_i_7_n_0;
    wire new_n7__8261_RESYNTH;
    wire new_n7__8359_RESYNTH;
    wire \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__6_n_0 ;
    wire adder_result_ext_o_carry__1_i_7_n_0;
    wire new_n7__8499_RESYNTH;
    wire new_n7__8379_RESYNTH;
    wire new_n7__8569_RESYNTH;
    wire \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__1_n_1 ;
    wire new_n7__8423_RESYNTH;
    wire adder_result_ext_o_carry__6_i_5_n_0;
    wire adder_result_ext_o_carry__6_i_8_n_0;
    wire adder_result_ext_o_carry__0_i_8_n_0;
    wire new_n7__8413_RESYNTH;
    wire new_n7__8549_RESYNTH;
    wire new_n7__8433_RESYNTH;
    wire new_n7__8271_RESYNTH;
    wire adder_result_ext_o_carry__3_i_6_n_0;
    wire new_n7__8621_RESYNTH;
    wire new_n7__8663_RESYNTH;
    wire adder_result_ext_o_carry__0_i_7_n_0;
    wire \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__4_n_2 ;
    wire \NLW_u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry_O_UNCONNECTED(0) ;
    wire \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__1_n_0 ;
    wire adder_result_ext_o_carry__2_i_8_n_0;
    wire \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry_n_2 ;
    wire adder_result_ext_o_carry__3_i_7_n_0;
    wire \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__0_n_1 ;
    wire adder_result_ext_o_carry__4_i_8_n_0;
    wire \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__4_n_3 ;
    wire adder_result_ext_o_carry__1_i_8_n_0;
    wire new_n7__8539_RESYNTH;
    wire adder_result_ext_o_carry__0_i_6_n_0;
    wire \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__3_n_3 ;
    wire new_n7__8251_RESYNTH;
    wire \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry_n_3 ;
    wire \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__1_n_3 ;
    wire \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__1_n_2 ;
    wire adder_result_ext_o_carry_i_6_n_0;
    wire \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry_n_1 ;
    wire \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__4_n_1 ;
    wire new_n7__8529_RESYNTH;
    wire \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__3_n_2 ;
    wire \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__2_n_1 ;
    wire adder_result_ext_o_carry__2_i_5_n_0;
    wire \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__3_n_0 ;

    HAL_XOR2 g10_4783_RESYNTH (
        .A(new_n16__8457_RESYNTH),
        .B(new_n7__8459_RESYNTH),
        .O(adder_result_ext_o_carry__4_i_5_n_0)
    );

    HAL_INV g00_1643_RESYNTH (
        .A(\u_ibex_core/ex_block_i/adder_in_a(9) ),
        .O(new_n7__8311_RESYNTH)
    );

    HAL_XOR2 g10_1638_RESYNTH (
        .A(new_n16__8299_RESYNTH),
        .B(new_n7__8301_RESYNTH),
        .O(adder_result_ext_o_carry__1_i_6_n_0)
    );

    HAL_XOR2 g10_7990_RESYNTH (
        .A(new_n16__8557_RESYNTH),
        .B(new_n7__8559_RESYNTH),
        .O(adder_result_ext_o_carry__6_i_7_n_0)
    );

    HAL_INV g00_7991_RESYNTH (
        .A(\u_ibex_core/ex_block_i/adder_in_a(28) ),
        .O(new_n7__8569_RESYNTH)
    );

    HAL_XOR2 g10_2127_RESYNTH (
        .A(new_n16__8357_RESYNTH),
        .B(new_n7__8359_RESYNTH),
        .O(adder_result_ext_o_carry__2_i_6_n_0)
    );

    CARRY4 \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__5  (
        .CI(\u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__4_n_0 ),
        .CYINIT(1'b0 ),
        .DI({
            \u_ibex_core/ex_block_i/adder_in_a(27) ,
            \u_ibex_core/ex_block_i/adder_in_a(26) ,
            \u_ibex_core/ex_block_i/adder_in_a(25) ,
            \u_ibex_core/ex_block_i/adder_in_a(24) 
        }),
        .S({
            adder_result_ext_o_carry__5_i_5_n_0,
            adder_result_ext_o_carry__5_i_6_n_0,
            adder_result_ext_o_carry__5_i_7_n_0,
            adder_result_ext_o_carry__5_i_8_n_0
        }),
        .CO({
            \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__5_n_0 ,
            \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__5_n_1 ,
            \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__5_n_2 ,
            \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__5_n_3 
        }),
        .O({
            \data_addr_o(26) ,
            \data_addr_o(25) ,
            \data_addr_o(24) ,
            \data_addr_o(23) 
        })
    );

    CARRY4 \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__6  (
        .CI(\u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__5_n_0 ),
        .CYINIT(1'b0 ),
        .DI({
            \u_ibex_core/ex_block_i/adder_in_a(31) ,
            \u_ibex_core/ex_block_i/adder_in_a(30) ,
            \u_ibex_core/ex_block_i/adder_in_a(29) ,
            \u_ibex_core/ex_block_i/adder_in_a(28) 
        }),
        .S({
            adder_result_ext_o_carry__6_i_5_n_0,
            adder_result_ext_o_carry__6_i_6_n_0,
            adder_result_ext_o_carry__6_i_7_n_0,
            adder_result_ext_o_carry__6_i_8_n_0
        }),
        .CO({
            \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__6_n_0 ,
            \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__6_n_1 ,
            \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__6_n_2 ,
            \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__6_n_3 
        }),
        .O({
            \data_addr_o(30) ,
            \data_addr_o(29) ,
            \data_addr_o(28) ,
            \data_addr_o(27) 
        })
    );

    CARRY4 \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__7  (
        .CI(\u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__6_n_0 ),
        .CYINIT(1'b0 ),
        .DI({
            1'b0 ,
            1'b0 ,
            1'b0 ,
            1'b0 
        }),
        .S({
            1'b0 ,
            1'b0 ,
            1'b0 ,
            adder_result_ext_o_carry__7_i_1_n_0
        }),
        .O({
            1'bz,
            1'bz,
            1'bz,
            \data_addr_o(31) 
        })
    );

    HAL_INV g00_5158_RESYNTH (
        .A(\u_ibex_core/ex_block_i/adder_in_a(25) ),
        .O(new_n7__8519_RESYNTH)
    );

    HAL_XOR2 g10_5152_RESYNTH (
        .A(new_n16__8507_RESYNTH),
        .B(new_n7__8509_RESYNTH),
        .O(adder_result_ext_o_carry__5_i_6_n_0)
    );

    HAL_INV g00_4785_RESYNTH (
        .A(\u_ibex_core/ex_block_i/adder_in_a(22) ),
        .O(new_n7__8469_RESYNTH)
    );

    HAL_XOR2 g10_8001_RESYNTH (
        .A(new_n16__8567_RESYNTH),
        .B(new_n7__8569_RESYNTH),
        .O(adder_result_ext_o_carry__6_i_8_n_0)
    );

    HAL_INV g00_4919_RESYNTH (
        .A(\u_ibex_core/ex_block_i/adder_in_a(20) ),
        .O(new_n7__8489_RESYNTH)
    );

    HAL_XOR2 g10_4912_RESYNTH (
        .A(new_n16__8477_RESYNTH),
        .B(new_n7__8479_RESYNTH),
        .O(adder_result_ext_o_carry__4_i_7_n_0)
    );

    HAL_INV g00_423_RESYNTH (
        .A(\u_ibex_core/ex_block_i/adder_in_a(7) ),
        .O(new_n7__8251_RESYNTH)
    );

    HAL_XOR2 g10_5070_RESYNTH (
        .A(new_n16__8497_RESYNTH),
        .B(new_n7__8499_RESYNTH),
        .O(adder_result_ext_o_carry__5_i_5_n_0)
    );

    HAL_INV g00_1694_RESYNTH (
        .A(\u_ibex_core/ex_block_i/adder_in_a(8) ),
        .O(new_n7__8321_RESYNTH)
    );

    HAL_XOR2 g10_4683_RESYNTH (
        .A(new_n16__8441_RESYNTH),
        .B(new_n7__8443_RESYNTH),
        .O(adder_result_ext_o_carry__3_i_8_n_0)
    );

    HAL_INV g00_445_RESYNTH (
        .A(\u_ibex_core/ex_block_i/adder_in_a(6) ),
        .O(new_n7__8261_RESYNTH)
    );

    HAL_INV g00_2154_RESYNTH (
        .A(\u_ibex_core/ex_block_i/adder_in_a(13) ),
        .O(new_n7__8369_RESYNTH)
    );

    HAL_XOR2 g10_1685_RESYNTH (
        .A(new_n16__8309_RESYNTH),
        .B(new_n7__8311_RESYNTH),
        .O(adder_result_ext_o_carry__1_i_7_n_0)
    );

    HAL_XOR2 g10_443_RESYNTH (
        .A(new_n16__8249_RESYNTH),
        .B(new_n7__8251_RESYNTH),
        .O(adder_result_ext_o_carry__0_i_5_n_0)
    );

    HAL_INV g00_2274_RESYNTH (
        .A(\u_ibex_core/ex_block_i/adder_in_a(12) ),
        .O(new_n7__8379_RESYNTH)
    );

    HAL_XOR2 g10_4560_RESYNTH (
        .A(new_n16__8421_RESYNTH),
        .B(new_n7__8423_RESYNTH),
        .O(adder_result_ext_o_carry__3_i_6_n_0)
    );

    HAL_INV g00_5084_RESYNTH (
        .A(\u_ibex_core/ex_block_i/adder_in_a(26) ),
        .O(new_n7__8509_RESYNTH)
    );

    HAL_INV g00_4563_RESYNTH (
        .A(\u_ibex_core/ex_block_i/adder_in_a(17) ),
        .O(new_n7__8433_RESYNTH)
    );

    HAL_XOR2 g10_1580_RESYNTH (
        .A(new_n16__8289_RESYNTH),
        .B(new_n7__8291_RESYNTH),
        .O(adder_result_ext_o_carry__1_i_5_n_0)
    );

    HAL_INV g00_1939_RESYNTH (
        .A(\u_ibex_core/ex_block_i/adder_in_a(15) ),
        .O(new_n7__8349_RESYNTH)
    );

    HAL_XOR2 g10_8062_RESYNTH (
        .A(new_n16__8619_RESYNTH),
        .B(new_n7__8621_RESYNTH),
        .O(adder_result_ext_o_carry_i_5_n_0)
    );

    HAL_INV g00_8052_RESYNTH (
        .A(\u_ibex_core/ex_block_i/adder_in_a(3) ),
        .O(new_n7__8621_RESYNTH)
    );

    HAL_XOR2 g10_2056_RESYNTH (
        .A(new_n16__8347_RESYNTH),
        .B(new_n7__8349_RESYNTH),
        .O(adder_result_ext_o_carry__2_i_5_n_0)
    );

    HAL_XOR2 g10_1456_RESYNTH (
        .A(new_n16__8279_RESYNTH),
        .B(new_n7__8281_RESYNTH),
        .O(adder_result_ext_o_carry__0_i_8_n_0)
    );

    HAL_XOR2 g10_4343_RESYNTH (
        .A(new_n16__8411_RESYNTH),
        .B(new_n7__8413_RESYNTH),
        .O(adder_result_ext_o_carry__3_i_5_n_0)
    );

    HAL_XOR2 g10_472_RESYNTH (
        .A(new_n16__8259_RESYNTH),
        .B(new_n7__8261_RESYNTH),
        .O(adder_result_ext_o_carry__0_i_6_n_0)
    );

    HAL_INV g00_473_RESYNTH (
        .A(\u_ibex_core/ex_block_i/adder_in_a(5) ),
        .O(new_n7__8271_RESYNTH)
    );

    HAL_INV g00_4856_RESYNTH (
        .A(\u_ibex_core/ex_block_i/adder_in_a(21) ),
        .O(new_n7__8479_RESYNTH)
    );

    HAL_XOR2 g10_7946_RESYNTH (
        .A(new_n16__8517_RESYNTH),
        .B(new_n7__8519_RESYNTH),
        .O(adder_result_ext_o_carry__5_i_7_n_0)
    );

    HAL_INV g00_1584_RESYNTH (
        .A(\u_ibex_core/ex_block_i/adder_in_a(10) ),
        .O(new_n7__8301_RESYNTH)
    );

    HAL_INV g00_7947_RESYNTH (
        .A(\u_ibex_core/ex_block_i/adder_in_a(24) ),
        .O(new_n7__8529_RESYNTH)
    );

    HAL_INV g00_4232_RESYNTH (
        .A(\u_ibex_core/ex_block_i/adder_in_a(19) ),
        .O(new_n7__8413_RESYNTH)
    );

    HAL_INV g00_1487_RESYNTH (
        .A(\u_ibex_core/ex_block_i/adder_in_a(11) ),
        .O(new_n7__8291_RESYNTH)
    );

    HAL_INV g00_4730_RESYNTH (
        .A(\u_ibex_core/ex_block_i/adder_in_a(23) ),
        .O(new_n7__8459_RESYNTH)
    );

    HAL_XOR2 g10_4849_RESYNTH (
        .A(new_n16__8467_RESYNTH),
        .B(new_n7__8469_RESYNTH),
        .O(adder_result_ext_o_carry__4_i_6_n_0)
    );

    HAL_XOR2 g10_1245_RESYNTH (
        .A(new_n16__8269_RESYNTH),
        .B(new_n7__8271_RESYNTH),
        .O(adder_result_ext_o_carry__0_i_7_n_0)
    );

    HAL_INV g00_8088_RESYNTH (
        .A(\u_ibex_core/ex_block_i/adder_in_a(2) ),
        .O(new_n7__8653_RESYNTH)
    );

    HAL_INV g00_4622_RESYNTH (
        .A(\u_ibex_core/ex_block_i/adder_in_a(16) ),
        .O(new_n7__8443_RESYNTH)
    );

    HAL_XOR2 g10_2220_RESYNTH (
        .A(new_n16__8367_RESYNTH),
        .B(new_n7__8369_RESYNTH),
        .O(adder_result_ext_o_carry__2_i_7_n_0)
    );

    HAL_INV g00_2065_RESYNTH (
        .A(\u_ibex_core/ex_block_i/adder_in_a(14) ),
        .O(new_n7__8359_RESYNTH)
    );

    HAL_INV g00_5007_RESYNTH (
        .A(\u_ibex_core/ex_block_i/adder_in_a(27) ),
        .O(new_n7__8499_RESYNTH)
    );

    HAL_XOR2 g10_7957_RESYNTH (
        .A(new_n16__8527_RESYNTH),
        .B(new_n7__8529_RESYNTH),
        .O(adder_result_ext_o_carry__5_i_8_n_0)
    );

    HAL_INV g00_4353_RESYNTH (
        .A(\u_ibex_core/ex_block_i/adder_in_a(18) ),
        .O(new_n7__8423_RESYNTH)
    );

    HAL_INV g00_7958_RESYNTH (
        .A(\u_ibex_core/ex_block_i/adder_in_a(31) ),
        .O(new_n7__8539_RESYNTH)
    );

    HAL_XOR2 g10_2586_RESYNTH (
        .A(new_n16__8377_RESYNTH),
        .B(new_n7__8379_RESYNTH),
        .O(adder_result_ext_o_carry__2_i_8_n_0)
    );

    HAL_XOR2 g10_4613_RESYNTH (
        .A(new_n16__8431_RESYNTH),
        .B(new_n7__8433_RESYNTH),
        .O(adder_result_ext_o_carry__3_i_7_n_0)
    );

    HAL_XOR2 g10_8109_RESYNTH (
        .A(new_n16__8661_RESYNTH),
        .B(new_n7__8663_RESYNTH),
        .O(adder_result_ext_o_carry_i_7_n_0)
    );

    HAL_INV g00_7980_RESYNTH (
        .A(\u_ibex_core/ex_block_i/adder_in_a(29) ),
        .O(new_n7__8559_RESYNTH)
    );

    HAL_XOR2 g10_4999_RESYNTH (
        .A(new_n16__8487_RESYNTH),
        .B(new_n7__8489_RESYNTH),
        .O(adder_result_ext_o_carry__4_i_8_n_0)
    );

    HAL_XOR2 g10_7979_RESYNTH (
        .A(new_n16__8547_RESYNTH),
        .B(new_n7__8549_RESYNTH),
        .O(adder_result_ext_o_carry__6_i_6_n_0)
    );

    CARRY4 \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__1  (
        .CI(\u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__0_n_0 ),
        .CYINIT(1'b0 ),
        .DI({
            \u_ibex_core/ex_block_i/adder_in_a(11) ,
            \u_ibex_core/ex_block_i/adder_in_a(10) ,
            \u_ibex_core/ex_block_i/adder_in_a(9) ,
            \u_ibex_core/ex_block_i/adder_in_a(8) 
        }),
        .S({
            adder_result_ext_o_carry__1_i_5_n_0,
            adder_result_ext_o_carry__1_i_6_n_0,
            adder_result_ext_o_carry__1_i_7_n_0,
            adder_result_ext_o_carry__1_i_8_n_0
        }),
        .CO({
            \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__1_n_0 ,
            \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__1_n_1 ,
            \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__1_n_2 ,
            \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__1_n_3 
        }),
        .O({
            \data_addr_o(10) ,
            \data_addr_o(9) ,
            \data_addr_o(8) ,
            \data_addr_o(7) 
        })
    );

    HAL_XOR2 g10_8098_RESYNTH (
        .A(new_n16__8651_RESYNTH),
        .B(new_n7__8653_RESYNTH),
        .O(adder_result_ext_o_carry_i_6_n_0)
    );

    CARRY4 \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__2  (
        .CI(\u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__1_n_0 ),
        .CYINIT(1'b0 ),
        .DI({
            \u_ibex_core/ex_block_i/adder_in_a(15) ,
            \u_ibex_core/ex_block_i/adder_in_a(14) ,
            \u_ibex_core/ex_block_i/adder_in_a(13) ,
            \u_ibex_core/ex_block_i/adder_in_a(12) 
        }),
        .S({
            adder_result_ext_o_carry__2_i_5_n_0,
            adder_result_ext_o_carry__2_i_6_n_0,
            adder_result_ext_o_carry__2_i_7_n_0,
            adder_result_ext_o_carry__2_i_8_n_0
        }),
        .CO({
            \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__2_n_0 ,
            \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__2_n_1 ,
            \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__2_n_2 ,
            \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__2_n_3 
        }),
        .O({
            \data_addr_o(14) ,
            \data_addr_o(13) ,
            \data_addr_o(12) ,
            \data_addr_o(11) 
        })
    );

    HAL_INV g00_8099_RESYNTH (
        .A(\u_ibex_core/ex_block_i/adder_in_a(1) ),
        .O(new_n7__8663_RESYNTH)
    );

    HAL_XOR2 g10_7968_RESYNTH (
        .A(new_n16__8537_RESYNTH),
        .B(new_n7__8539_RESYNTH),
        .O(adder_result_ext_o_carry__6_i_5_n_0)
    );

    HAL_INV g00_1250_RESYNTH (
        .A(\u_ibex_core/ex_block_i/adder_in_a(4) ),
        .O(new_n7__8281_RESYNTH)
    );

    CARRY4 \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__3  (
        .CI(\u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__2_n_0 ),
        .CYINIT(1'b0 ),
        .DI({
            \u_ibex_core/ex_block_i/adder_in_a(19) ,
            \u_ibex_core/ex_block_i/adder_in_a(18) ,
            \u_ibex_core/ex_block_i/adder_in_a(17) ,
            \u_ibex_core/ex_block_i/adder_in_a(16) 
        }),
        .S({
            adder_result_ext_o_carry__3_i_5_n_0,
            adder_result_ext_o_carry__3_i_6_n_0,
            adder_result_ext_o_carry__3_i_7_n_0,
            adder_result_ext_o_carry__3_i_8_n_0
        }),
        .CO({
            \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__3_n_0 ,
            \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__3_n_1 ,
            \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__3_n_2 ,
            \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__3_n_3 
        }),
        .O({
            \data_addr_o(18) ,
            \data_addr_o(17) ,
            \data_addr_o(16) ,
            \data_addr_o(15) 
        })
    );

    HAL_INV g00_7969_RESYNTH (
        .A(\u_ibex_core/ex_block_i/adder_in_a(30) ),
        .O(new_n7__8549_RESYNTH)
    );

    CARRY4 \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__4  (
        .CI(\u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__3_n_0 ),
        .CYINIT(1'b0 ),
        .DI({
            \u_ibex_core/ex_block_i/adder_in_a(23) ,
            \u_ibex_core/ex_block_i/adder_in_a(22) ,
            \u_ibex_core/ex_block_i/adder_in_a(21) ,
            \u_ibex_core/ex_block_i/adder_in_a(20) 
        }),
        .S({
            adder_result_ext_o_carry__4_i_5_n_0,
            adder_result_ext_o_carry__4_i_6_n_0,
            adder_result_ext_o_carry__4_i_7_n_0,
            adder_result_ext_o_carry__4_i_8_n_0
        }),
        .CO({
            \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__4_n_0 ,
            \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__4_n_1 ,
            \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__4_n_2 ,
            \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__4_n_3 
        }),
        .O({
            \data_addr_o(22) ,
            \data_addr_o(21) ,
            \data_addr_o(20) ,
            \data_addr_o(19) 
        })
    );

    HAL_XOR2 g10_1769_RESYNTH (
        .A(new_n16__8319_RESYNTH),
        .B(new_n7__8321_RESYNTH),
        .O(adder_result_ext_o_carry__1_i_8_n_0)
    );

    CARRY4 \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry  (
        .CI(1'b0 ),
        .CYINIT(1'b0 ),
        .DI({
            \u_ibex_core/ex_block_i/adder_in_a(3) ,
            \u_ibex_core/ex_block_i/adder_in_a(2) ,
            \u_ibex_core/ex_block_i/adder_in_a(1) ,
            \u_ibex_core/ex_block_i/adder_in_b(0) 
        }),
        .S({
            adder_result_ext_o_carry_i_5_n_0,
            adder_result_ext_o_carry_i_6_n_0,
            adder_result_ext_o_carry_i_7_n_0,
            adder_result_ext_o_carry_i_8_n_0
        }),
        .CO({
            \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry_n_0 ,
            \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry_n_1 ,
            \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry_n_2 ,
            \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry_n_3 
        }),
        .O({
            \data_addr_o(2) ,
            \u_ibex_core/alu_adder_result_ex(1) ,
            \u_ibex_core/alu_adder_result_ex(0) ,
            \NLW_u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry_O_UNCONNECTED(0) 
        })
    );

    CARRY4 \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__0  (
        .CI(\u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry_n_0 ),
        .CYINIT(1'b0 ),
        .DI({
            \u_ibex_core/ex_block_i/adder_in_a(7) ,
            \u_ibex_core/ex_block_i/adder_in_a(6) ,
            \u_ibex_core/ex_block_i/adder_in_a(5) ,
            \u_ibex_core/ex_block_i/adder_in_a(4) 
        }),
        .S({
            adder_result_ext_o_carry__0_i_5_n_0,
            adder_result_ext_o_carry__0_i_6_n_0,
            adder_result_ext_o_carry__0_i_7_n_0,
            adder_result_ext_o_carry__0_i_8_n_0
        }),
        .CO({
            \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__0_n_0 ,
            \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__0_n_1 ,
            \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__0_n_2 ,
            \u_ibex_core/ex_block_i/alu_i/adder_result_ext_o_carry__0_n_3 
        }),
        .O({
            \data_addr_o(6) ,
            \data_addr_o(5) ,
            \data_addr_o(4) ,
            \data_addr_o(3) 
        })
    );
endmodule

