`timescale 1 ps/1 ps
module top(\edge/pdata_2_3y(11) ,\edge/pdata_2_3y(9) ,\edge/pdata_2_3y(0) ,\edge/pdata_2_3y(18) ,\edge/pdata_2_3y(3) ,\edge/pdata_2_3y(16) ,\edge/pdata_2_3y(8) ,\edge/pdata_2_3y(2) ,\edge/pdata_2_3y(6) ,\edge/pdata_2_3y(4) ,\edge/pdata_2_3y(1) ,\edge/pdata_2_3y(14) ,\edge/pdata_2_3y(23) ,\edge/pdata_2_3y(10) ,\edge/pdata_2_3y(21) ,\edge/pdata_2_3y(19) ,\edge/pdata_2_3y(17) ,\edge/pdata_2_3y(15) ,\edge/pdata_2_3y(13) ,\edge/pdata_2_3y(12) ,\edge/pdata_2_3y(7) ,\edge/pdata_2_3y(20) ,\edge/pdata_2_3y(22) ,\edge/pdata_2_3y(5) ,\edge/filterV/plusOp101_out(29) ,\edge/filterV/plusOp101_out(27) ,\edge/filterV/plusOp101_out(18) ,\edge/filterV/plusOp101_out(25) ,\edge/filterV/plusOp101_out(23) ,\edge/filterV/plusOp101_out(31) ,\edge/filterV/plusOp101_out(30) ,\edge/filterV/plusOp101_out(17) ,\edge/filterV/plusOp101_out(9) ,\edge/filterV/plusOp101_out(12) ,\edge/filterV/plusOp101_out(7) ,\edge/filterV/plusOp101_out(11) ,\edge/filterV/plusOp101_out(22) ,\edge/filterV/plusOp101_out(21) ,\edge/filterV/plusOp101_out(8) ,\edge/filterV/plusOp101_out(20) ,\edge/filterV/plusOp101_out(26) ,\edge/filterV/plusOp101_out(13) ,\edge/filterV/plusOp101_out(28) ,\edge/filterV/plusOp101_out(15) ,\edge/filterV/plusOp101_out(16) ,\edge/filterV/plusOp101_out(14) ,\edge/filterV/plusOp101_out(10) ,\edge/filterV/plusOp101_out(24) ,\edge/filterV/plusOp101_out(19) );
    input \edge/pdata_2_3y(11) ;
    input \edge/pdata_2_3y(9) ;
    input \edge/pdata_2_3y(0) ;
    input \edge/pdata_2_3y(18) ;
    input \edge/pdata_2_3y(3) ;
    input \edge/pdata_2_3y(16) ;
    input \edge/pdata_2_3y(8) ;
    input \edge/pdata_2_3y(2) ;
    input \edge/pdata_2_3y(6) ;
    input \edge/pdata_2_3y(4) ;
    input \edge/pdata_2_3y(1) ;
    input \edge/pdata_2_3y(14) ;
    input \edge/pdata_2_3y(23) ;
    input \edge/pdata_2_3y(10) ;
    input \edge/pdata_2_3y(21) ;
    input \edge/pdata_2_3y(19) ;
    input \edge/pdata_2_3y(17) ;
    input \edge/pdata_2_3y(15) ;
    input \edge/pdata_2_3y(13) ;
    input \edge/pdata_2_3y(12) ;
    input \edge/pdata_2_3y(7) ;
    input \edge/pdata_2_3y(20) ;
    input \edge/pdata_2_3y(22) ;
    input \edge/pdata_2_3y(5) ;
    output \edge/filterV/plusOp101_out(29) ;
    output \edge/filterV/plusOp101_out(27) ;
    output \edge/filterV/plusOp101_out(18) ;
    output \edge/filterV/plusOp101_out(25) ;
    output \edge/filterV/plusOp101_out(23) ;
    output \edge/filterV/plusOp101_out(31) ;
    output \edge/filterV/plusOp101_out(30) ;
    output \edge/filterV/plusOp101_out(17) ;
    output \edge/filterV/plusOp101_out(9) ;
    output \edge/filterV/plusOp101_out(12) ;
    output \edge/filterV/plusOp101_out(7) ;
    output \edge/filterV/plusOp101_out(11) ;
    output \edge/filterV/plusOp101_out(22) ;
    output \edge/filterV/plusOp101_out(21) ;
    output \edge/filterV/plusOp101_out(8) ;
    output \edge/filterV/plusOp101_out(20) ;
    output \edge/filterV/plusOp101_out(26) ;
    output \edge/filterV/plusOp101_out(13) ;
    output \edge/filterV/plusOp101_out(28) ;
    output \edge/filterV/plusOp101_out(15) ;
    output \edge/filterV/plusOp101_out(16) ;
    output \edge/filterV/plusOp101_out(14) ;
    output \edge/filterV/plusOp101_out(10) ;
    output \edge/filterV/plusOp101_out(24) ;
    output \edge/filterV/plusOp101_out(19) ;
    wire \p2ya_reg[18]_i_1_n_2 ;
    wire \p2ya[31]_i_2_n_0 ;
    wire \p2ya_reg[18]_i_1_n_1 ;
    wire \p2ya[30]_i_5_n_0 ;
    wire \p2ya_reg[18]_i_1_n_0 ;
    wire \p2ya[30]_i_4_n_0 ;
    wire \p2ya[18]_i_4_n_0 ;
    wire \p2ya_reg[10]_i_1_n_0 ;
    wire \p2ya[18]_i_2_n_0 ;
    wire \p2ya[10]_i_3_n_0 ;
    wire \p2ya_reg[14]_i_1__0_n_0 ;
    wire \p2ya[26]_i_4_n_0 ;
    wire \p2ya[14]_i_4_n_0 ;
    wire \p2ya_reg[18]_i_1_n_3 ;
    wire \p2ya[14]_i_2_n_0 ;
    wire \p2ya_reg[10]_i_1_n_3 ;
    wire \p2ya[22]_i_3_n_0 ;
    wire \p2ya_reg[10]_i_1_n_2 ;
    wire \p2ya[22]_i_2_n_0 ;
    wire \p2ya_reg[10]_i_1_n_1 ;
    wire \p2ya[18]_i_5_n_0 ;
    wire \p2ya_reg[14]_i_1__0_n_1 ;
    wire \p2ya[26]_i_5_n_0 ;
    wire \p2ya[10]_i_2_n_0 ;
    wire \p2ya_reg[30]_i_1_n_1 ;
    wire \p2ya[26]_i_3_n_0 ;
    wire \p2ya_reg[22]_i_1_n_2 ;
    wire \p2ya[14]_i_5_n_0 ;
    wire \p2ya_reg[22]_i_1_n_0 ;
    wire \p2ya_reg[30]_i_1_n_0 ;
    wire \p2ya[18]_i_3_n_0 ;
    wire \p2ya_reg[26]_i_1_n_0 ;
    wire \p2ya_reg[26]_i_1_n_3 ;
    wire \p2ya_reg[26]_i_1_n_2 ;
    wire \p2ya_reg[26]_i_1_n_1 ;
    wire \p2ya[26]_i_2_n_0 ;
    wire \p2ya_reg[30]_i_1_n_3 ;
    wire \p2ya[22]_i_5_n_0 ;
    wire \p2ya_reg[30]_i_1_n_2 ;
    wire \p2ya[14]_i_3_n_0 ;
    wire \p2ya_reg[22]_i_1_n_3 ;
    wire \p2ya_reg[22]_i_1_n_1 ;
    wire \p2ya[30]_i_2_n_0 ;
    wire \p2ya_reg[14]_i_1__0_n_2 ;
    wire \p2ya[10]_i_4_n_0 ;
    wire \p2ya[30]_i_3_n_0 ;
    wire \p2ya_reg[14]_i_1__0_n_3 ;
    wire \p2ya[22]_i_4_n_0 ;

    HAL_INV _4749__11_NEW_GATE (
        .A(\edge/pdata_2_3y(1) ),
        .O(\p2ya[10]_i_4_n_0 )
    );

    HAL_XNOR2 _4892__5711_NEW_GATE (
        .A(\edge/pdata_2_3y(4) ),
        .B(\edge/pdata_2_3y(6) ),
        .O(\p2ya[14]_i_3_n_0 )
    );

    HAL_XNOR2 _4894__5713_NEW_GATE (
        .A(\edge/pdata_2_3y(4) ),
        .B(\edge/pdata_2_3y(2) ),
        .O(\p2ya[14]_i_5_n_0 )
    );

    HAL_XNOR2 _4900__5719_NEW_GATE (
        .A(\edge/pdata_2_3y(16) ),
        .B(\edge/pdata_2_3y(18) ),
        .O(\p2ya[26]_i_3_n_0 )
    );

    HAL_XNOR2 _4915__5818_NEW_GATE (
        .A(\edge/pdata_2_3y(3) ),
        .B(\edge/pdata_2_3y(1) ),
        .O(\p2ya[10]_i_2_n_0 )
    );

    HAL_XNOR2 _4947__5861_NEW_GATE (
        .A(\edge/pdata_2_3y(6) ),
        .B(\edge/pdata_2_3y(8) ),
        .O(\p2ya[18]_i_5_n_0 )
    );

    HAL_XNOR2 _4959__5873_NEW_GATE (
        .A(\edge/pdata_2_3y(16) ),
        .B(\edge/pdata_2_3y(14) ),
        .O(\p2ya[26]_i_5_n_0 )
    );

    HAL_XNOR2 _4960__5874_NEW_GATE (
        .A(\edge/pdata_2_3y(20) ),
        .B(\edge/pdata_2_3y(22) ),
        .O(\p2ya[30]_i_3_n_0 )
    );

    HAL_XNOR2 _4962__5876_NEW_GATE (
        .A(\edge/pdata_2_3y(14) ),
        .B(\edge/pdata_2_3y(12) ),
        .O(\p2ya[22]_i_3_n_0 )
    );

    HAL_XNOR2 _4964__5878_NEW_GATE (
        .A(\edge/pdata_2_3y(8) ),
        .B(\edge/pdata_2_3y(10) ),
        .O(\p2ya[18]_i_3_n_0 )
    );

    CARRY4 \p2ya_reg[10]_i_1  (
        .CI(1'b0 ),
        .CYINIT(1'b0 ),
        .DI({
            \edge/pdata_2_3y(1) ,
            \edge/pdata_2_3y(0) ,
            1'b0 ,
            1'b1 
        }),
        .S({
            \p2ya[10]_i_2_n_0 ,
            \p2ya[10]_i_3_n_0 ,
            \p2ya[10]_i_4_n_0 ,
            \edge/pdata_2_3y(0) 
        }),
        .CO({
            \p2ya_reg[10]_i_1_n_0 ,
            \p2ya_reg[10]_i_1_n_1 ,
            \p2ya_reg[10]_i_1_n_2 ,
            \p2ya_reg[10]_i_1_n_3 
        }),
        .O({
            \edge/filterV/plusOp101_out(10) ,
            \edge/filterV/plusOp101_out(9) ,
            \edge/filterV/plusOp101_out(8) ,
            \edge/filterV/plusOp101_out(7) 
        })
    );

    CARRY4 \p2ya_reg[14]_i_1__0  (
        .CI(\p2ya_reg[10]_i_1_n_0 ),
        .CYINIT(1'b0 ),
        .DI({
            \edge/pdata_2_3y(5) ,
            \edge/pdata_2_3y(4) ,
            \edge/pdata_2_3y(3) ,
            \edge/pdata_2_3y(2) 
        }),
        .S({
            \p2ya[14]_i_2_n_0 ,
            \p2ya[14]_i_3_n_0 ,
            \p2ya[14]_i_4_n_0 ,
            \p2ya[14]_i_5_n_0 
        }),
        .CO({
            \p2ya_reg[14]_i_1__0_n_0 ,
            \p2ya_reg[14]_i_1__0_n_1 ,
            \p2ya_reg[14]_i_1__0_n_2 ,
            \p2ya_reg[14]_i_1__0_n_3 
        }),
        .O({
            \edge/filterV/plusOp101_out(14) ,
            \edge/filterV/plusOp101_out(13) ,
            \edge/filterV/plusOp101_out(12) ,
            \edge/filterV/plusOp101_out(11) 
        })
    );

    CARRY4 \p2ya_reg[18]_i_1  (
        .CI(\p2ya_reg[14]_i_1__0_n_0 ),
        .CYINIT(1'b0 ),
        .DI({
            \edge/pdata_2_3y(9) ,
            \edge/pdata_2_3y(8) ,
            \edge/pdata_2_3y(7) ,
            \edge/pdata_2_3y(6) 
        }),
        .S({
            \p2ya[18]_i_2_n_0 ,
            \p2ya[18]_i_3_n_0 ,
            \p2ya[18]_i_4_n_0 ,
            \p2ya[18]_i_5_n_0 
        }),
        .CO({
            \p2ya_reg[18]_i_1_n_0 ,
            \p2ya_reg[18]_i_1_n_1 ,
            \p2ya_reg[18]_i_1_n_2 ,
            \p2ya_reg[18]_i_1_n_3 
        }),
        .O({
            \edge/filterV/plusOp101_out(18) ,
            \edge/filterV/plusOp101_out(17) ,
            \edge/filterV/plusOp101_out(16) ,
            \edge/filterV/plusOp101_out(15) 
        })
    );

    CARRY4 \p2ya_reg[22]_i_1  (
        .CI(\p2ya_reg[18]_i_1_n_0 ),
        .CYINIT(1'b0 ),
        .DI({
            \edge/pdata_2_3y(13) ,
            \edge/pdata_2_3y(12) ,
            \edge/pdata_2_3y(11) ,
            \edge/pdata_2_3y(10) 
        }),
        .S({
            \p2ya[22]_i_2_n_0 ,
            \p2ya[22]_i_3_n_0 ,
            \p2ya[22]_i_4_n_0 ,
            \p2ya[22]_i_5_n_0 
        }),
        .CO({
            \p2ya_reg[22]_i_1_n_0 ,
            \p2ya_reg[22]_i_1_n_1 ,
            \p2ya_reg[22]_i_1_n_2 ,
            \p2ya_reg[22]_i_1_n_3 
        }),
        .O({
            \edge/filterV/plusOp101_out(22) ,
            \edge/filterV/plusOp101_out(21) ,
            \edge/filterV/plusOp101_out(20) ,
            \edge/filterV/plusOp101_out(19) 
        })
    );

    CARRY4 \p2ya_reg[26]_i_1  (
        .CI(\p2ya_reg[22]_i_1_n_0 ),
        .CYINIT(1'b0 ),
        .DI({
            \edge/pdata_2_3y(17) ,
            \edge/pdata_2_3y(16) ,
            \edge/pdata_2_3y(15) ,
            \edge/pdata_2_3y(14) 
        }),
        .S({
            \p2ya[26]_i_2_n_0 ,
            \p2ya[26]_i_3_n_0 ,
            \p2ya[26]_i_4_n_0 ,
            \p2ya[26]_i_5_n_0 
        }),
        .CO({
            \p2ya_reg[26]_i_1_n_0 ,
            \p2ya_reg[26]_i_1_n_1 ,
            \p2ya_reg[26]_i_1_n_2 ,
            \p2ya_reg[26]_i_1_n_3 
        }),
        .O({
            \edge/filterV/plusOp101_out(26) ,
            \edge/filterV/plusOp101_out(25) ,
            \edge/filterV/plusOp101_out(24) ,
            \edge/filterV/plusOp101_out(23) 
        })
    );

    CARRY4 \p2ya_reg[30]_i_1  (
        .CI(\p2ya_reg[26]_i_1_n_0 ),
        .CYINIT(1'b0 ),
        .DI({
            \edge/pdata_2_3y(21) ,
            \edge/pdata_2_3y(20) ,
            \edge/pdata_2_3y(19) ,
            \edge/pdata_2_3y(18) 
        }),
        .S({
            \p2ya[30]_i_2_n_0 ,
            \p2ya[30]_i_3_n_0 ,
            \p2ya[30]_i_4_n_0 ,
            \p2ya[30]_i_5_n_0 
        }),
        .CO({
            \p2ya_reg[30]_i_1_n_0 ,
            \p2ya_reg[30]_i_1_n_1 ,
            \p2ya_reg[30]_i_1_n_2 ,
            \p2ya_reg[30]_i_1_n_3 
        }),
        .O({
            \edge/filterV/plusOp101_out(30) ,
            \edge/filterV/plusOp101_out(29) ,
            \edge/filterV/plusOp101_out(28) ,
            \edge/filterV/plusOp101_out(27) 
        })
    );

    CARRY4 \p2ya_reg[31]_i_1  (
        .CI(\p2ya_reg[30]_i_1_n_0 ),
        .CYINIT(1'b0 ),
        .DI({
            1'b0 ,
            1'b0 ,
            1'b0 ,
            1'b0 
        }),
        .S({
            1'b0 ,
            1'b0 ,
            1'b0 ,
            \p2ya[31]_i_2_n_0 
        }),
        .O({
            1'bz,
            1'bz,
            1'bz,
            \edge/filterV/plusOp101_out(31) 
        })
    );

    HAL_XNOR2 _4983__6199_NEW_GATE (
        .A(\edge/pdata_2_3y(22) ),
        .B(\edge/pdata_2_3y(23) ),
        .O(\p2ya[31]_i_2_n_0 )
    );

    HAL_XNOR2 _4985__6202_NEW_GATE (
        .A(\edge/pdata_2_3y(12) ),
        .B(\edge/pdata_2_3y(10) ),
        .O(\p2ya[22]_i_5_n_0 )
    );

    HAL_XNOR2 _4986__6271_NEW_GATE (
        .A(\edge/pdata_2_3y(18) ),
        .B(\edge/pdata_2_3y(20) ),
        .O(\p2ya[30]_i_5_n_0 )
    );

    HAL_XNOR2 _4998__6283_NEW_GATE (
        .A(\edge/pdata_2_3y(23) ),
        .B(\edge/pdata_2_3y(21) ),
        .O(\p2ya[30]_i_2_n_0 )
    );

    HAL_XNOR2 _5001__6286_NEW_GATE (
        .A(\edge/pdata_2_3y(3) ),
        .B(\edge/pdata_2_3y(5) ),
        .O(\p2ya[14]_i_4_n_0 )
    );

    HAL_XNOR2 _5017__6315_NEW_GATE (
        .A(\edge/pdata_2_3y(5) ),
        .B(\edge/pdata_2_3y(7) ),
        .O(\p2ya[14]_i_2_n_0 )
    );

    HAL_XNOR2 _5024__6322_NEW_GATE (
        .A(\edge/pdata_2_3y(17) ),
        .B(\edge/pdata_2_3y(19) ),
        .O(\p2ya[26]_i_2_n_0 )
    );

    HAL_XNOR2 _5032__6330_NEW_GATE (
        .A(\edge/pdata_2_3y(13) ),
        .B(\edge/pdata_2_3y(15) ),
        .O(\p2ya[22]_i_2_n_0 )
    );

    HAL_XNOR2 _5076__6589_NEW_GATE (
        .A(\edge/pdata_2_3y(17) ),
        .B(\edge/pdata_2_3y(15) ),
        .O(\p2ya[26]_i_4_n_0 )
    );

    HAL_XNOR2 _5077__6590_NEW_GATE (
        .A(\edge/pdata_2_3y(7) ),
        .B(\edge/pdata_2_3y(9) ),
        .O(\p2ya[18]_i_4_n_0 )
    );

    HAL_XNOR2 _5089__6636_NEW_GATE (
        .A(\edge/pdata_2_3y(21) ),
        .B(\edge/pdata_2_3y(19) ),
        .O(\p2ya[30]_i_4_n_0 )
    );

    HAL_XNOR2 _5090__6637_NEW_GATE (
        .A(\edge/pdata_2_3y(9) ),
        .B(\edge/pdata_2_3y(11) ),
        .O(\p2ya[18]_i_2_n_0 )
    );

    HAL_XNOR2 _5092__6639_NEW_GATE (
        .A(\edge/pdata_2_3y(2) ),
        .B(\edge/pdata_2_3y(0) ),
        .O(\p2ya[10]_i_3_n_0 )
    );

    HAL_XNOR2 _5104__6765_NEW_GATE (
        .A(\edge/pdata_2_3y(13) ),
        .B(\edge/pdata_2_3y(11) ),
        .O(\p2ya[22]_i_4_n_0 )
    );
endmodule

